magic
tech sky130A
magscale 1 2
timestamp 1586552775
<< viali >>
rect 1625 3545 1659 3579
rect 797 3477 831 3511
rect 1257 3477 1291 3511
rect 1809 3477 1843 3511
rect 2545 3409 2579 3443
rect 1441 3341 1475 3375
rect 2177 3273 2211 3307
rect 2361 3273 2395 3307
rect 889 3205 923 3239
rect 2085 3205 2119 3239
rect 1349 2865 1383 2899
rect 1717 2865 1751 2899
rect 2269 2865 2303 2899
rect 2821 2865 2855 2899
rect 797 2797 831 2831
rect 1165 2797 1199 2831
rect 1625 2797 1659 2831
rect 3005 2797 3039 2831
rect 2085 2661 2119 2695
rect 3189 2661 3223 2695
rect 797 2457 831 2491
rect 2913 2457 2947 2491
rect 3097 2457 3131 2491
rect 1073 2389 1107 2423
rect 3281 2321 3315 2355
rect 1993 2253 2027 2287
rect 2361 2253 2395 2287
rect 2637 2253 2671 2287
rect 3465 2253 3499 2287
rect 889 2185 923 2219
rect 1257 2117 1291 2151
rect 1441 2117 1475 2151
rect 1809 2117 1843 2151
rect 2269 2117 2303 2151
rect 3649 2117 3683 2151
rect 3005 1913 3039 1947
rect 3097 1913 3131 1947
rect 705 1777 739 1811
rect 1073 1709 1107 1743
rect 2453 1709 2487 1743
rect 3373 1641 3407 1675
rect 3557 1573 3591 1607
rect 3189 1233 3223 1267
rect 705 1165 739 1199
rect 1441 1165 1475 1199
rect 1809 1165 1843 1199
rect 981 1097 1015 1131
rect 1349 1029 1383 1063
rect 3649 1029 3683 1063
rect 3649 825 3683 859
rect 797 689 831 723
rect 3557 689 3591 723
rect 1165 621 1199 655
rect 2545 621 2579 655
rect 3097 553 3131 587
<< metal1 >>
rect 400 3690 4080 3712
rect 400 3638 1046 3690
rect 1098 3638 1110 3690
rect 1162 3638 1174 3690
rect 1226 3638 1238 3690
rect 1290 3638 1302 3690
rect 1354 3638 4080 3690
rect 400 3616 4080 3638
rect 1613 3579 1671 3585
rect 1613 3545 1625 3579
rect 1659 3576 1671 3579
rect 3174 3576 3180 3588
rect 1659 3548 3180 3576
rect 1659 3545 1671 3548
rect 1613 3539 1671 3545
rect 785 3511 843 3517
rect 785 3477 797 3511
rect 831 3508 843 3511
rect 1245 3511 1303 3517
rect 1245 3508 1257 3511
rect 831 3480 1257 3508
rect 831 3477 843 3480
rect 785 3471 843 3477
rect 1245 3477 1257 3480
rect 1291 3508 1303 3511
rect 1702 3508 1708 3520
rect 1291 3480 1708 3508
rect 1291 3477 1303 3480
rect 1245 3471 1303 3477
rect 1702 3468 1708 3480
rect 1760 3508 1766 3520
rect 1797 3511 1855 3517
rect 1797 3508 1809 3511
rect 1760 3480 1809 3508
rect 1760 3468 1766 3480
rect 1797 3477 1809 3480
rect 1843 3477 1855 3511
rect 1797 3471 1855 3477
rect 1334 3332 1340 3384
rect 1392 3372 1398 3384
rect 1429 3375 1487 3381
rect 1429 3372 1441 3375
rect 1392 3344 1441 3372
rect 1392 3332 1398 3344
rect 1429 3341 1441 3344
rect 1475 3372 1487 3375
rect 1904 3372 1932 3548
rect 3174 3536 3180 3548
rect 3232 3536 3238 3588
rect 2346 3400 2352 3452
rect 2404 3440 2410 3452
rect 2533 3443 2591 3449
rect 2533 3440 2545 3443
rect 2404 3412 2545 3440
rect 2404 3400 2410 3412
rect 2533 3409 2545 3412
rect 2579 3409 2591 3443
rect 2533 3403 2591 3409
rect 1475 3344 1932 3372
rect 1475 3341 1487 3344
rect 1429 3335 1487 3341
rect 1886 3264 1892 3316
rect 1944 3304 1950 3316
rect 2165 3307 2223 3313
rect 2165 3304 2177 3307
rect 1944 3276 2177 3304
rect 1944 3264 1950 3276
rect 2165 3273 2177 3276
rect 2211 3304 2223 3307
rect 2349 3307 2407 3313
rect 2349 3304 2361 3307
rect 2211 3276 2361 3304
rect 2211 3273 2223 3276
rect 2165 3267 2223 3273
rect 2349 3273 2361 3276
rect 2395 3273 2407 3307
rect 2349 3267 2407 3273
rect 598 3196 604 3248
rect 656 3236 662 3248
rect 877 3239 935 3245
rect 877 3236 889 3239
rect 656 3208 889 3236
rect 656 3196 662 3208
rect 877 3205 889 3208
rect 923 3205 935 3239
rect 877 3199 935 3205
rect 2073 3239 2131 3245
rect 2073 3205 2085 3239
rect 2119 3236 2131 3239
rect 2438 3236 2444 3248
rect 2119 3208 2444 3236
rect 2119 3205 2131 3208
rect 2073 3199 2131 3205
rect 2438 3196 2444 3208
rect 2496 3196 2502 3248
rect 400 3146 4080 3168
rect 400 3094 2546 3146
rect 2598 3094 2610 3146
rect 2662 3094 2674 3146
rect 2726 3094 2738 3146
rect 2790 3094 2802 3146
rect 2854 3094 4080 3146
rect 400 3072 4080 3094
rect 1426 2924 1432 2976
rect 1484 2964 1490 2976
rect 1484 2936 2300 2964
rect 1484 2924 1490 2936
rect 2272 2908 2300 2936
rect 874 2856 880 2908
rect 932 2896 938 2908
rect 1334 2896 1340 2908
rect 932 2868 1340 2896
rect 932 2856 938 2868
rect 1334 2856 1340 2868
rect 1392 2856 1398 2908
rect 1702 2896 1708 2908
rect 1663 2868 1708 2896
rect 1702 2856 1708 2868
rect 1760 2856 1766 2908
rect 2254 2896 2260 2908
rect 2167 2868 2260 2896
rect 2254 2856 2260 2868
rect 2312 2856 2318 2908
rect 2438 2856 2444 2908
rect 2496 2896 2502 2908
rect 2809 2899 2867 2905
rect 2809 2896 2821 2899
rect 2496 2868 2821 2896
rect 2496 2856 2502 2868
rect 2809 2865 2821 2868
rect 2855 2896 2867 2899
rect 3174 2896 3180 2908
rect 2855 2868 3180 2896
rect 2855 2865 2867 2868
rect 2809 2859 2867 2865
rect 3174 2856 3180 2868
rect 3232 2856 3238 2908
rect 782 2828 788 2840
rect 743 2800 788 2828
rect 782 2788 788 2800
rect 840 2788 846 2840
rect 1150 2828 1156 2840
rect 1111 2800 1156 2828
rect 1150 2788 1156 2800
rect 1208 2788 1214 2840
rect 1610 2828 1616 2840
rect 1571 2800 1616 2828
rect 1610 2788 1616 2800
rect 1668 2788 1674 2840
rect 2993 2831 3051 2837
rect 2993 2797 3005 2831
rect 3039 2828 3051 2831
rect 3082 2828 3088 2840
rect 3039 2800 3088 2828
rect 3039 2797 3051 2800
rect 2993 2791 3051 2797
rect 3082 2788 3088 2800
rect 3140 2828 3146 2840
rect 4094 2828 4100 2840
rect 3140 2800 4100 2828
rect 3140 2788 3146 2800
rect 4094 2788 4100 2800
rect 4152 2788 4158 2840
rect 2070 2692 2076 2704
rect 2031 2664 2076 2692
rect 2070 2652 2076 2664
rect 2128 2652 2134 2704
rect 3174 2692 3180 2704
rect 3135 2664 3180 2692
rect 3174 2652 3180 2664
rect 3232 2652 3238 2704
rect 400 2602 4080 2624
rect 400 2550 1046 2602
rect 1098 2550 1110 2602
rect 1162 2550 1174 2602
rect 1226 2550 1238 2602
rect 1290 2550 1302 2602
rect 1354 2550 4080 2602
rect 400 2528 4080 2550
rect 785 2491 843 2497
rect 785 2457 797 2491
rect 831 2488 843 2491
rect 874 2488 880 2500
rect 831 2460 880 2488
rect 831 2457 843 2460
rect 785 2451 843 2457
rect 874 2448 880 2460
rect 932 2448 938 2500
rect 2254 2448 2260 2500
rect 2312 2488 2318 2500
rect 2901 2491 2959 2497
rect 2901 2488 2913 2491
rect 2312 2460 2913 2488
rect 2312 2448 2318 2460
rect 2901 2457 2913 2460
rect 2947 2457 2959 2491
rect 3082 2488 3088 2500
rect 3043 2460 3088 2488
rect 2901 2451 2959 2457
rect 3082 2448 3088 2460
rect 3140 2448 3146 2500
rect 966 2380 972 2432
rect 1024 2420 1030 2432
rect 1061 2423 1119 2429
rect 1061 2420 1073 2423
rect 1024 2392 1073 2420
rect 1024 2380 1030 2392
rect 1061 2389 1073 2392
rect 1107 2389 1119 2423
rect 1061 2383 1119 2389
rect 2070 2352 2076 2364
rect 1812 2324 2076 2352
rect 414 2176 420 2228
rect 472 2216 478 2228
rect 877 2219 935 2225
rect 877 2216 889 2219
rect 472 2188 889 2216
rect 472 2176 478 2188
rect 877 2185 889 2188
rect 923 2216 935 2219
rect 1610 2216 1616 2228
rect 923 2188 1616 2216
rect 923 2185 935 2188
rect 877 2179 935 2185
rect 1610 2176 1616 2188
rect 1668 2176 1674 2228
rect 782 2108 788 2160
rect 840 2148 846 2160
rect 1245 2151 1303 2157
rect 1245 2148 1257 2151
rect 840 2120 1257 2148
rect 840 2108 846 2120
rect 1245 2117 1257 2120
rect 1291 2148 1303 2151
rect 1429 2151 1487 2157
rect 1429 2148 1441 2151
rect 1291 2120 1441 2148
rect 1291 2117 1303 2120
rect 1245 2111 1303 2117
rect 1429 2117 1441 2120
rect 1475 2117 1487 2151
rect 1429 2111 1487 2117
rect 1518 2108 1524 2160
rect 1576 2148 1582 2160
rect 1812 2157 1840 2324
rect 2070 2312 2076 2324
rect 2128 2352 2134 2364
rect 2990 2352 2996 2364
rect 2128 2324 2996 2352
rect 2128 2312 2134 2324
rect 2364 2293 2392 2324
rect 2990 2312 2996 2324
rect 3048 2352 3054 2364
rect 3269 2355 3327 2361
rect 3269 2352 3281 2355
rect 3048 2324 3281 2352
rect 3048 2312 3054 2324
rect 3269 2321 3281 2324
rect 3315 2321 3327 2355
rect 3269 2315 3327 2321
rect 1981 2287 2039 2293
rect 1981 2253 1993 2287
rect 2027 2284 2039 2287
rect 2349 2287 2407 2293
rect 2027 2256 2300 2284
rect 2027 2253 2039 2256
rect 1981 2247 2039 2253
rect 2272 2160 2300 2256
rect 2349 2253 2361 2287
rect 2395 2253 2407 2287
rect 2349 2247 2407 2253
rect 2625 2287 2683 2293
rect 2625 2253 2637 2287
rect 2671 2284 2683 2287
rect 2898 2284 2904 2296
rect 2671 2256 2904 2284
rect 2671 2253 2683 2256
rect 2625 2247 2683 2253
rect 2898 2244 2904 2256
rect 2956 2284 2962 2296
rect 3453 2287 3511 2293
rect 3453 2284 3465 2287
rect 2956 2256 3465 2284
rect 2956 2244 2962 2256
rect 3453 2253 3465 2256
rect 3499 2253 3511 2287
rect 3453 2247 3511 2253
rect 1797 2151 1855 2157
rect 1797 2148 1809 2151
rect 1576 2120 1809 2148
rect 1576 2108 1582 2120
rect 1797 2117 1809 2120
rect 1843 2117 1855 2151
rect 2254 2148 2260 2160
rect 2215 2120 2260 2148
rect 1797 2111 1855 2117
rect 2254 2108 2260 2120
rect 2312 2108 2318 2160
rect 2346 2108 2352 2160
rect 2404 2148 2410 2160
rect 3637 2151 3695 2157
rect 3637 2148 3649 2151
rect 2404 2120 3649 2148
rect 2404 2108 2410 2120
rect 3637 2117 3649 2120
rect 3683 2117 3695 2151
rect 3637 2111 3695 2117
rect 400 2058 4080 2080
rect 400 2006 2546 2058
rect 2598 2006 2610 2058
rect 2662 2006 2674 2058
rect 2726 2006 2738 2058
rect 2790 2006 2802 2058
rect 2854 2006 4080 2058
rect 400 1984 4080 2006
rect 2990 1944 2996 1956
rect 2951 1916 2996 1944
rect 2990 1904 2996 1916
rect 3048 1944 3054 1956
rect 3085 1947 3143 1953
rect 3085 1944 3097 1947
rect 3048 1916 3097 1944
rect 3048 1904 3054 1916
rect 3085 1913 3097 1916
rect 3131 1913 3143 1947
rect 3085 1907 3143 1913
rect 1426 1836 1432 1888
rect 1484 1836 1490 1888
rect 693 1811 751 1817
rect 693 1777 705 1811
rect 739 1808 751 1811
rect 782 1808 788 1820
rect 739 1780 788 1808
rect 739 1777 751 1780
rect 693 1771 751 1777
rect 782 1768 788 1780
rect 840 1768 846 1820
rect 598 1700 604 1752
rect 656 1740 662 1752
rect 1061 1743 1119 1749
rect 1061 1740 1073 1743
rect 656 1712 1073 1740
rect 656 1700 662 1712
rect 708 1604 736 1712
rect 1061 1709 1073 1712
rect 1107 1709 1119 1743
rect 1061 1703 1119 1709
rect 1610 1700 1616 1752
rect 1668 1740 1674 1752
rect 2346 1740 2352 1752
rect 1668 1712 2352 1740
rect 1668 1700 1674 1712
rect 2346 1700 2352 1712
rect 2404 1740 2410 1752
rect 2441 1743 2499 1749
rect 2441 1740 2453 1743
rect 2404 1712 2453 1740
rect 2404 1700 2410 1712
rect 2441 1709 2453 1712
rect 2487 1709 2499 1743
rect 2441 1703 2499 1709
rect 2806 1632 2812 1684
rect 2864 1672 2870 1684
rect 3361 1675 3419 1681
rect 3361 1672 3373 1675
rect 2864 1644 3373 1672
rect 2864 1632 2870 1644
rect 3361 1641 3373 1644
rect 3407 1641 3419 1675
rect 3361 1635 3419 1641
rect 3542 1604 3548 1616
rect 708 1576 3548 1604
rect 3542 1564 3548 1576
rect 3600 1564 3606 1616
rect 400 1514 4080 1536
rect 400 1462 1046 1514
rect 1098 1462 1110 1514
rect 1162 1462 1174 1514
rect 1226 1462 1238 1514
rect 1290 1462 1302 1514
rect 1354 1462 4080 1514
rect 400 1440 4080 1462
rect 3174 1264 3180 1276
rect 3135 1236 3180 1264
rect 3174 1224 3180 1236
rect 3232 1224 3238 1276
rect 693 1199 751 1205
rect 693 1165 705 1199
rect 739 1196 751 1199
rect 1334 1196 1340 1208
rect 739 1168 1340 1196
rect 739 1165 751 1168
rect 693 1159 751 1165
rect 1334 1156 1340 1168
rect 1392 1156 1398 1208
rect 1429 1199 1487 1205
rect 1429 1165 1441 1199
rect 1475 1196 1487 1199
rect 1702 1196 1708 1208
rect 1475 1168 1708 1196
rect 1475 1165 1487 1168
rect 1429 1159 1487 1165
rect 1702 1156 1708 1168
rect 1760 1156 1766 1208
rect 1797 1199 1855 1205
rect 1797 1165 1809 1199
rect 1843 1196 1855 1199
rect 1886 1196 1892 1208
rect 1843 1168 1892 1196
rect 1843 1165 1855 1168
rect 1797 1159 1855 1165
rect 1886 1156 1892 1168
rect 1944 1156 1950 1208
rect 969 1131 1027 1137
rect 969 1097 981 1131
rect 1015 1128 1027 1131
rect 1518 1128 1524 1140
rect 1015 1100 1524 1128
rect 1015 1097 1027 1100
rect 969 1091 1027 1097
rect 1518 1088 1524 1100
rect 1576 1088 1582 1140
rect 2806 1088 2812 1140
rect 2864 1088 2870 1140
rect 782 1020 788 1072
rect 840 1060 846 1072
rect 1337 1063 1395 1069
rect 1337 1060 1349 1063
rect 840 1032 1349 1060
rect 840 1020 846 1032
rect 1337 1029 1349 1032
rect 1383 1060 1395 1063
rect 1702 1060 1708 1072
rect 1383 1032 1708 1060
rect 1383 1029 1395 1032
rect 1337 1023 1395 1029
rect 1702 1020 1708 1032
rect 1760 1060 1766 1072
rect 3082 1060 3088 1072
rect 1760 1032 3088 1060
rect 1760 1020 1766 1032
rect 3082 1020 3088 1032
rect 3140 1020 3146 1072
rect 3634 1020 3640 1072
rect 3692 1060 3698 1072
rect 3692 1032 3737 1060
rect 3692 1020 3698 1032
rect 400 970 4080 992
rect 400 918 2546 970
rect 2598 918 2610 970
rect 2662 918 2674 970
rect 2726 918 2738 970
rect 2790 918 2802 970
rect 2854 918 4080 970
rect 400 896 4080 918
rect 3634 856 3640 868
rect 1536 828 3640 856
rect 1536 800 1564 828
rect 3634 816 3640 828
rect 3692 816 3698 868
rect 1518 748 1524 800
rect 1576 748 1582 800
rect 782 720 788 732
rect 743 692 788 720
rect 782 680 788 692
rect 840 680 846 732
rect 3542 720 3548 732
rect 3503 692 3548 720
rect 3542 680 3548 692
rect 3600 680 3606 732
rect 1153 655 1211 661
rect 1153 621 1165 655
rect 1199 652 1211 655
rect 1610 652 1616 664
rect 1199 624 1616 652
rect 1199 621 1211 624
rect 1153 615 1211 621
rect 1610 612 1616 624
rect 1668 612 1674 664
rect 1886 612 1892 664
rect 1944 652 1950 664
rect 2533 655 2591 661
rect 2533 652 2545 655
rect 1944 624 2545 652
rect 1944 612 1950 624
rect 2533 621 2545 624
rect 2579 621 2591 655
rect 2533 615 2591 621
rect 3082 584 3088 596
rect 2995 556 3088 584
rect 3082 544 3088 556
rect 3140 584 3146 596
rect 4094 584 4100 596
rect 3140 556 4100 584
rect 3140 544 3146 556
rect 4094 544 4100 556
rect 4152 544 4158 596
rect 400 426 4080 448
rect 400 374 1046 426
rect 1098 374 1110 426
rect 1162 374 1174 426
rect 1226 374 1238 426
rect 1290 374 1302 426
rect 1354 374 4080 426
rect 400 352 4080 374
<< via1 >>
rect 1046 3638 1098 3690
rect 1110 3638 1162 3690
rect 1174 3638 1226 3690
rect 1238 3638 1290 3690
rect 1302 3638 1354 3690
rect 1708 3468 1760 3520
rect 1340 3332 1392 3384
rect 3180 3536 3232 3588
rect 2352 3400 2404 3452
rect 1892 3264 1944 3316
rect 604 3196 656 3248
rect 2444 3196 2496 3248
rect 2546 3094 2598 3146
rect 2610 3094 2662 3146
rect 2674 3094 2726 3146
rect 2738 3094 2790 3146
rect 2802 3094 2854 3146
rect 1432 2924 1484 2976
rect 880 2856 932 2908
rect 1340 2899 1392 2908
rect 1340 2865 1349 2899
rect 1349 2865 1383 2899
rect 1383 2865 1392 2899
rect 1340 2856 1392 2865
rect 1708 2899 1760 2908
rect 1708 2865 1717 2899
rect 1717 2865 1751 2899
rect 1751 2865 1760 2899
rect 1708 2856 1760 2865
rect 2260 2899 2312 2908
rect 2260 2865 2269 2899
rect 2269 2865 2303 2899
rect 2303 2865 2312 2899
rect 2260 2856 2312 2865
rect 2444 2856 2496 2908
rect 3180 2856 3232 2908
rect 788 2831 840 2840
rect 788 2797 797 2831
rect 797 2797 831 2831
rect 831 2797 840 2831
rect 788 2788 840 2797
rect 1156 2831 1208 2840
rect 1156 2797 1165 2831
rect 1165 2797 1199 2831
rect 1199 2797 1208 2831
rect 1156 2788 1208 2797
rect 1616 2831 1668 2840
rect 1616 2797 1625 2831
rect 1625 2797 1659 2831
rect 1659 2797 1668 2831
rect 1616 2788 1668 2797
rect 3088 2788 3140 2840
rect 4100 2788 4152 2840
rect 2076 2695 2128 2704
rect 2076 2661 2085 2695
rect 2085 2661 2119 2695
rect 2119 2661 2128 2695
rect 2076 2652 2128 2661
rect 3180 2695 3232 2704
rect 3180 2661 3189 2695
rect 3189 2661 3223 2695
rect 3223 2661 3232 2695
rect 3180 2652 3232 2661
rect 1046 2550 1098 2602
rect 1110 2550 1162 2602
rect 1174 2550 1226 2602
rect 1238 2550 1290 2602
rect 1302 2550 1354 2602
rect 880 2448 932 2500
rect 2260 2448 2312 2500
rect 3088 2491 3140 2500
rect 3088 2457 3097 2491
rect 3097 2457 3131 2491
rect 3131 2457 3140 2491
rect 3088 2448 3140 2457
rect 972 2380 1024 2432
rect 420 2176 472 2228
rect 1616 2176 1668 2228
rect 788 2108 840 2160
rect 1524 2108 1576 2160
rect 2076 2312 2128 2364
rect 2996 2312 3048 2364
rect 2904 2244 2956 2296
rect 2260 2151 2312 2160
rect 2260 2117 2269 2151
rect 2269 2117 2303 2151
rect 2303 2117 2312 2151
rect 2260 2108 2312 2117
rect 2352 2108 2404 2160
rect 2546 2006 2598 2058
rect 2610 2006 2662 2058
rect 2674 2006 2726 2058
rect 2738 2006 2790 2058
rect 2802 2006 2854 2058
rect 2996 1947 3048 1956
rect 2996 1913 3005 1947
rect 3005 1913 3039 1947
rect 3039 1913 3048 1947
rect 2996 1904 3048 1913
rect 1432 1836 1484 1888
rect 788 1768 840 1820
rect 604 1700 656 1752
rect 1616 1700 1668 1752
rect 2352 1700 2404 1752
rect 2812 1632 2864 1684
rect 3548 1607 3600 1616
rect 3548 1573 3557 1607
rect 3557 1573 3591 1607
rect 3591 1573 3600 1607
rect 3548 1564 3600 1573
rect 1046 1462 1098 1514
rect 1110 1462 1162 1514
rect 1174 1462 1226 1514
rect 1238 1462 1290 1514
rect 1302 1462 1354 1514
rect 3180 1267 3232 1276
rect 3180 1233 3189 1267
rect 3189 1233 3223 1267
rect 3223 1233 3232 1267
rect 3180 1224 3232 1233
rect 1340 1156 1392 1208
rect 1708 1156 1760 1208
rect 1892 1156 1944 1208
rect 1524 1088 1576 1140
rect 2812 1088 2864 1140
rect 788 1020 840 1072
rect 1708 1020 1760 1072
rect 3088 1020 3140 1072
rect 3640 1063 3692 1072
rect 3640 1029 3649 1063
rect 3649 1029 3683 1063
rect 3683 1029 3692 1063
rect 3640 1020 3692 1029
rect 2546 918 2598 970
rect 2610 918 2662 970
rect 2674 918 2726 970
rect 2738 918 2790 970
rect 2802 918 2854 970
rect 3640 859 3692 868
rect 3640 825 3649 859
rect 3649 825 3683 859
rect 3683 825 3692 859
rect 3640 816 3692 825
rect 1524 748 1576 800
rect 788 723 840 732
rect 788 689 797 723
rect 797 689 831 723
rect 831 689 840 723
rect 788 680 840 689
rect 3548 723 3600 732
rect 3548 689 3557 723
rect 3557 689 3591 723
rect 3591 689 3600 723
rect 3548 680 3600 689
rect 1616 612 1668 664
rect 1892 612 1944 664
rect 3088 587 3140 596
rect 3088 553 3097 587
rect 3097 553 3131 587
rect 3131 553 3140 587
rect 3088 544 3140 553
rect 4100 544 4152 596
rect 1046 374 1098 426
rect 1110 374 1162 426
rect 1174 374 1226 426
rect 1238 374 1290 426
rect 1302 374 1354 426
<< metal2 >>
rect 1310 4119 1422 4543
rect 3150 4119 3262 4543
rect 1352 3882 1380 4119
rect 1352 3854 1472 3882
rect 1040 3692 1360 3712
rect 1040 3690 1052 3692
rect 1108 3690 1132 3692
rect 1188 3690 1212 3692
rect 1268 3690 1292 3692
rect 1348 3690 1360 3692
rect 1040 3638 1046 3690
rect 1108 3638 1110 3690
rect 1290 3638 1292 3690
rect 1354 3638 1360 3690
rect 1040 3636 1052 3638
rect 1108 3636 1132 3638
rect 1188 3636 1212 3638
rect 1268 3636 1292 3638
rect 1348 3636 1360 3638
rect 1040 3616 1360 3636
rect 1340 3384 1392 3390
rect 1340 3326 1392 3332
rect 604 3248 656 3254
rect 604 3190 656 3196
rect 420 2228 472 2234
rect 420 2170 472 2176
rect 432 424 460 2170
rect 616 1758 644 3190
rect 1154 2944 1210 2953
rect 880 2908 932 2914
rect 1352 2914 1380 3326
rect 1444 2982 1472 3854
rect 3192 3594 3220 4119
rect 3180 3588 3232 3594
rect 3180 3530 3232 3536
rect 1708 3520 1760 3526
rect 1708 3462 1760 3468
rect 1432 2976 1484 2982
rect 1432 2918 1484 2924
rect 1720 2914 1748 3462
rect 2352 3452 2404 3458
rect 2352 3394 2404 3400
rect 1892 3316 1944 3322
rect 1892 3258 1944 3264
rect 1154 2879 1210 2888
rect 1340 2908 1392 2914
rect 880 2850 932 2856
rect 788 2840 840 2846
rect 788 2782 840 2788
rect 800 2166 828 2782
rect 892 2506 920 2850
rect 1168 2846 1196 2879
rect 1340 2850 1392 2856
rect 1708 2908 1760 2914
rect 1708 2850 1760 2856
rect 1156 2840 1208 2846
rect 984 2800 1156 2828
rect 880 2500 932 2506
rect 880 2442 932 2448
rect 984 2438 1012 2800
rect 1156 2782 1208 2788
rect 1616 2840 1668 2846
rect 1616 2782 1668 2788
rect 1040 2604 1360 2624
rect 1040 2602 1052 2604
rect 1108 2602 1132 2604
rect 1188 2602 1212 2604
rect 1268 2602 1292 2604
rect 1348 2602 1360 2604
rect 1040 2550 1046 2602
rect 1108 2550 1110 2602
rect 1290 2550 1292 2602
rect 1354 2550 1360 2602
rect 1040 2548 1052 2550
rect 1108 2548 1132 2550
rect 1188 2548 1212 2550
rect 1268 2548 1292 2550
rect 1348 2548 1360 2550
rect 1040 2528 1360 2548
rect 972 2432 1024 2438
rect 972 2374 1024 2380
rect 1628 2234 1656 2782
rect 1616 2228 1668 2234
rect 1616 2170 1668 2176
rect 788 2160 840 2166
rect 1524 2160 1576 2166
rect 788 2102 840 2108
rect 1444 2120 1524 2148
rect 800 1826 828 2102
rect 1444 1894 1472 2120
rect 1524 2102 1576 2108
rect 1432 1888 1484 1894
rect 1432 1830 1484 1836
rect 788 1820 840 1826
rect 788 1762 840 1768
rect 604 1752 656 1758
rect 604 1694 656 1700
rect 800 1078 828 1762
rect 1040 1516 1360 1536
rect 1040 1514 1052 1516
rect 1108 1514 1132 1516
rect 1188 1514 1212 1516
rect 1268 1514 1292 1516
rect 1348 1514 1360 1516
rect 1040 1462 1046 1514
rect 1108 1462 1110 1514
rect 1290 1462 1292 1514
rect 1354 1462 1360 1514
rect 1040 1460 1052 1462
rect 1108 1460 1132 1462
rect 1188 1460 1212 1462
rect 1268 1460 1292 1462
rect 1348 1460 1360 1462
rect 1040 1440 1360 1460
rect 1340 1208 1392 1214
rect 1444 1196 1472 1830
rect 1616 1752 1668 1758
rect 1616 1694 1668 1700
rect 1392 1168 1472 1196
rect 1340 1150 1392 1156
rect 1524 1140 1576 1146
rect 1524 1082 1576 1088
rect 788 1072 840 1078
rect 788 1014 840 1020
rect 800 738 828 1014
rect 1536 806 1564 1082
rect 1524 800 1576 806
rect 1524 742 1576 748
rect 788 732 840 738
rect 788 674 840 680
rect 1628 670 1656 1694
rect 1904 1214 1932 3258
rect 2260 2908 2312 2914
rect 2260 2850 2312 2856
rect 2076 2704 2128 2710
rect 2076 2646 2128 2652
rect 2088 2370 2116 2646
rect 2272 2506 2300 2850
rect 2260 2500 2312 2506
rect 2260 2442 2312 2448
rect 2076 2364 2128 2370
rect 2076 2306 2128 2312
rect 2364 2166 2392 3394
rect 2444 3248 2496 3254
rect 2444 3190 2496 3196
rect 2456 2914 2484 3190
rect 2540 3148 2860 3168
rect 2540 3146 2552 3148
rect 2608 3146 2632 3148
rect 2688 3146 2712 3148
rect 2768 3146 2792 3148
rect 2848 3146 2860 3148
rect 2540 3094 2546 3146
rect 2608 3094 2610 3146
rect 2790 3094 2792 3146
rect 2854 3094 2860 3146
rect 2540 3092 2552 3094
rect 2608 3092 2632 3094
rect 2688 3092 2712 3094
rect 2768 3092 2792 3094
rect 2848 3092 2860 3094
rect 2540 3072 2860 3092
rect 4098 2944 4154 2953
rect 2444 2908 2496 2914
rect 2444 2850 2496 2856
rect 3180 2908 3232 2914
rect 4098 2879 4154 2888
rect 3180 2850 3232 2856
rect 3088 2840 3140 2846
rect 3088 2782 3140 2788
rect 3100 2506 3128 2782
rect 3192 2710 3220 2850
rect 4112 2846 4140 2879
rect 4100 2840 4152 2846
rect 4100 2782 4152 2788
rect 3180 2704 3232 2710
rect 3180 2646 3232 2652
rect 3088 2500 3140 2506
rect 3088 2442 3140 2448
rect 2996 2364 3048 2370
rect 2996 2306 3048 2312
rect 2904 2296 2956 2302
rect 2904 2238 2956 2244
rect 2260 2160 2312 2166
rect 2260 2102 2312 2108
rect 2352 2160 2404 2166
rect 2352 2102 2404 2108
rect 1708 1208 1760 1214
rect 1708 1150 1760 1156
rect 1892 1208 1944 1214
rect 1892 1150 1944 1156
rect 1720 1078 1748 1150
rect 1708 1072 1760 1078
rect 1708 1014 1760 1020
rect 1904 670 1932 1150
rect 1616 664 1668 670
rect 1616 606 1668 612
rect 1892 664 1944 670
rect 1892 606 1944 612
rect 1040 428 1360 448
rect 1040 426 1052 428
rect 1108 426 1132 428
rect 1188 426 1212 428
rect 1268 426 1292 428
rect 1348 426 1360 428
rect 390 0 502 424
rect 1040 374 1046 426
rect 1108 374 1110 426
rect 1290 374 1292 426
rect 1354 374 1360 426
rect 2272 424 2300 2102
rect 2364 1758 2392 2102
rect 2540 2060 2860 2080
rect 2540 2058 2552 2060
rect 2608 2058 2632 2060
rect 2688 2058 2712 2060
rect 2768 2058 2792 2060
rect 2848 2058 2860 2060
rect 2540 2006 2546 2058
rect 2608 2006 2610 2058
rect 2790 2006 2792 2058
rect 2854 2006 2860 2058
rect 2540 2004 2552 2006
rect 2608 2004 2632 2006
rect 2688 2004 2712 2006
rect 2768 2004 2792 2006
rect 2848 2004 2860 2006
rect 2540 1984 2860 2004
rect 2352 1752 2404 1758
rect 2352 1694 2404 1700
rect 2812 1684 2864 1690
rect 2916 1672 2944 2238
rect 3008 1962 3036 2306
rect 2996 1956 3048 1962
rect 2996 1898 3048 1904
rect 2864 1644 2944 1672
rect 2812 1626 2864 1632
rect 2824 1146 2852 1626
rect 3192 1282 3220 2646
rect 3548 1616 3600 1622
rect 3548 1558 3600 1564
rect 3180 1276 3232 1282
rect 3180 1218 3232 1224
rect 2812 1140 2864 1146
rect 2812 1082 2864 1088
rect 3088 1072 3140 1078
rect 3088 1014 3140 1020
rect 2540 972 2860 992
rect 2540 970 2552 972
rect 2608 970 2632 972
rect 2688 970 2712 972
rect 2768 970 2792 972
rect 2848 970 2860 972
rect 2540 918 2546 970
rect 2608 918 2610 970
rect 2790 918 2792 970
rect 2854 918 2860 970
rect 2540 916 2552 918
rect 2608 916 2632 918
rect 2688 916 2712 918
rect 2768 916 2792 918
rect 2848 916 2860 918
rect 2540 896 2860 916
rect 3100 602 3128 1014
rect 3560 738 3588 1558
rect 3640 1072 3692 1078
rect 3640 1014 3692 1020
rect 3652 874 3680 1014
rect 3640 868 3692 874
rect 3640 810 3692 816
rect 3548 732 3600 738
rect 3548 674 3600 680
rect 3088 596 3140 602
rect 3088 538 3140 544
rect 4100 596 4152 602
rect 4100 538 4152 544
rect 4112 424 4140 538
rect 1040 372 1052 374
rect 1108 372 1132 374
rect 1188 372 1212 374
rect 1268 372 1292 374
rect 1348 372 1360 374
rect 1040 352 1360 372
rect 2230 0 2342 424
rect 4070 0 4182 424
<< via2 >>
rect 1052 3690 1108 3692
rect 1132 3690 1188 3692
rect 1212 3690 1268 3692
rect 1292 3690 1348 3692
rect 1052 3638 1098 3690
rect 1098 3638 1108 3690
rect 1132 3638 1162 3690
rect 1162 3638 1174 3690
rect 1174 3638 1188 3690
rect 1212 3638 1226 3690
rect 1226 3638 1238 3690
rect 1238 3638 1268 3690
rect 1292 3638 1302 3690
rect 1302 3638 1348 3690
rect 1052 3636 1108 3638
rect 1132 3636 1188 3638
rect 1212 3636 1268 3638
rect 1292 3636 1348 3638
rect 1154 2888 1210 2944
rect 1052 2602 1108 2604
rect 1132 2602 1188 2604
rect 1212 2602 1268 2604
rect 1292 2602 1348 2604
rect 1052 2550 1098 2602
rect 1098 2550 1108 2602
rect 1132 2550 1162 2602
rect 1162 2550 1174 2602
rect 1174 2550 1188 2602
rect 1212 2550 1226 2602
rect 1226 2550 1238 2602
rect 1238 2550 1268 2602
rect 1292 2550 1302 2602
rect 1302 2550 1348 2602
rect 1052 2548 1108 2550
rect 1132 2548 1188 2550
rect 1212 2548 1268 2550
rect 1292 2548 1348 2550
rect 1052 1514 1108 1516
rect 1132 1514 1188 1516
rect 1212 1514 1268 1516
rect 1292 1514 1348 1516
rect 1052 1462 1098 1514
rect 1098 1462 1108 1514
rect 1132 1462 1162 1514
rect 1162 1462 1174 1514
rect 1174 1462 1188 1514
rect 1212 1462 1226 1514
rect 1226 1462 1238 1514
rect 1238 1462 1268 1514
rect 1292 1462 1302 1514
rect 1302 1462 1348 1514
rect 1052 1460 1108 1462
rect 1132 1460 1188 1462
rect 1212 1460 1268 1462
rect 1292 1460 1348 1462
rect 2552 3146 2608 3148
rect 2632 3146 2688 3148
rect 2712 3146 2768 3148
rect 2792 3146 2848 3148
rect 2552 3094 2598 3146
rect 2598 3094 2608 3146
rect 2632 3094 2662 3146
rect 2662 3094 2674 3146
rect 2674 3094 2688 3146
rect 2712 3094 2726 3146
rect 2726 3094 2738 3146
rect 2738 3094 2768 3146
rect 2792 3094 2802 3146
rect 2802 3094 2848 3146
rect 2552 3092 2608 3094
rect 2632 3092 2688 3094
rect 2712 3092 2768 3094
rect 2792 3092 2848 3094
rect 4098 2888 4154 2944
rect 1052 426 1108 428
rect 1132 426 1188 428
rect 1212 426 1268 428
rect 1292 426 1348 428
rect 1052 374 1098 426
rect 1098 374 1108 426
rect 1132 374 1162 426
rect 1162 374 1174 426
rect 1174 374 1188 426
rect 1212 374 1226 426
rect 1226 374 1238 426
rect 1238 374 1268 426
rect 1292 374 1302 426
rect 1302 374 1348 426
rect 2552 2058 2608 2060
rect 2632 2058 2688 2060
rect 2712 2058 2768 2060
rect 2792 2058 2848 2060
rect 2552 2006 2598 2058
rect 2598 2006 2608 2058
rect 2632 2006 2662 2058
rect 2662 2006 2674 2058
rect 2674 2006 2688 2058
rect 2712 2006 2726 2058
rect 2726 2006 2738 2058
rect 2738 2006 2768 2058
rect 2792 2006 2802 2058
rect 2802 2006 2848 2058
rect 2552 2004 2608 2006
rect 2632 2004 2688 2006
rect 2712 2004 2768 2006
rect 2792 2004 2848 2006
rect 2552 970 2608 972
rect 2632 970 2688 972
rect 2712 970 2768 972
rect 2792 970 2848 972
rect 2552 918 2598 970
rect 2598 918 2608 970
rect 2632 918 2662 970
rect 2662 918 2674 970
rect 2674 918 2688 970
rect 2712 918 2726 970
rect 2726 918 2738 970
rect 2738 918 2768 970
rect 2792 918 2802 970
rect 2802 918 2848 970
rect 2552 916 2608 918
rect 2632 916 2688 918
rect 2712 916 2768 918
rect 2792 916 2848 918
rect 1052 372 1108 374
rect 1132 372 1188 374
rect 1212 372 1268 374
rect 1292 372 1348 374
<< metal3 >>
rect 1040 3696 1360 3712
rect 1040 3632 1048 3696
rect 1112 3632 1128 3696
rect 1192 3632 1208 3696
rect 1272 3632 1288 3696
rect 1352 3632 1360 3696
rect 1040 3616 1360 3632
rect 2540 3152 2860 3168
rect 2540 3088 2548 3152
rect 2612 3088 2628 3152
rect 2692 3088 2708 3152
rect 2772 3088 2788 3152
rect 2852 3088 2860 3152
rect 2540 3072 2860 3088
rect 0 2946 440 3036
rect 4103 2949 4543 3036
rect 1149 2946 1215 2949
rect 0 2944 1215 2946
rect 0 2888 1154 2944
rect 1210 2888 1215 2944
rect 0 2886 1215 2888
rect 0 2796 440 2886
rect 1149 2883 1215 2886
rect 4093 2944 4543 2949
rect 4093 2888 4098 2944
rect 4154 2888 4543 2944
rect 4093 2883 4543 2888
rect 4103 2796 4543 2883
rect 1040 2608 1360 2624
rect 1040 2544 1048 2608
rect 1112 2544 1128 2608
rect 1192 2544 1208 2608
rect 1272 2544 1288 2608
rect 1352 2544 1360 2608
rect 1040 2528 1360 2544
rect 2540 2064 2860 2080
rect 2540 2000 2548 2064
rect 2612 2000 2628 2064
rect 2692 2000 2708 2064
rect 2772 2000 2788 2064
rect 2852 2000 2860 2064
rect 2540 1984 2860 2000
rect 1040 1520 1360 1536
rect 1040 1456 1048 1520
rect 1112 1456 1128 1520
rect 1192 1456 1208 1520
rect 1272 1456 1288 1520
rect 1352 1456 1360 1520
rect 1040 1440 1360 1456
rect 2540 976 2860 992
rect 2540 912 2548 976
rect 2612 912 2628 976
rect 2692 912 2708 976
rect 2772 912 2788 976
rect 2852 912 2860 976
rect 2540 896 2860 912
rect 1040 432 1360 448
rect 1040 368 1048 432
rect 1112 368 1128 432
rect 1192 368 1208 432
rect 1272 368 1288 432
rect 1352 368 1360 432
rect 1040 352 1360 368
<< via3 >>
rect 1048 3692 1112 3696
rect 1048 3636 1052 3692
rect 1052 3636 1108 3692
rect 1108 3636 1112 3692
rect 1048 3632 1112 3636
rect 1128 3692 1192 3696
rect 1128 3636 1132 3692
rect 1132 3636 1188 3692
rect 1188 3636 1192 3692
rect 1128 3632 1192 3636
rect 1208 3692 1272 3696
rect 1208 3636 1212 3692
rect 1212 3636 1268 3692
rect 1268 3636 1272 3692
rect 1208 3632 1272 3636
rect 1288 3692 1352 3696
rect 1288 3636 1292 3692
rect 1292 3636 1348 3692
rect 1348 3636 1352 3692
rect 1288 3632 1352 3636
rect 2548 3148 2612 3152
rect 2548 3092 2552 3148
rect 2552 3092 2608 3148
rect 2608 3092 2612 3148
rect 2548 3088 2612 3092
rect 2628 3148 2692 3152
rect 2628 3092 2632 3148
rect 2632 3092 2688 3148
rect 2688 3092 2692 3148
rect 2628 3088 2692 3092
rect 2708 3148 2772 3152
rect 2708 3092 2712 3148
rect 2712 3092 2768 3148
rect 2768 3092 2772 3148
rect 2708 3088 2772 3092
rect 2788 3148 2852 3152
rect 2788 3092 2792 3148
rect 2792 3092 2848 3148
rect 2848 3092 2852 3148
rect 2788 3088 2852 3092
rect 1048 2604 1112 2608
rect 1048 2548 1052 2604
rect 1052 2548 1108 2604
rect 1108 2548 1112 2604
rect 1048 2544 1112 2548
rect 1128 2604 1192 2608
rect 1128 2548 1132 2604
rect 1132 2548 1188 2604
rect 1188 2548 1192 2604
rect 1128 2544 1192 2548
rect 1208 2604 1272 2608
rect 1208 2548 1212 2604
rect 1212 2548 1268 2604
rect 1268 2548 1272 2604
rect 1208 2544 1272 2548
rect 1288 2604 1352 2608
rect 1288 2548 1292 2604
rect 1292 2548 1348 2604
rect 1348 2548 1352 2604
rect 1288 2544 1352 2548
rect 2548 2060 2612 2064
rect 2548 2004 2552 2060
rect 2552 2004 2608 2060
rect 2608 2004 2612 2060
rect 2548 2000 2612 2004
rect 2628 2060 2692 2064
rect 2628 2004 2632 2060
rect 2632 2004 2688 2060
rect 2688 2004 2692 2060
rect 2628 2000 2692 2004
rect 2708 2060 2772 2064
rect 2708 2004 2712 2060
rect 2712 2004 2768 2060
rect 2768 2004 2772 2060
rect 2708 2000 2772 2004
rect 2788 2060 2852 2064
rect 2788 2004 2792 2060
rect 2792 2004 2848 2060
rect 2848 2004 2852 2060
rect 2788 2000 2852 2004
rect 1048 1516 1112 1520
rect 1048 1460 1052 1516
rect 1052 1460 1108 1516
rect 1108 1460 1112 1516
rect 1048 1456 1112 1460
rect 1128 1516 1192 1520
rect 1128 1460 1132 1516
rect 1132 1460 1188 1516
rect 1188 1460 1192 1516
rect 1128 1456 1192 1460
rect 1208 1516 1272 1520
rect 1208 1460 1212 1516
rect 1212 1460 1268 1516
rect 1268 1460 1272 1516
rect 1208 1456 1272 1460
rect 1288 1516 1352 1520
rect 1288 1460 1292 1516
rect 1292 1460 1348 1516
rect 1348 1460 1352 1516
rect 1288 1456 1352 1460
rect 2548 972 2612 976
rect 2548 916 2552 972
rect 2552 916 2608 972
rect 2608 916 2612 972
rect 2548 912 2612 916
rect 2628 972 2692 976
rect 2628 916 2632 972
rect 2632 916 2688 972
rect 2688 916 2692 972
rect 2628 912 2692 916
rect 2708 972 2772 976
rect 2708 916 2712 972
rect 2712 916 2768 972
rect 2768 916 2772 972
rect 2708 912 2772 916
rect 2788 972 2852 976
rect 2788 916 2792 972
rect 2792 916 2848 972
rect 2848 916 2852 972
rect 2788 912 2852 916
rect 1048 428 1112 432
rect 1048 372 1052 428
rect 1052 372 1108 428
rect 1108 372 1112 428
rect 1048 368 1112 372
rect 1128 428 1192 432
rect 1128 372 1132 428
rect 1132 372 1188 428
rect 1188 372 1192 428
rect 1128 368 1192 372
rect 1208 428 1272 432
rect 1208 372 1212 428
rect 1212 372 1268 428
rect 1268 372 1272 428
rect 1208 368 1272 372
rect 1288 428 1352 432
rect 1288 372 1292 428
rect 1292 372 1348 428
rect 1348 372 1352 428
rect 1288 368 1352 372
<< metal4 >>
rect 1040 3696 1360 3712
rect 1040 3632 1048 3696
rect 1112 3632 1128 3696
rect 1192 3632 1208 3696
rect 1272 3632 1288 3696
rect 1352 3632 1360 3696
rect 1040 2608 1360 3632
rect 1040 2544 1048 2608
rect 1112 2544 1128 2608
rect 1192 2544 1208 2608
rect 1272 2544 1288 2608
rect 1352 2544 1360 2608
rect 1040 1520 1360 2544
rect 1040 1456 1048 1520
rect 1112 1456 1128 1520
rect 1192 1456 1208 1520
rect 1272 1456 1288 1520
rect 1352 1456 1360 1520
rect 1040 1318 1360 1456
rect 1040 1082 1082 1318
rect 1318 1082 1360 1318
rect 1040 432 1360 1082
rect 1040 368 1048 432
rect 1112 368 1128 432
rect 1192 368 1208 432
rect 1272 368 1288 432
rect 1352 368 1360 432
rect 2540 3152 2860 3664
rect 2540 3088 2548 3152
rect 2612 3088 2628 3152
rect 2692 3088 2708 3152
rect 2772 3088 2788 3152
rect 2852 3088 2860 3152
rect 2540 2818 2860 3088
rect 2540 2582 2582 2818
rect 2818 2582 2860 2818
rect 2540 2064 2860 2582
rect 2540 2000 2548 2064
rect 2612 2000 2628 2064
rect 2692 2000 2708 2064
rect 2772 2000 2788 2064
rect 2852 2000 2860 2064
rect 2540 976 2860 2000
rect 2540 912 2548 976
rect 2612 912 2628 976
rect 2692 912 2708 976
rect 2772 912 2788 976
rect 2852 912 2860 976
rect 2540 400 2860 912
rect 1040 352 1360 368
<< via4 >>
rect 1082 1082 1318 1318
rect 2582 2582 2818 2818
<< metal5 >>
rect 400 2818 4080 2860
rect 400 2582 2582 2818
rect 2818 2582 4080 2818
rect 400 2540 4080 2582
rect 400 1318 4080 1360
rect 400 1082 1082 1318
rect 1318 1082 4080 1318
rect 400 1040 4080 1082
use sky130_fd_sc_hd__decap_3  PHY_2 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 400 0 1 944
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1586547711
transform 1 0 400 0 -1 944
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 1228 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL1380x0 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 676 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _10_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 676 0 1 944
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1586547711
transform 1 0 3804 0 1 944
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1586547711
transform 1 0 3804 0 -1 944
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1586547711
transform 1 0 3620 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1586547711
transform 1 0 2976 0 -1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1586547711
transform 1 0 3620 0 -1 944
box 0 -48 184 592
use sky130_fd_sc_hd__conb_1  _11_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 3344 0 -1 944
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_12 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 3252 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL13800x0
timestamp 1586547711
transform 1 0 3160 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__dfstp_4  _12_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 1412 0 1 944
box 0 -48 2208 592
use sky130_fd_sc_hd__dfstp_4  _13_
timestamp 1586547711
transform 1 0 768 0 -1 944
box 0 -48 2208 592
use sky130_fd_sc_hd__dfstp_4  _14_
timestamp 1586547711
transform 1 0 676 0 -1 2032
box 0 -48 2208 592
use sky130_fd_sc_hd__fill_1  FILL16560x5440
timestamp 1586547711
transform 1 0 3712 0 -1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_13
timestamp 1586547711
transform 1 0 3252 0 -1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1586547711
transform 1 0 3528 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1586547711
transform 1 0 3344 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1586547711
transform 1 0 3068 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1586547711
transform 1 0 2884 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1586547711
transform 1 0 3804 0 -1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1586547711
transform 1 0 400 0 -1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1586547711
transform 1 0 400 0 1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1586547711
transform 1 0 676 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1586547711
transform 1 0 860 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1586547711
transform 1 0 1044 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1586547711
transform 1 0 1228 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1586547711
transform 1 0 1412 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL5980x8160
timestamp 1586547711
transform 1 0 1596 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _05_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 1688 0 1 2032
box 0 -48 460 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1586547711
transform 1 0 2148 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _09_
timestamp 1586547711
transform 1 0 2332 0 1 2032
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1586547711
transform 1 0 2884 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1586547711
transform 1 0 3068 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1586547711
transform 1 0 3252 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1586547711
transform 1 0 3436 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1586547711
transform 1 0 3620 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1586547711
transform 1 0 3804 0 1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1586547711
transform 1 0 400 0 -1 3120
box 0 -48 276 592
use sky130_fd_sc_hd__o22a_4  _08_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 676 0 -1 3120
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1586547711
transform 1 0 1964 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL8740x10880
timestamp 1586547711
transform 1 0 2148 0 -1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__nor2_4  _06_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 2240 0 -1 3120
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1586547711
transform 1 0 3804 0 -1 3120
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1586547711
transform 1 0 3068 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_14
timestamp 1586547711
transform 1 0 3252 0 -1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL16560x10880
timestamp 1586547711
transform 1 0 3712 0 -1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL14720x10880 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 3344 0 -1 3120
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1586547711
transform 1 0 400 0 1 3120
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1586547711
transform 1 0 676 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1586547711
transform 1 0 860 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL3220x13600
timestamp 1586547711
transform 1 0 1044 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _07_
timestamp 1586547711
transform 1 0 1136 0 1 3120
box 0 -48 460 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1586547711
transform 1 0 1596 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1586547711
transform 1 0 1780 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1586547711
transform 1 0 1964 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1586547711
transform 1 0 2148 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1586547711
transform 1 0 2332 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1586547711
transform 1 0 2516 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL11500x13600 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 2700 0 1 3120
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_15
timestamp 1586547711
transform 1 0 3252 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL16560x13600
timestamp 1586547711
transform 1 0 3712 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL14720x13600
timestamp 1586547711
transform 1 0 3344 0 1 3120
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1586547711
transform 1 0 3804 0 1 3120
box 0 -48 276 592
<< labels >>
rlabel metal2 s 3150 4119 3262 4543 6 ext_clk_sel
port 0 nsew default input
rlabel metal2 s 390 0 502 424 8 ext_clk
port 1 nsew default input
rlabel metal3 s 0 2796 440 3036 4 pll_clk
port 2 nsew default input
rlabel metal2 s 2230 0 2342 424 8 reset
port 3 nsew default input
rlabel metal2 s 1310 4119 1422 4543 6 ext_reset
port 4 nsew default input
rlabel metal2 s 4070 0 4182 424 8 clk
port 5 nsew default tristate
rlabel metal3 s 4103 2796 4543 3036 6 resetn
port 6 nsew default tristate
flabel metal5 s 3748 1088 4036 1336 0 FreeSans 1600 0 0 0 vdd1v8
port 7 nsew
flabel metal5 s 3720 2578 4008 2826 0 FreeSans 1600 0 0 0 vss
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 4543 4543
<< end >>
