magic
tech sky130A
timestamp 1586445093
<< checkpaint >>
rect 197 197 2545 2553
use s8iom0s8_com_bus_slice_1um  FILLER_5
timestamp 0
transform 1 0 204 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_6
timestamp 0
transform 1 0 205 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_7
timestamp 0
transform 1 0 206 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_8
timestamp 0
transform 1 0 207 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_9
timestamp 0
transform 1 0 208 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_10
timestamp 0
transform 1 0 209 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_11
timestamp 0
transform 1 0 210 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_12
timestamp 0
transform 1 0 211 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_13
timestamp 0
transform 1 0 212 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_14
timestamp 0
transform 1 0 213 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_15
timestamp 0
transform 1 0 214 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_16
timestamp 0
transform 1 0 215 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_17
timestamp 0
transform 1 0 216 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_18
timestamp 0
transform 1 0 217 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_19
timestamp 0
transform 1 0 218 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_20
timestamp 0
transform 1 0 219 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_21
timestamp 0
transform 1 0 220 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_22
timestamp 0
transform 1 0 221 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_23
timestamp 0
transform 1 0 222 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_24
timestamp 0
transform 1 0 223 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_25
timestamp 0
transform 1 0 224 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_26
timestamp 0
transform 1 0 225 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_27
timestamp 0
transform 1 0 226 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_28
timestamp 0
transform 1 0 227 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_29
timestamp 0
transform 1 0 228 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_30
timestamp 0
transform 1 0 229 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_31
timestamp 0
transform 1 0 230 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_32
timestamp 0
transform 1 0 231 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_33
timestamp 0
transform 1 0 232 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_34
timestamp 0
transform 1 0 233 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_35
timestamp 0
transform 1 0 234 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_36
timestamp 0
transform 1 0 235 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_37
timestamp 0
transform 1 0 236 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_38
timestamp 0
transform 1 0 237 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_39
timestamp 0
transform 1 0 238 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_40
timestamp 0
transform 1 0 239 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_41
timestamp 0
transform 1 0 240 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_42
timestamp 0
transform 1 0 241 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_43
timestamp 0
transform 1 0 242 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_44
timestamp 0
transform 1 0 243 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_45
timestamp 0
transform 1 0 244 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_46
timestamp 0
transform 1 0 245 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_47
timestamp 0
transform 1 0 246 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_48
timestamp 0
transform 1 0 247 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_49
timestamp 0
transform 1 0 248 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_50
timestamp 0
transform 1 0 249 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_51
timestamp 0
transform 1 0 250 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_52
timestamp 0
transform 1 0 251 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_53
timestamp 0
transform 1 0 252 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_54
timestamp 0
transform 1 0 253 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_55
timestamp 0
transform 1 0 254 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_56
timestamp 0
transform 1 0 255 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_57
timestamp 0
transform 1 0 256 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_58
timestamp 0
transform 1 0 257 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_59
timestamp 0
transform 1 0 258 0 1 2552
box 0 0 1 1
use s8iom0_vdda_hvc_pad  vdd3v3hclamp[0]
timestamp 0
transform 1 0 259 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_61
timestamp 0
transform 1 0 334 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_62
timestamp 0
transform 1 0 335 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_63
timestamp 0
transform 1 0 336 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_64
timestamp 0
transform 1 0 337 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_65
timestamp 0
transform 1 0 338 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_66
timestamp 0
transform 1 0 339 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_67
timestamp 0
transform 1 0 340 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_68
timestamp 0
transform 1 0 341 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_69
timestamp 0
transform 1 0 342 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_70
timestamp 0
transform 1 0 343 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_71
timestamp 0
transform 1 0 344 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_72
timestamp 0
transform 1 0 345 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_73
timestamp 0
transform 1 0 346 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_74
timestamp 0
transform 1 0 347 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_75
timestamp 0
transform 1 0 348 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_76
timestamp 0
transform 1 0 349 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_77
timestamp 0
transform 1 0 350 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_78
timestamp 0
transform 1 0 351 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_79
timestamp 0
transform 1 0 352 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_80
timestamp 0
transform 1 0 353 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_81
timestamp 0
transform 1 0 354 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_82
timestamp 0
transform 1 0 355 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_83
timestamp 0
transform 1 0 356 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_84
timestamp 0
transform 1 0 357 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_85
timestamp 0
transform 1 0 358 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_86
timestamp 0
transform 1 0 359 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_87
timestamp 0
transform 1 0 360 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_88
timestamp 0
transform 1 0 361 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_89
timestamp 0
transform 1 0 362 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_90
timestamp 0
transform 1 0 363 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_91
timestamp 0
transform 1 0 364 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_92
timestamp 0
transform 1 0 365 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_93
timestamp 0
transform 1 0 366 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_94
timestamp 0
transform 1 0 367 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_95
timestamp 0
transform 1 0 368 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_96
timestamp 0
transform 1 0 369 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_97
timestamp 0
transform 1 0 370 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_98
timestamp 0
transform 1 0 371 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_99
timestamp 0
transform 1 0 372 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_100
timestamp 0
transform 1 0 373 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_101
timestamp 0
transform 1 0 374 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_102
timestamp 0
transform 1 0 375 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_103
timestamp 0
transform 1 0 376 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_104
timestamp 0
transform 1 0 377 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_105
timestamp 0
transform 1 0 378 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_106
timestamp 0
transform 1 0 379 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_107
timestamp 0
transform 1 0 380 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_108
timestamp 0
transform 1 0 381 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_109
timestamp 0
transform 1 0 382 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_110
timestamp 0
transform 1 0 383 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_111
timestamp 0
transform 1 0 384 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_112
timestamp 0
transform 1 0 385 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_113
timestamp 0
transform 1 0 386 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_114
timestamp 0
transform 1 0 387 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_115
timestamp 0
transform 1 0 388 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_116
timestamp 0
transform 1 0 389 0 1 2552
box 0 0 1 1
use s8iom0_vdda_lvc_pad  vdd3v3lclamp[0]
timestamp 0
transform 1 0 390 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_118
timestamp 0
transform 1 0 465 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_119
timestamp 0
transform 1 0 466 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_120
timestamp 0
transform 1 0 467 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_121
timestamp 0
transform 1 0 468 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_122
timestamp 0
transform 1 0 469 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_123
timestamp 0
transform 1 0 470 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_124
timestamp 0
transform 1 0 471 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_125
timestamp 0
transform 1 0 472 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_126
timestamp 0
transform 1 0 473 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_127
timestamp 0
transform 1 0 474 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_128
timestamp 0
transform 1 0 475 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_129
timestamp 0
transform 1 0 476 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_130
timestamp 0
transform 1 0 477 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_131
timestamp 0
transform 1 0 478 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_132
timestamp 0
transform 1 0 479 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_133
timestamp 0
transform 1 0 480 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_134
timestamp 0
transform 1 0 481 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_135
timestamp 0
transform 1 0 482 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_136
timestamp 0
transform 1 0 483 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_137
timestamp 0
transform 1 0 484 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_138
timestamp 0
transform 1 0 485 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_139
timestamp 0
transform 1 0 486 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_140
timestamp 0
transform 1 0 487 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_141
timestamp 0
transform 1 0 488 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_142
timestamp 0
transform 1 0 489 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_143
timestamp 0
transform 1 0 490 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_144
timestamp 0
transform 1 0 491 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_145
timestamp 0
transform 1 0 492 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_146
timestamp 0
transform 1 0 493 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_147
timestamp 0
transform 1 0 494 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_148
timestamp 0
transform 1 0 495 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_149
timestamp 0
transform 1 0 496 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_150
timestamp 0
transform 1 0 497 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_151
timestamp 0
transform 1 0 498 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_152
timestamp 0
transform 1 0 499 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_153
timestamp 0
transform 1 0 500 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_154
timestamp 0
transform 1 0 501 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_155
timestamp 0
transform 1 0 502 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_156
timestamp 0
transform 1 0 503 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_157
timestamp 0
transform 1 0 504 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_158
timestamp 0
transform 1 0 505 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_159
timestamp 0
transform 1 0 506 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_160
timestamp 0
transform 1 0 507 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_161
timestamp 0
transform 1 0 508 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_162
timestamp 0
transform 1 0 509 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_163
timestamp 0
transform 1 0 510 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_164
timestamp 0
transform 1 0 511 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_165
timestamp 0
transform 1 0 512 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_166
timestamp 0
transform 1 0 513 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_167
timestamp 0
transform 1 0 514 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_168
timestamp 0
transform 1 0 515 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_169
timestamp 0
transform 1 0 516 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_170
timestamp 0
transform 1 0 517 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_171
timestamp 0
transform 1 0 518 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_172
timestamp 0
transform 1 0 519 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_173
timestamp 0
transform 1 0 520 0 1 2552
box 0 0 1 1
use s8iom0_vccd_hvc_pad  vdd1v8hclamp[0]
timestamp 0
transform 1 0 521 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_175
timestamp 0
transform 1 0 596 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_176
timestamp 0
transform 1 0 597 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_177
timestamp 0
transform 1 0 598 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_178
timestamp 0
transform 1 0 599 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_179
timestamp 0
transform 1 0 600 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_180
timestamp 0
transform 1 0 601 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_181
timestamp 0
transform 1 0 602 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_182
timestamp 0
transform 1 0 603 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_183
timestamp 0
transform 1 0 604 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_184
timestamp 0
transform 1 0 605 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_185
timestamp 0
transform 1 0 606 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_186
timestamp 0
transform 1 0 607 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_187
timestamp 0
transform 1 0 608 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_188
timestamp 0
transform 1 0 609 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_189
timestamp 0
transform 1 0 610 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_190
timestamp 0
transform 1 0 611 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_191
timestamp 0
transform 1 0 612 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_192
timestamp 0
transform 1 0 613 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_193
timestamp 0
transform 1 0 614 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_194
timestamp 0
transform 1 0 615 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_195
timestamp 0
transform 1 0 616 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_196
timestamp 0
transform 1 0 617 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_197
timestamp 0
transform 1 0 618 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_198
timestamp 0
transform 1 0 619 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_199
timestamp 0
transform 1 0 620 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_200
timestamp 0
transform 1 0 621 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_201
timestamp 0
transform 1 0 622 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_202
timestamp 0
transform 1 0 623 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_203
timestamp 0
transform 1 0 624 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_204
timestamp 0
transform 1 0 625 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_205
timestamp 0
transform 1 0 626 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_206
timestamp 0
transform 1 0 627 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_207
timestamp 0
transform 1 0 628 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_208
timestamp 0
transform 1 0 629 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_209
timestamp 0
transform 1 0 630 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_210
timestamp 0
transform 1 0 631 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_211
timestamp 0
transform 1 0 632 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_212
timestamp 0
transform 1 0 633 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_213
timestamp 0
transform 1 0 634 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_214
timestamp 0
transform 1 0 635 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_215
timestamp 0
transform 1 0 636 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_216
timestamp 0
transform 1 0 637 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_217
timestamp 0
transform 1 0 638 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_218
timestamp 0
transform 1 0 639 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_219
timestamp 0
transform 1 0 640 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_220
timestamp 0
transform 1 0 641 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_221
timestamp 0
transform 1 0 642 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_222
timestamp 0
transform 1 0 643 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_223
timestamp 0
transform 1 0 644 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_224
timestamp 0
transform 1 0 645 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_225
timestamp 0
transform 1 0 646 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_226
timestamp 0
transform 1 0 647 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_227
timestamp 0
transform 1 0 648 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_228
timestamp 0
transform 1 0 649 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_229
timestamp 0
transform 1 0 650 0 1 2552
box 0 0 1 1
use s8iom0_vssa_hvc_pad  vsshclamp[0]
timestamp 0
transform 1 0 651 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_231
timestamp 0
transform 1 0 726 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_232
timestamp 0
transform 1 0 727 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_233
timestamp 0
transform 1 0 728 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_234
timestamp 0
transform 1 0 729 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_235
timestamp 0
transform 1 0 730 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_236
timestamp 0
transform 1 0 731 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_237
timestamp 0
transform 1 0 732 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_238
timestamp 0
transform 1 0 733 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_239
timestamp 0
transform 1 0 734 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_240
timestamp 0
transform 1 0 735 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_241
timestamp 0
transform 1 0 736 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_242
timestamp 0
transform 1 0 737 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_243
timestamp 0
transform 1 0 738 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_244
timestamp 0
transform 1 0 739 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_245
timestamp 0
transform 1 0 740 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_246
timestamp 0
transform 1 0 741 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_247
timestamp 0
transform 1 0 742 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_248
timestamp 0
transform 1 0 743 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_249
timestamp 0
transform 1 0 744 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_250
timestamp 0
transform 1 0 745 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_251
timestamp 0
transform 1 0 746 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_252
timestamp 0
transform 1 0 747 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_253
timestamp 0
transform 1 0 748 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_254
timestamp 0
transform 1 0 749 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_255
timestamp 0
transform 1 0 750 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_256
timestamp 0
transform 1 0 751 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_257
timestamp 0
transform 1 0 752 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_258
timestamp 0
transform 1 0 753 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_259
timestamp 0
transform 1 0 754 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_260
timestamp 0
transform 1 0 755 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_261
timestamp 0
transform 1 0 756 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_262
timestamp 0
transform 1 0 757 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_263
timestamp 0
transform 1 0 758 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_264
timestamp 0
transform 1 0 759 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_265
timestamp 0
transform 1 0 760 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_266
timestamp 0
transform 1 0 761 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_267
timestamp 0
transform 1 0 762 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_268
timestamp 0
transform 1 0 763 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_269
timestamp 0
transform 1 0 764 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_270
timestamp 0
transform 1 0 765 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_271
timestamp 0
transform 1 0 766 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_272
timestamp 0
transform 1 0 767 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_273
timestamp 0
transform 1 0 768 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_274
timestamp 0
transform 1 0 769 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_275
timestamp 0
transform 1 0 770 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_276
timestamp 0
transform 1 0 771 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_277
timestamp 0
transform 1 0 772 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_278
timestamp 0
transform 1 0 773 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_279
timestamp 0
transform 1 0 774 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_280
timestamp 0
transform 1 0 775 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_281
timestamp 0
transform 1 0 776 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_282
timestamp 0
transform 1 0 777 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_283
timestamp 0
transform 1 0 778 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_284
timestamp 0
transform 1 0 779 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_285
timestamp 0
transform 1 0 780 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_286
timestamp 0
transform 1 0 781 0 1 2552
box 0 0 1 1
use s8iom0_vssa_lvc_pad  vssalclamp
timestamp 0
transform 1 0 782 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_288
timestamp 0
transform 1 0 857 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_289
timestamp 0
transform 1 0 858 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_290
timestamp 0
transform 1 0 859 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_291
timestamp 0
transform 1 0 860 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_292
timestamp 0
transform 1 0 861 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_293
timestamp 0
transform 1 0 862 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_294
timestamp 0
transform 1 0 863 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_295
timestamp 0
transform 1 0 864 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_296
timestamp 0
transform 1 0 865 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_297
timestamp 0
transform 1 0 866 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_298
timestamp 0
transform 1 0 867 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_299
timestamp 0
transform 1 0 868 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_300
timestamp 0
transform 1 0 869 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_301
timestamp 0
transform 1 0 870 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_302
timestamp 0
transform 1 0 871 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_303
timestamp 0
transform 1 0 872 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_304
timestamp 0
transform 1 0 873 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_305
timestamp 0
transform 1 0 874 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_306
timestamp 0
transform 1 0 875 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_307
timestamp 0
transform 1 0 876 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_308
timestamp 0
transform 1 0 877 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_309
timestamp 0
transform 1 0 878 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_310
timestamp 0
transform 1 0 879 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_311
timestamp 0
transform 1 0 880 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_312
timestamp 0
transform 1 0 881 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_313
timestamp 0
transform 1 0 882 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_314
timestamp 0
transform 1 0 883 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_315
timestamp 0
transform 1 0 884 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_316
timestamp 0
transform 1 0 885 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_317
timestamp 0
transform 1 0 886 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_318
timestamp 0
transform 1 0 887 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_319
timestamp 0
transform 1 0 888 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_320
timestamp 0
transform 1 0 889 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_321
timestamp 0
transform 1 0 890 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_322
timestamp 0
transform 1 0 891 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_323
timestamp 0
transform 1 0 892 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_324
timestamp 0
transform 1 0 893 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_325
timestamp 0
transform 1 0 894 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_326
timestamp 0
transform 1 0 895 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_327
timestamp 0
transform 1 0 896 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_328
timestamp 0
transform 1 0 897 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_329
timestamp 0
transform 1 0 898 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_330
timestamp 0
transform 1 0 899 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_331
timestamp 0
transform 1 0 900 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_332
timestamp 0
transform 1 0 901 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_333
timestamp 0
transform 1 0 902 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_334
timestamp 0
transform 1 0 903 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_335
timestamp 0
transform 1 0 904 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_336
timestamp 0
transform 1 0 905 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_337
timestamp 0
transform 1 0 906 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_338
timestamp 0
transform 1 0 907 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_339
timestamp 0
transform 1 0 908 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_340
timestamp 0
transform 1 0 909 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_341
timestamp 0
transform 1 0 910 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_342
timestamp 0
transform 1 0 911 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_343
timestamp 0
transform 1 0 912 0 1 2552
box 0 0 1 1
use s8iom0_gpiov2_pad  gpio_pad[8]
timestamp 0
transform 1 0 913 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_345
timestamp 0
transform 1 0 993 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_346
timestamp 0
transform 1 0 994 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_347
timestamp 0
transform 1 0 995 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_348
timestamp 0
transform 1 0 996 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_349
timestamp 0
transform 1 0 997 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_350
timestamp 0
transform 1 0 998 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_351
timestamp 0
transform 1 0 999 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_352
timestamp 0
transform 1 0 1000 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_353
timestamp 0
transform 1 0 1001 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_354
timestamp 0
transform 1 0 1002 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_355
timestamp 0
transform 1 0 1003 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_356
timestamp 0
transform 1 0 1004 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_357
timestamp 0
transform 1 0 1005 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_358
timestamp 0
transform 1 0 1006 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_359
timestamp 0
transform 1 0 1007 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_360
timestamp 0
transform 1 0 1008 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_361
timestamp 0
transform 1 0 1009 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_362
timestamp 0
transform 1 0 1010 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_363
timestamp 0
transform 1 0 1011 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_364
timestamp 0
transform 1 0 1012 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_365
timestamp 0
transform 1 0 1013 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_366
timestamp 0
transform 1 0 1014 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_367
timestamp 0
transform 1 0 1015 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_368
timestamp 0
transform 1 0 1016 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_369
timestamp 0
transform 1 0 1017 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_370
timestamp 0
transform 1 0 1018 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_371
timestamp 0
transform 1 0 1019 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_372
timestamp 0
transform 1 0 1020 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_373
timestamp 0
transform 1 0 1021 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_374
timestamp 0
transform 1 0 1022 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_375
timestamp 0
transform 1 0 1023 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_376
timestamp 0
transform 1 0 1024 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_377
timestamp 0
transform 1 0 1025 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_378
timestamp 0
transform 1 0 1026 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_379
timestamp 0
transform 1 0 1027 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_380
timestamp 0
transform 1 0 1028 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_381
timestamp 0
transform 1 0 1029 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_382
timestamp 0
transform 1 0 1030 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_383
timestamp 0
transform 1 0 1031 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_384
timestamp 0
transform 1 0 1032 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_385
timestamp 0
transform 1 0 1033 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_386
timestamp 0
transform 1 0 1034 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_387
timestamp 0
transform 1 0 1035 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_388
timestamp 0
transform 1 0 1036 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_389
timestamp 0
transform 1 0 1037 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_390
timestamp 0
transform 1 0 1038 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_391
timestamp 0
transform 1 0 1039 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_392
timestamp 0
transform 1 0 1040 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_393
timestamp 0
transform 1 0 1041 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_394
timestamp 0
transform 1 0 1042 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_395
timestamp 0
transform 1 0 1043 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_396
timestamp 0
transform 1 0 1044 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_397
timestamp 0
transform 1 0 1045 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_398
timestamp 0
transform 1 0 1046 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_399
timestamp 0
transform 1 0 1047 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_400
timestamp 0
transform 1 0 1048 0 1 2552
box 0 0 1 1
use s8iom0_gpiov2_pad  gpio_pad[7]
timestamp 0
transform 1 0 1049 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_402
timestamp 0
transform 1 0 1129 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_403
timestamp 0
transform 1 0 1130 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_404
timestamp 0
transform 1 0 1131 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_405
timestamp 0
transform 1 0 1132 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_406
timestamp 0
transform 1 0 1133 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_407
timestamp 0
transform 1 0 1134 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_408
timestamp 0
transform 1 0 1135 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_409
timestamp 0
transform 1 0 1136 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_410
timestamp 0
transform 1 0 1137 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_411
timestamp 0
transform 1 0 1138 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_412
timestamp 0
transform 1 0 1139 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_413
timestamp 0
transform 1 0 1140 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_414
timestamp 0
transform 1 0 1141 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_415
timestamp 0
transform 1 0 1142 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_416
timestamp 0
transform 1 0 1143 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_417
timestamp 0
transform 1 0 1144 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_418
timestamp 0
transform 1 0 1145 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_419
timestamp 0
transform 1 0 1146 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_420
timestamp 0
transform 1 0 1147 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_421
timestamp 0
transform 1 0 1148 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_422
timestamp 0
transform 1 0 1149 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_423
timestamp 0
transform 1 0 1150 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_424
timestamp 0
transform 1 0 1151 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_425
timestamp 0
transform 1 0 1152 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_426
timestamp 0
transform 1 0 1153 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_427
timestamp 0
transform 1 0 1154 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_428
timestamp 0
transform 1 0 1155 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_429
timestamp 0
transform 1 0 1156 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_430
timestamp 0
transform 1 0 1157 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_431
timestamp 0
transform 1 0 1158 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_432
timestamp 0
transform 1 0 1159 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_433
timestamp 0
transform 1 0 1160 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_434
timestamp 0
transform 1 0 1161 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_435
timestamp 0
transform 1 0 1162 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_436
timestamp 0
transform 1 0 1163 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_437
timestamp 0
transform 1 0 1164 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_438
timestamp 0
transform 1 0 1165 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_439
timestamp 0
transform 1 0 1166 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_440
timestamp 0
transform 1 0 1167 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_441
timestamp 0
transform 1 0 1168 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_442
timestamp 0
transform 1 0 1169 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_443
timestamp 0
transform 1 0 1170 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_444
timestamp 0
transform 1 0 1171 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_445
timestamp 0
transform 1 0 1172 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_446
timestamp 0
transform 1 0 1173 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_447
timestamp 0
transform 1 0 1174 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_448
timestamp 0
transform 1 0 1175 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_449
timestamp 0
transform 1 0 1176 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_450
timestamp 0
transform 1 0 1177 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_451
timestamp 0
transform 1 0 1178 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_452
timestamp 0
transform 1 0 1179 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_453
timestamp 0
transform 1 0 1180 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_454
timestamp 0
transform 1 0 1181 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_455
timestamp 0
transform 1 0 1182 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_456
timestamp 0
transform 1 0 1183 0 1 2552
box 0 0 1 1
use s8iom0_gpiov2_pad  gpio_pad[6]
timestamp 0
transform 1 0 1184 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_458
timestamp 0
transform 1 0 1264 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_459
timestamp 0
transform 1 0 1265 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_460
timestamp 0
transform 1 0 1266 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_461
timestamp 0
transform 1 0 1267 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_462
timestamp 0
transform 1 0 1268 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_463
timestamp 0
transform 1 0 1269 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_464
timestamp 0
transform 1 0 1270 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_465
timestamp 0
transform 1 0 1271 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_466
timestamp 0
transform 1 0 1272 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_467
timestamp 0
transform 1 0 1273 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_468
timestamp 0
transform 1 0 1274 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_469
timestamp 0
transform 1 0 1275 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_470
timestamp 0
transform 1 0 1276 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_471
timestamp 0
transform 1 0 1277 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_472
timestamp 0
transform 1 0 1278 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_473
timestamp 0
transform 1 0 1279 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_474
timestamp 0
transform 1 0 1280 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_475
timestamp 0
transform 1 0 1281 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_476
timestamp 0
transform 1 0 1282 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_477
timestamp 0
transform 1 0 1283 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_478
timestamp 0
transform 1 0 1284 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_479
timestamp 0
transform 1 0 1285 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_480
timestamp 0
transform 1 0 1286 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_481
timestamp 0
transform 1 0 1287 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_482
timestamp 0
transform 1 0 1288 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_483
timestamp 0
transform 1 0 1289 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_484
timestamp 0
transform 1 0 1290 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_485
timestamp 0
transform 1 0 1291 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_486
timestamp 0
transform 1 0 1292 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_487
timestamp 0
transform 1 0 1293 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_488
timestamp 0
transform 1 0 1294 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_489
timestamp 0
transform 1 0 1295 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_490
timestamp 0
transform 1 0 1296 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_491
timestamp 0
transform 1 0 1297 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_492
timestamp 0
transform 1 0 1298 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_493
timestamp 0
transform 1 0 1299 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_494
timestamp 0
transform 1 0 1300 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_495
timestamp 0
transform 1 0 1301 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_496
timestamp 0
transform 1 0 1302 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_497
timestamp 0
transform 1 0 1303 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_498
timestamp 0
transform 1 0 1304 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_499
timestamp 0
transform 1 0 1305 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_500
timestamp 0
transform 1 0 1306 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_501
timestamp 0
transform 1 0 1307 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_502
timestamp 0
transform 1 0 1308 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_503
timestamp 0
transform 1 0 1309 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_504
timestamp 0
transform 1 0 1310 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_505
timestamp 0
transform 1 0 1311 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_506
timestamp 0
transform 1 0 1312 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_507
timestamp 0
transform 1 0 1313 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_508
timestamp 0
transform 1 0 1314 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_509
timestamp 0
transform 1 0 1315 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_510
timestamp 0
transform 1 0 1316 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_511
timestamp 0
transform 1 0 1317 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_512
timestamp 0
transform 1 0 1318 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_513
timestamp 0
transform 1 0 1319 0 1 2552
box 0 0 1 1
use s8iom0_gpiov2_pad  gpio_pad[5]
timestamp 0
transform 1 0 1320 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_515
timestamp 0
transform 1 0 1400 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_516
timestamp 0
transform 1 0 1401 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_517
timestamp 0
transform 1 0 1402 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_518
timestamp 0
transform 1 0 1403 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_519
timestamp 0
transform 1 0 1404 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_520
timestamp 0
transform 1 0 1405 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_521
timestamp 0
transform 1 0 1406 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_522
timestamp 0
transform 1 0 1407 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_523
timestamp 0
transform 1 0 1408 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_524
timestamp 0
transform 1 0 1409 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_525
timestamp 0
transform 1 0 1410 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_526
timestamp 0
transform 1 0 1411 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_527
timestamp 0
transform 1 0 1412 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_528
timestamp 0
transform 1 0 1413 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_529
timestamp 0
transform 1 0 1414 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_530
timestamp 0
transform 1 0 1415 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_531
timestamp 0
transform 1 0 1416 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_532
timestamp 0
transform 1 0 1417 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_533
timestamp 0
transform 1 0 1418 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_534
timestamp 0
transform 1 0 1419 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_535
timestamp 0
transform 1 0 1420 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_536
timestamp 0
transform 1 0 1421 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_537
timestamp 0
transform 1 0 1422 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_538
timestamp 0
transform 1 0 1423 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_539
timestamp 0
transform 1 0 1424 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_540
timestamp 0
transform 1 0 1425 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_541
timestamp 0
transform 1 0 1426 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_542
timestamp 0
transform 1 0 1427 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_543
timestamp 0
transform 1 0 1428 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_544
timestamp 0
transform 1 0 1429 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_545
timestamp 0
transform 1 0 1430 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_546
timestamp 0
transform 1 0 1431 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_547
timestamp 0
transform 1 0 1432 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_548
timestamp 0
transform 1 0 1433 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_549
timestamp 0
transform 1 0 1434 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_550
timestamp 0
transform 1 0 1435 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_551
timestamp 0
transform 1 0 1436 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_552
timestamp 0
transform 1 0 1437 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_553
timestamp 0
transform 1 0 1438 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_554
timestamp 0
transform 1 0 1439 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_555
timestamp 0
transform 1 0 1440 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_556
timestamp 0
transform 1 0 1441 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_557
timestamp 0
transform 1 0 1442 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_558
timestamp 0
transform 1 0 1443 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_559
timestamp 0
transform 1 0 1444 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_560
timestamp 0
transform 1 0 1445 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_561
timestamp 0
transform 1 0 1446 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_562
timestamp 0
transform 1 0 1447 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_563
timestamp 0
transform 1 0 1448 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_564
timestamp 0
transform 1 0 1449 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_565
timestamp 0
transform 1 0 1450 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_566
timestamp 0
transform 1 0 1451 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_567
timestamp 0
transform 1 0 1452 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_568
timestamp 0
transform 1 0 1453 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_569
timestamp 0
transform 1 0 1454 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_570
timestamp 0
transform 1 0 1455 0 1 2552
box 0 0 1 1
use s8iom0_gpiov2_pad  gpio_pad[15]
timestamp 0
transform 1 0 1456 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_572
timestamp 0
transform 1 0 1536 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_573
timestamp 0
transform 1 0 1537 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_574
timestamp 0
transform 1 0 1538 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_575
timestamp 0
transform 1 0 1539 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_576
timestamp 0
transform 1 0 1540 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_577
timestamp 0
transform 1 0 1541 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_578
timestamp 0
transform 1 0 1542 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_579
timestamp 0
transform 1 0 1543 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_580
timestamp 0
transform 1 0 1544 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_581
timestamp 0
transform 1 0 1545 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_582
timestamp 0
transform 1 0 1546 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_583
timestamp 0
transform 1 0 1547 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_584
timestamp 0
transform 1 0 1548 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_585
timestamp 0
transform 1 0 1549 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_586
timestamp 0
transform 1 0 1550 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_587
timestamp 0
transform 1 0 1551 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_588
timestamp 0
transform 1 0 1552 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_589
timestamp 0
transform 1 0 1553 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_590
timestamp 0
transform 1 0 1554 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_591
timestamp 0
transform 1 0 1555 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_592
timestamp 0
transform 1 0 1556 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_593
timestamp 0
transform 1 0 1557 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_594
timestamp 0
transform 1 0 1558 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_595
timestamp 0
transform 1 0 1559 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_596
timestamp 0
transform 1 0 1560 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_597
timestamp 0
transform 1 0 1561 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_598
timestamp 0
transform 1 0 1562 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_599
timestamp 0
transform 1 0 1563 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_600
timestamp 0
transform 1 0 1564 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_601
timestamp 0
transform 1 0 1565 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_602
timestamp 0
transform 1 0 1566 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_603
timestamp 0
transform 1 0 1567 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_604
timestamp 0
transform 1 0 1568 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_605
timestamp 0
transform 1 0 1569 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_606
timestamp 0
transform 1 0 1570 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_607
timestamp 0
transform 1 0 1571 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_608
timestamp 0
transform 1 0 1572 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_609
timestamp 0
transform 1 0 1573 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_610
timestamp 0
transform 1 0 1574 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_611
timestamp 0
transform 1 0 1575 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_612
timestamp 0
transform 1 0 1576 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_613
timestamp 0
transform 1 0 1577 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_614
timestamp 0
transform 1 0 1578 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_615
timestamp 0
transform 1 0 1579 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_616
timestamp 0
transform 1 0 1580 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_617
timestamp 0
transform 1 0 1581 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_618
timestamp 0
transform 1 0 1582 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_619
timestamp 0
transform 1 0 1583 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_620
timestamp 0
transform 1 0 1584 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_621
timestamp 0
transform 1 0 1585 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_622
timestamp 0
transform 1 0 1586 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_623
timestamp 0
transform 1 0 1587 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_624
timestamp 0
transform 1 0 1588 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_625
timestamp 0
transform 1 0 1589 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_626
timestamp 0
transform 1 0 1590 0 1 2552
box 0 0 1 1
use s8iom0_gpiov2_pad  gpio_pad[14]
timestamp 0
transform 1 0 1591 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_628
timestamp 0
transform 1 0 1671 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_629
timestamp 0
transform 1 0 1672 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_630
timestamp 0
transform 1 0 1673 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_631
timestamp 0
transform 1 0 1674 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_632
timestamp 0
transform 1 0 1675 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_633
timestamp 0
transform 1 0 1676 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_634
timestamp 0
transform 1 0 1677 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_635
timestamp 0
transform 1 0 1678 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_636
timestamp 0
transform 1 0 1679 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_637
timestamp 0
transform 1 0 1680 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_638
timestamp 0
transform 1 0 1681 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_639
timestamp 0
transform 1 0 1682 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_640
timestamp 0
transform 1 0 1683 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_641
timestamp 0
transform 1 0 1684 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_642
timestamp 0
transform 1 0 1685 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_643
timestamp 0
transform 1 0 1686 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_644
timestamp 0
transform 1 0 1687 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_645
timestamp 0
transform 1 0 1688 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_646
timestamp 0
transform 1 0 1689 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_647
timestamp 0
transform 1 0 1690 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_648
timestamp 0
transform 1 0 1691 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_649
timestamp 0
transform 1 0 1692 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_650
timestamp 0
transform 1 0 1693 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_651
timestamp 0
transform 1 0 1694 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_652
timestamp 0
transform 1 0 1695 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_653
timestamp 0
transform 1 0 1696 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_654
timestamp 0
transform 1 0 1697 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_655
timestamp 0
transform 1 0 1698 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_656
timestamp 0
transform 1 0 1699 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_657
timestamp 0
transform 1 0 1700 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_658
timestamp 0
transform 1 0 1701 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_659
timestamp 0
transform 1 0 1702 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_660
timestamp 0
transform 1 0 1703 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_661
timestamp 0
transform 1 0 1704 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_662
timestamp 0
transform 1 0 1705 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_663
timestamp 0
transform 1 0 1706 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_664
timestamp 0
transform 1 0 1707 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_665
timestamp 0
transform 1 0 1708 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_666
timestamp 0
transform 1 0 1709 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_667
timestamp 0
transform 1 0 1710 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_668
timestamp 0
transform 1 0 1711 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_669
timestamp 0
transform 1 0 1712 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_670
timestamp 0
transform 1 0 1713 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_671
timestamp 0
transform 1 0 1714 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_672
timestamp 0
transform 1 0 1715 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_673
timestamp 0
transform 1 0 1716 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_674
timestamp 0
transform 1 0 1717 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_675
timestamp 0
transform 1 0 1718 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_676
timestamp 0
transform 1 0 1719 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_677
timestamp 0
transform 1 0 1720 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_678
timestamp 0
transform 1 0 1721 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_679
timestamp 0
transform 1 0 1722 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_680
timestamp 0
transform 1 0 1723 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_681
timestamp 0
transform 1 0 1724 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_682
timestamp 0
transform 1 0 1725 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_683
timestamp 0
transform 1 0 1726 0 1 2552
box 0 0 1 1
use s8iom0_gpiov2_pad  gpio_pad[13]
timestamp 0
transform 1 0 1727 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_685
timestamp 0
transform 1 0 1807 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_686
timestamp 0
transform 1 0 1808 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_687
timestamp 0
transform 1 0 1809 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_688
timestamp 0
transform 1 0 1810 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_689
timestamp 0
transform 1 0 1811 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_690
timestamp 0
transform 1 0 1812 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_691
timestamp 0
transform 1 0 1813 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_692
timestamp 0
transform 1 0 1814 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_693
timestamp 0
transform 1 0 1815 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_694
timestamp 0
transform 1 0 1816 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_695
timestamp 0
transform 1 0 1817 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_696
timestamp 0
transform 1 0 1818 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_697
timestamp 0
transform 1 0 1819 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_698
timestamp 0
transform 1 0 1820 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_699
timestamp 0
transform 1 0 1821 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_700
timestamp 0
transform 1 0 1822 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_701
timestamp 0
transform 1 0 1823 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_702
timestamp 0
transform 1 0 1824 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_703
timestamp 0
transform 1 0 1825 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_704
timestamp 0
transform 1 0 1826 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_705
timestamp 0
transform 1 0 1827 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_706
timestamp 0
transform 1 0 1828 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_707
timestamp 0
transform 1 0 1829 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_708
timestamp 0
transform 1 0 1830 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_709
timestamp 0
transform 1 0 1831 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_710
timestamp 0
transform 1 0 1832 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_711
timestamp 0
transform 1 0 1833 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_712
timestamp 0
transform 1 0 1834 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_713
timestamp 0
transform 1 0 1835 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_714
timestamp 0
transform 1 0 1836 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_715
timestamp 0
transform 1 0 1837 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_716
timestamp 0
transform 1 0 1838 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_717
timestamp 0
transform 1 0 1839 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_718
timestamp 0
transform 1 0 1840 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_719
timestamp 0
transform 1 0 1841 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_720
timestamp 0
transform 1 0 1842 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_721
timestamp 0
transform 1 0 1843 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_722
timestamp 0
transform 1 0 1844 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_723
timestamp 0
transform 1 0 1845 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_724
timestamp 0
transform 1 0 1846 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_725
timestamp 0
transform 1 0 1847 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_726
timestamp 0
transform 1 0 1848 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_727
timestamp 0
transform 1 0 1849 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_728
timestamp 0
transform 1 0 1850 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_729
timestamp 0
transform 1 0 1851 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_730
timestamp 0
transform 1 0 1852 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_731
timestamp 0
transform 1 0 1853 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_732
timestamp 0
transform 1 0 1854 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_733
timestamp 0
transform 1 0 1855 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_734
timestamp 0
transform 1 0 1856 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_735
timestamp 0
transform 1 0 1857 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_736
timestamp 0
transform 1 0 1858 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_737
timestamp 0
transform 1 0 1859 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_738
timestamp 0
transform 1 0 1860 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_739
timestamp 0
transform 1 0 1861 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_740
timestamp 0
transform 1 0 1862 0 1 2552
box 0 0 1 1
use s8iom0_gpiov2_pad  gpio_pad[12]
timestamp 0
transform 1 0 1863 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_742
timestamp 0
transform 1 0 1943 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_743
timestamp 0
transform 1 0 1944 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_744
timestamp 0
transform 1 0 1945 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_745
timestamp 0
transform 1 0 1946 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_746
timestamp 0
transform 1 0 1947 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_747
timestamp 0
transform 1 0 1948 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_748
timestamp 0
transform 1 0 1949 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_749
timestamp 0
transform 1 0 1950 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_750
timestamp 0
transform 1 0 1951 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_751
timestamp 0
transform 1 0 1952 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_752
timestamp 0
transform 1 0 1953 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_753
timestamp 0
transform 1 0 1954 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_754
timestamp 0
transform 1 0 1955 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_755
timestamp 0
transform 1 0 1956 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_756
timestamp 0
transform 1 0 1957 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_757
timestamp 0
transform 1 0 1958 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_758
timestamp 0
transform 1 0 1959 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_759
timestamp 0
transform 1 0 1960 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_760
timestamp 0
transform 1 0 1961 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_761
timestamp 0
transform 1 0 1962 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_762
timestamp 0
transform 1 0 1963 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_763
timestamp 0
transform 1 0 1964 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_764
timestamp 0
transform 1 0 1965 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_765
timestamp 0
transform 1 0 1966 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_766
timestamp 0
transform 1 0 1967 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_767
timestamp 0
transform 1 0 1968 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_768
timestamp 0
transform 1 0 1969 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_769
timestamp 0
transform 1 0 1970 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_770
timestamp 0
transform 1 0 1971 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_771
timestamp 0
transform 1 0 1972 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_772
timestamp 0
transform 1 0 1973 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_773
timestamp 0
transform 1 0 1974 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_774
timestamp 0
transform 1 0 1975 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_775
timestamp 0
transform 1 0 1976 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_776
timestamp 0
transform 1 0 1977 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_777
timestamp 0
transform 1 0 1978 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_778
timestamp 0
transform 1 0 1979 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_779
timestamp 0
transform 1 0 1980 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_780
timestamp 0
transform 1 0 1981 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_781
timestamp 0
transform 1 0 1982 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_782
timestamp 0
transform 1 0 1983 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_783
timestamp 0
transform 1 0 1984 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_784
timestamp 0
transform 1 0 1985 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_785
timestamp 0
transform 1 0 1986 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_786
timestamp 0
transform 1 0 1987 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_787
timestamp 0
transform 1 0 1988 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_788
timestamp 0
transform 1 0 1989 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_789
timestamp 0
transform 1 0 1990 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_790
timestamp 0
transform 1 0 1991 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_791
timestamp 0
transform 1 0 1992 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_792
timestamp 0
transform 1 0 1993 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_793
timestamp 0
transform 1 0 1994 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_794
timestamp 0
transform 1 0 1995 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_795
timestamp 0
transform 1 0 1996 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_796
timestamp 0
transform 1 0 1997 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_797
timestamp 0
transform 1 0 1998 0 1 2552
box 0 0 1 1
use s8iom0_gpiov2_pad  irq_pad
timestamp 0
transform 1 0 1999 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_799
timestamp 0
transform 1 0 2079 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_800
timestamp 0
transform 1 0 2080 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_801
timestamp 0
transform 1 0 2081 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_802
timestamp 0
transform 1 0 2082 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_803
timestamp 0
transform 1 0 2083 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_804
timestamp 0
transform 1 0 2084 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_805
timestamp 0
transform 1 0 2085 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_806
timestamp 0
transform 1 0 2086 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_807
timestamp 0
transform 1 0 2087 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_808
timestamp 0
transform 1 0 2088 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_809
timestamp 0
transform 1 0 2089 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_810
timestamp 0
transform 1 0 2090 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_811
timestamp 0
transform 1 0 2091 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_812
timestamp 0
transform 1 0 2092 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_813
timestamp 0
transform 1 0 2093 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_814
timestamp 0
transform 1 0 2094 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_815
timestamp 0
transform 1 0 2095 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_816
timestamp 0
transform 1 0 2096 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_817
timestamp 0
transform 1 0 2097 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_818
timestamp 0
transform 1 0 2098 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_819
timestamp 0
transform 1 0 2099 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_820
timestamp 0
transform 1 0 2100 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_821
timestamp 0
transform 1 0 2101 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_822
timestamp 0
transform 1 0 2102 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_823
timestamp 0
transform 1 0 2103 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_824
timestamp 0
transform 1 0 2104 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_825
timestamp 0
transform 1 0 2105 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_826
timestamp 0
transform 1 0 2106 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_827
timestamp 0
transform 1 0 2107 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_828
timestamp 0
transform 1 0 2108 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_829
timestamp 0
transform 1 0 2109 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_830
timestamp 0
transform 1 0 2110 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_831
timestamp 0
transform 1 0 2111 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_832
timestamp 0
transform 1 0 2112 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_833
timestamp 0
transform 1 0 2113 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_834
timestamp 0
transform 1 0 2114 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_835
timestamp 0
transform 1 0 2115 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_836
timestamp 0
transform 1 0 2116 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_837
timestamp 0
transform 1 0 2117 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_838
timestamp 0
transform 1 0 2118 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_839
timestamp 0
transform 1 0 2119 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_840
timestamp 0
transform 1 0 2120 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_841
timestamp 0
transform 1 0 2121 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_842
timestamp 0
transform 1 0 2122 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_843
timestamp 0
transform 1 0 2123 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_844
timestamp 0
transform 1 0 2124 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_845
timestamp 0
transform 1 0 2125 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_846
timestamp 0
transform 1 0 2126 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_847
timestamp 0
transform 1 0 2127 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_848
timestamp 0
transform 1 0 2128 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_849
timestamp 0
transform 1 0 2129 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_850
timestamp 0
transform 1 0 2130 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_851
timestamp 0
transform 1 0 2131 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_852
timestamp 0
transform 1 0 2132 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_853
timestamp 0
transform 1 0 2133 0 1 2552
box 0 0 1 1
use s8iom0_gpiov2_pad  SDO_pad
timestamp 0
transform 1 0 2134 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_855
timestamp 0
transform 1 0 2214 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_856
timestamp 0
transform 1 0 2215 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_857
timestamp 0
transform 1 0 2216 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_858
timestamp 0
transform 1 0 2217 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_859
timestamp 0
transform 1 0 2218 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_860
timestamp 0
transform 1 0 2219 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_861
timestamp 0
transform 1 0 2220 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_862
timestamp 0
transform 1 0 2221 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_863
timestamp 0
transform 1 0 2222 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_864
timestamp 0
transform 1 0 2223 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_865
timestamp 0
transform 1 0 2224 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_866
timestamp 0
transform 1 0 2225 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_867
timestamp 0
transform 1 0 2226 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_868
timestamp 0
transform 1 0 2227 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_869
timestamp 0
transform 1 0 2228 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_870
timestamp 0
transform 1 0 2229 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_871
timestamp 0
transform 1 0 2230 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_872
timestamp 0
transform 1 0 2231 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_873
timestamp 0
transform 1 0 2232 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_874
timestamp 0
transform 1 0 2233 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_875
timestamp 0
transform 1 0 2234 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_876
timestamp 0
transform 1 0 2235 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_877
timestamp 0
transform 1 0 2236 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_878
timestamp 0
transform 1 0 2237 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_879
timestamp 0
transform 1 0 2238 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_880
timestamp 0
transform 1 0 2239 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_881
timestamp 0
transform 1 0 2240 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_882
timestamp 0
transform 1 0 2241 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_883
timestamp 0
transform 1 0 2242 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_884
timestamp 0
transform 1 0 2243 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_885
timestamp 0
transform 1 0 2244 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_886
timestamp 0
transform 1 0 2245 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_887
timestamp 0
transform 1 0 2246 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_888
timestamp 0
transform 1 0 2247 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_889
timestamp 0
transform 1 0 2248 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_890
timestamp 0
transform 1 0 2249 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_891
timestamp 0
transform 1 0 2250 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_892
timestamp 0
transform 1 0 2251 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_893
timestamp 0
transform 1 0 2252 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_894
timestamp 0
transform 1 0 2253 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_895
timestamp 0
transform 1 0 2254 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_896
timestamp 0
transform 1 0 2255 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_897
timestamp 0
transform 1 0 2256 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_898
timestamp 0
transform 1 0 2257 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_899
timestamp 0
transform 1 0 2258 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_900
timestamp 0
transform 1 0 2259 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_901
timestamp 0
transform 1 0 2260 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_902
timestamp 0
transform 1 0 2261 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_903
timestamp 0
transform 1 0 2262 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_904
timestamp 0
transform 1 0 2263 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_905
timestamp 0
transform 1 0 2264 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_906
timestamp 0
transform 1 0 2265 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_907
timestamp 0
transform 1 0 2266 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_908
timestamp 0
transform 1 0 2267 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_909
timestamp 0
transform 1 0 2268 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_910
timestamp 0
transform 1 0 2269 0 1 2552
box 0 0 1 1
use s8iom0_gpiov2_pad  SDI_pad
timestamp 0
transform 1 0 2270 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_912
timestamp 0
transform 1 0 2350 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_913
timestamp 0
transform 1 0 2351 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_914
timestamp 0
transform 1 0 2352 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_915
timestamp 0
transform 1 0 2353 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_916
timestamp 0
transform 1 0 2354 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_917
timestamp 0
transform 1 0 2355 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_918
timestamp 0
transform 1 0 2356 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_919
timestamp 0
transform 1 0 2357 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_920
timestamp 0
transform 1 0 2358 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_921
timestamp 0
transform 1 0 2359 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_922
timestamp 0
transform 1 0 2360 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_923
timestamp 0
transform 1 0 2361 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_924
timestamp 0
transform 1 0 2362 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_925
timestamp 0
transform 1 0 2363 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_926
timestamp 0
transform 1 0 2364 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_927
timestamp 0
transform 1 0 2365 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_928
timestamp 0
transform 1 0 2366 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_929
timestamp 0
transform 1 0 2367 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_930
timestamp 0
transform 1 0 2368 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_931
timestamp 0
transform 1 0 2369 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_932
timestamp 0
transform 1 0 2370 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_933
timestamp 0
transform 1 0 2371 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_934
timestamp 0
transform 1 0 2372 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_935
timestamp 0
transform 1 0 2373 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_936
timestamp 0
transform 1 0 2374 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_937
timestamp 0
transform 1 0 2375 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_938
timestamp 0
transform 1 0 2376 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_939
timestamp 0
transform 1 0 2377 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_940
timestamp 0
transform 1 0 2378 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_941
timestamp 0
transform 1 0 2379 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_942
timestamp 0
transform 1 0 2380 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_943
timestamp 0
transform 1 0 2381 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_944
timestamp 0
transform 1 0 2382 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_945
timestamp 0
transform 1 0 2383 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_946
timestamp 0
transform 1 0 2384 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_947
timestamp 0
transform 1 0 2385 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_948
timestamp 0
transform 1 0 2386 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_949
timestamp 0
transform 1 0 2387 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_950
timestamp 0
transform 1 0 2388 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_951
timestamp 0
transform 1 0 2389 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_952
timestamp 0
transform 1 0 2390 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_953
timestamp 0
transform 1 0 2391 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_954
timestamp 0
transform 1 0 2392 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_955
timestamp 0
transform 1 0 2393 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_956
timestamp 0
transform 1 0 2394 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_957
timestamp 0
transform 1 0 2395 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_958
timestamp 0
transform 1 0 2396 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_959
timestamp 0
transform 1 0 2397 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_960
timestamp 0
transform 1 0 2398 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_961
timestamp 0
transform 1 0 2399 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_962
timestamp 0
transform 1 0 2400 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_963
timestamp 0
transform 1 0 2401 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_964
timestamp 0
transform 1 0 2402 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_965
timestamp 0
transform 1 0 2403 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_966
timestamp 0
transform 1 0 2404 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_967
timestamp 0
transform 1 0 2405 0 1 2552
box 0 0 1 1
use s8iom0_gpiov2_pad  flash_csb_pad
timestamp 0
transform 1 0 2406 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_969
timestamp 0
transform 1 0 2486 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_970
timestamp 0
transform 1 0 2487 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_971
timestamp 0
transform 1 0 2488 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_972
timestamp 0
transform 1 0 2489 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_973
timestamp 0
transform 1 0 2490 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_974
timestamp 0
transform 1 0 2491 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_975
timestamp 0
transform 1 0 2492 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_976
timestamp 0
transform 1 0 2493 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_977
timestamp 0
transform 1 0 2494 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_978
timestamp 0
transform 1 0 2495 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_979
timestamp 0
transform 1 0 2496 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_980
timestamp 0
transform 1 0 2497 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_981
timestamp 0
transform 1 0 2498 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_982
timestamp 0
transform 1 0 2499 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_983
timestamp 0
transform 1 0 2500 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_984
timestamp 0
transform 1 0 2501 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_985
timestamp 0
transform 1 0 2502 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_986
timestamp 0
transform 1 0 2503 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_987
timestamp 0
transform 1 0 2504 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_988
timestamp 0
transform 1 0 2505 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_989
timestamp 0
transform 1 0 2506 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_990
timestamp 0
transform 1 0 2507 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_991
timestamp 0
transform 1 0 2508 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_992
timestamp 0
transform 1 0 2509 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_993
timestamp 0
transform 1 0 2510 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_994
timestamp 0
transform 1 0 2511 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_995
timestamp 0
transform 1 0 2512 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_996
timestamp 0
transform 1 0 2513 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_997
timestamp 0
transform 1 0 2514 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_998
timestamp 0
transform 1 0 2515 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_999
timestamp 0
transform 1 0 2516 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1000
timestamp 0
transform 1 0 2517 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1001
timestamp 0
transform 1 0 2518 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1002
timestamp 0
transform 1 0 2519 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1003
timestamp 0
transform 1 0 2520 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1004
timestamp 0
transform 1 0 2521 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1005
timestamp 0
transform 1 0 2522 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1006
timestamp 0
transform 1 0 2523 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1007
timestamp 0
transform 1 0 2524 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1008
timestamp 0
transform 1 0 2525 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1009
timestamp 0
transform 1 0 2526 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1010
timestamp 0
transform 1 0 2527 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1011
timestamp 0
transform 1 0 2528 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1012
timestamp 0
transform 1 0 2529 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1013
timestamp 0
transform 1 0 2530 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1014
timestamp 0
transform 1 0 2531 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1015
timestamp 0
transform 1 0 2532 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1016
timestamp 0
transform 1 0 2533 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1017
timestamp 0
transform 1 0 2534 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1018
timestamp 0
transform 1 0 2535 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1019
timestamp 0
transform 1 0 2536 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1020
timestamp 0
transform 1 0 2537 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1021
timestamp 0
transform 1 0 2538 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1022
timestamp 0
transform 1 0 2539 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1023
timestamp 0
transform 1 0 2540 0 1 2552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1024
timestamp 0
transform 1 0 2541 0 1 2552
box 0 0 1 1
use s8iom0_corner_pad  corner[2]
timestamp 0
transform 0 -1 204 1 0 2550
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3268
timestamp 0
transform 0 -1 198 1 0 2549
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3267
timestamp 0
transform 0 -1 198 1 0 2548
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3266
timestamp 0
transform 0 -1 198 1 0 2547
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3265
timestamp 0
transform 0 -1 198 1 0 2546
box 0 0 1 1
use s8iom0_corner_pad  corner[3]
timestamp 0
transform 1 0 2542 0 1 2546
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3264
timestamp 0
transform 0 -1 198 1 0 2545
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3263
timestamp 0
transform 0 -1 198 1 0 2544
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3262
timestamp 0
transform 0 -1 198 1 0 2543
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3261
timestamp 0
transform 0 -1 198 1 0 2542
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3260
timestamp 0
transform 0 -1 198 1 0 2541
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3259
timestamp 0
transform 0 -1 198 1 0 2540
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3258
timestamp 0
transform 0 -1 198 1 0 2539
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3257
timestamp 0
transform 0 -1 198 1 0 2538
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3256
timestamp 0
transform 0 -1 198 1 0 2537
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3255
timestamp 0
transform 0 -1 198 1 0 2536
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3254
timestamp 0
transform 0 -1 198 1 0 2535
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3253
timestamp 0
transform 0 -1 198 1 0 2534
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3252
timestamp 0
transform 0 -1 198 1 0 2533
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3251
timestamp 0
transform 0 -1 198 1 0 2532
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3250
timestamp 0
transform 0 -1 198 1 0 2531
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3249
timestamp 0
transform 0 -1 198 1 0 2530
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3248
timestamp 0
transform 0 -1 198 1 0 2529
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3247
timestamp 0
transform 0 -1 198 1 0 2528
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3246
timestamp 0
transform 0 -1 198 1 0 2527
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3245
timestamp 0
transform 0 -1 198 1 0 2526
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3244
timestamp 0
transform 0 -1 198 1 0 2525
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3243
timestamp 0
transform 0 -1 198 1 0 2524
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3242
timestamp 0
transform 0 -1 198 1 0 2523
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3241
timestamp 0
transform 0 -1 198 1 0 2522
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3240
timestamp 0
transform 0 -1 198 1 0 2521
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3239
timestamp 0
transform 0 -1 198 1 0 2520
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3238
timestamp 0
transform 0 -1 198 1 0 2519
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3237
timestamp 0
transform 0 -1 198 1 0 2518
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3236
timestamp 0
transform 0 -1 198 1 0 2517
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3235
timestamp 0
transform 0 -1 198 1 0 2516
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3234
timestamp 0
transform 0 -1 198 1 0 2515
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3233
timestamp 0
transform 0 -1 198 1 0 2514
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3232
timestamp 0
transform 0 -1 198 1 0 2513
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3231
timestamp 0
transform 0 -1 198 1 0 2512
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3230
timestamp 0
transform 0 -1 198 1 0 2511
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3229
timestamp 0
transform 0 -1 198 1 0 2510
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3228
timestamp 0
transform 0 -1 198 1 0 2509
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3227
timestamp 0
transform 0 -1 198 1 0 2508
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3226
timestamp 0
transform 0 -1 198 1 0 2507
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3225
timestamp 0
transform 0 -1 198 1 0 2506
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3224
timestamp 0
transform 0 -1 198 1 0 2505
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3223
timestamp 0
transform 0 -1 198 1 0 2504
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3222
timestamp 0
transform 0 -1 198 1 0 2503
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3221
timestamp 0
transform 0 -1 198 1 0 2502
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3220
timestamp 0
transform 0 -1 198 1 0 2501
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3219
timestamp 0
transform 0 -1 198 1 0 2500
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3218
timestamp 0
transform 0 -1 198 1 0 2499
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3217
timestamp 0
transform 0 -1 198 1 0 2498
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3216
timestamp 0
transform 0 -1 198 1 0 2497
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3215
timestamp 0
transform 0 -1 198 1 0 2496
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3214
timestamp 0
transform 0 -1 198 1 0 2495
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3213
timestamp 0
transform 0 -1 198 1 0 2494
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3212
timestamp 0
transform 0 -1 198 1 0 2493
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3211
timestamp 0
transform 0 -1 198 1 0 2492
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4770
timestamp 0
transform 0 1 2544 -1 0 2546
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4769
timestamp 0
transform 0 1 2544 -1 0 2545
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4768
timestamp 0
transform 0 1 2544 -1 0 2544
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4767
timestamp 0
transform 0 1 2544 -1 0 2543
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4766
timestamp 0
transform 0 1 2544 -1 0 2542
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4765
timestamp 0
transform 0 1 2544 -1 0 2541
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4764
timestamp 0
transform 0 1 2544 -1 0 2540
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4763
timestamp 0
transform 0 1 2544 -1 0 2539
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4762
timestamp 0
transform 0 1 2544 -1 0 2538
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4761
timestamp 0
transform 0 1 2544 -1 0 2537
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4760
timestamp 0
transform 0 1 2544 -1 0 2536
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4759
timestamp 0
transform 0 1 2544 -1 0 2535
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4758
timestamp 0
transform 0 1 2544 -1 0 2534
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4757
timestamp 0
transform 0 1 2544 -1 0 2533
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4756
timestamp 0
transform 0 1 2544 -1 0 2532
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4755
timestamp 0
transform 0 1 2544 -1 0 2531
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4754
timestamp 0
transform 0 1 2544 -1 0 2530
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4753
timestamp 0
transform 0 1 2544 -1 0 2529
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4752
timestamp 0
transform 0 1 2544 -1 0 2528
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4751
timestamp 0
transform 0 1 2544 -1 0 2527
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4750
timestamp 0
transform 0 1 2544 -1 0 2526
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4749
timestamp 0
transform 0 1 2544 -1 0 2525
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4748
timestamp 0
transform 0 1 2544 -1 0 2524
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4747
timestamp 0
transform 0 1 2544 -1 0 2523
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4746
timestamp 0
transform 0 1 2544 -1 0 2522
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4745
timestamp 0
transform 0 1 2544 -1 0 2521
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4744
timestamp 0
transform 0 1 2544 -1 0 2520
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4743
timestamp 0
transform 0 1 2544 -1 0 2519
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4742
timestamp 0
transform 0 1 2544 -1 0 2518
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4741
timestamp 0
transform 0 1 2544 -1 0 2517
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4740
timestamp 0
transform 0 1 2544 -1 0 2516
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4739
timestamp 0
transform 0 1 2544 -1 0 2515
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4738
timestamp 0
transform 0 1 2544 -1 0 2514
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4737
timestamp 0
transform 0 1 2544 -1 0 2513
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4736
timestamp 0
transform 0 1 2544 -1 0 2512
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4735
timestamp 0
transform 0 1 2544 -1 0 2511
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4734
timestamp 0
transform 0 1 2544 -1 0 2510
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4733
timestamp 0
transform 0 1 2544 -1 0 2509
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4732
timestamp 0
transform 0 1 2544 -1 0 2508
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4731
timestamp 0
transform 0 1 2544 -1 0 2507
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4730
timestamp 0
transform 0 1 2544 -1 0 2506
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4729
timestamp 0
transform 0 1 2544 -1 0 2505
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4728
timestamp 0
transform 0 1 2544 -1 0 2504
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4727
timestamp 0
transform 0 1 2544 -1 0 2503
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4726
timestamp 0
transform 0 1 2544 -1 0 2502
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4725
timestamp 0
transform 0 1 2544 -1 0 2501
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4724
timestamp 0
transform 0 1 2544 -1 0 2500
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4723
timestamp 0
transform 0 1 2544 -1 0 2499
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4722
timestamp 0
transform 0 1 2544 -1 0 2498
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4721
timestamp 0
transform 0 1 2544 -1 0 2497
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4720
timestamp 0
transform 0 1 2544 -1 0 2496
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4719
timestamp 0
transform 0 1 2544 -1 0 2495
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4718
timestamp 0
transform 0 1 2544 -1 0 2494
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4717
timestamp 0
transform 0 1 2544 -1 0 2493
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4716
timestamp 0
transform 0 1 2544 -1 0 2492
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4715
timestamp 0
transform 0 1 2544 -1 0 2491
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4714
timestamp 0
transform 0 1 2544 -1 0 2490
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4713
timestamp 0
transform 0 1 2544 -1 0 2489
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4712
timestamp 0
transform 0 1 2544 -1 0 2488
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4711
timestamp 0
transform 0 1 2544 -1 0 2487
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4710
timestamp 0
transform 0 1 2544 -1 0 2486
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4709
timestamp 0
transform 0 1 2544 -1 0 2485
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4708
timestamp 0
transform 0 1 2544 -1 0 2484
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4707
timestamp 0
transform 0 1 2544 -1 0 2483
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4706
timestamp 0
transform 0 1 2544 -1 0 2482
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4705
timestamp 0
transform 0 1 2544 -1 0 2481
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4704
timestamp 0
transform 0 1 2544 -1 0 2480
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4703
timestamp 0
transform 0 1 2544 -1 0 2479
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4702
timestamp 0
transform 0 1 2544 -1 0 2478
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4701
timestamp 0
transform 0 1 2544 -1 0 2477
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4700
timestamp 0
transform 0 1 2544 -1 0 2476
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4699
timestamp 0
transform 0 1 2544 -1 0 2475
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4698
timestamp 0
transform 0 1 2544 -1 0 2474
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4697
timestamp 0
transform 0 1 2544 -1 0 2473
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4696
timestamp 0
transform 0 1 2544 -1 0 2472
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4695
timestamp 0
transform 0 1 2544 -1 0 2471
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4694
timestamp 0
transform 0 1 2544 -1 0 2470
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4693
timestamp 0
transform 0 1 2544 -1 0 2469
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4692
timestamp 0
transform 0 1 2544 -1 0 2468
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4691
timestamp 0
transform 0 1 2544 -1 0 2467
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4690
timestamp 0
transform 0 1 2544 -1 0 2466
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4689
timestamp 0
transform 0 1 2544 -1 0 2465
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4688
timestamp 0
transform 0 1 2544 -1 0 2464
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4687
timestamp 0
transform 0 1 2544 -1 0 2463
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4686
timestamp 0
transform 0 1 2544 -1 0 2462
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4685
timestamp 0
transform 0 1 2544 -1 0 2461
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4684
timestamp 0
transform 0 1 2544 -1 0 2460
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4683
timestamp 0
transform 0 1 2544 -1 0 2459
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4682
timestamp 0
transform 0 1 2544 -1 0 2458
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4681
timestamp 0
transform 0 1 2544 -1 0 2457
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4680
timestamp 0
transform 0 1 2544 -1 0 2456
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4679
timestamp 0
transform 0 1 2544 -1 0 2455
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4678
timestamp 0
transform 0 1 2544 -1 0 2454
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4677
timestamp 0
transform 0 1 2544 -1 0 2453
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4676
timestamp 0
transform 0 1 2544 -1 0 2452
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4675
timestamp 0
transform 0 1 2544 -1 0 2451
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4674
timestamp 0
transform 0 1 2544 -1 0 2450
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4673
timestamp 0
transform 0 1 2544 -1 0 2449
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4672
timestamp 0
transform 0 1 2544 -1 0 2448
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4671
timestamp 0
transform 0 1 2544 -1 0 2447
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4670
timestamp 0
transform 0 1 2544 -1 0 2446
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4669
timestamp 0
transform 0 1 2544 -1 0 2445
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4668
timestamp 0
transform 0 1 2544 -1 0 2444
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4667
timestamp 0
transform 0 1 2544 -1 0 2443
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4666
timestamp 0
transform 0 1 2544 -1 0 2442
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4665
timestamp 0
transform 0 1 2544 -1 0 2441
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4664
timestamp 0
transform 0 1 2544 -1 0 2440
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4663
timestamp 0
transform 0 1 2544 -1 0 2439
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4662
timestamp 0
transform 0 1 2544 -1 0 2438
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4661
timestamp 0
transform 0 1 2544 -1 0 2437
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4660
timestamp 0
transform 0 1 2544 -1 0 2436
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4659
timestamp 0
transform 0 1 2544 -1 0 2435
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4658
timestamp 0
transform 0 1 2544 -1 0 2434
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4657
timestamp 0
transform 0 1 2544 -1 0 2433
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4656
timestamp 0
transform 0 1 2544 -1 0 2432
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4655
timestamp 0
transform 0 1 2544 -1 0 2431
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4654
timestamp 0
transform 0 1 2544 -1 0 2430
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4653
timestamp 0
transform 0 1 2544 -1 0 2429
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4652
timestamp 0
transform 0 1 2544 -1 0 2428
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4651
timestamp 0
transform 0 1 2544 -1 0 2427
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4650
timestamp 0
transform 0 1 2544 -1 0 2426
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4649
timestamp 0
transform 0 1 2544 -1 0 2425
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4648
timestamp 0
transform 0 1 2544 -1 0 2424
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4647
timestamp 0
transform 0 1 2544 -1 0 2423
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4646
timestamp 0
transform 0 1 2544 -1 0 2422
box 0 0 1 1
use s8iom0_gpiov2_pad  gpio_pad[11]
timestamp 0
transform 0 1 2544 -1 0 2421
box 0 0 1 1
use s8iom0s8_top_gpio_ovtv2  ser_tx_pad
timestamp 0
transform 0 -1 200 1 0 2352
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3209
timestamp 0
transform 0 -1 198 1 0 2351
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3208
timestamp 0
transform 0 -1 198 1 0 2350
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3207
timestamp 0
transform 0 -1 198 1 0 2349
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3206
timestamp 0
transform 0 -1 198 1 0 2348
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3205
timestamp 0
transform 0 -1 198 1 0 2347
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3204
timestamp 0
transform 0 -1 198 1 0 2346
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3203
timestamp 0
transform 0 -1 198 1 0 2345
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3202
timestamp 0
transform 0 -1 198 1 0 2344
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3201
timestamp 0
transform 0 -1 198 1 0 2343
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3200
timestamp 0
transform 0 -1 198 1 0 2342
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3199
timestamp 0
transform 0 -1 198 1 0 2341
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3198
timestamp 0
transform 0 -1 198 1 0 2340
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3197
timestamp 0
transform 0 -1 198 1 0 2339
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3196
timestamp 0
transform 0 -1 198 1 0 2338
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3195
timestamp 0
transform 0 -1 198 1 0 2337
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3194
timestamp 0
transform 0 -1 198 1 0 2336
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3193
timestamp 0
transform 0 -1 198 1 0 2335
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3192
timestamp 0
transform 0 -1 198 1 0 2334
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3191
timestamp 0
transform 0 -1 198 1 0 2333
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3190
timestamp 0
transform 0 -1 198 1 0 2332
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3189
timestamp 0
transform 0 -1 198 1 0 2331
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3188
timestamp 0
transform 0 -1 198 1 0 2330
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3187
timestamp 0
transform 0 -1 198 1 0 2329
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3186
timestamp 0
transform 0 -1 198 1 0 2328
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3185
timestamp 0
transform 0 -1 198 1 0 2327
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3184
timestamp 0
transform 0 -1 198 1 0 2326
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3183
timestamp 0
transform 0 -1 198 1 0 2325
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3182
timestamp 0
transform 0 -1 198 1 0 2324
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3181
timestamp 0
transform 0 -1 198 1 0 2323
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3180
timestamp 0
transform 0 -1 198 1 0 2322
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3179
timestamp 0
transform 0 -1 198 1 0 2321
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3178
timestamp 0
transform 0 -1 198 1 0 2320
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3177
timestamp 0
transform 0 -1 198 1 0 2319
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3176
timestamp 0
transform 0 -1 198 1 0 2318
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3175
timestamp 0
transform 0 -1 198 1 0 2317
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3174
timestamp 0
transform 0 -1 198 1 0 2316
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3173
timestamp 0
transform 0 -1 198 1 0 2315
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3172
timestamp 0
transform 0 -1 198 1 0 2314
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3171
timestamp 0
transform 0 -1 198 1 0 2313
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3170
timestamp 0
transform 0 -1 198 1 0 2312
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3169
timestamp 0
transform 0 -1 198 1 0 2311
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3168
timestamp 0
transform 0 -1 198 1 0 2310
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3167
timestamp 0
transform 0 -1 198 1 0 2309
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3166
timestamp 0
transform 0 -1 198 1 0 2308
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3165
timestamp 0
transform 0 -1 198 1 0 2307
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3164
timestamp 0
transform 0 -1 198 1 0 2306
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3163
timestamp 0
transform 0 -1 198 1 0 2305
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3162
timestamp 0
transform 0 -1 198 1 0 2304
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3161
timestamp 0
transform 0 -1 198 1 0 2303
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3160
timestamp 0
transform 0 -1 198 1 0 2302
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3159
timestamp 0
transform 0 -1 198 1 0 2301
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3158
timestamp 0
transform 0 -1 198 1 0 2300
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3157
timestamp 0
transform 0 -1 198 1 0 2299
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3156
timestamp 0
transform 0 -1 198 1 0 2298
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3155
timestamp 0
transform 0 -1 198 1 0 2297
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3154
timestamp 0
transform 0 -1 198 1 0 2296
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3153
timestamp 0
transform 0 -1 198 1 0 2295
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4644
timestamp 0
transform 0 1 2544 -1 0 2341
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4643
timestamp 0
transform 0 1 2544 -1 0 2340
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4642
timestamp 0
transform 0 1 2544 -1 0 2339
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4641
timestamp 0
transform 0 1 2544 -1 0 2338
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4640
timestamp 0
transform 0 1 2544 -1 0 2337
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4639
timestamp 0
transform 0 1 2544 -1 0 2336
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4638
timestamp 0
transform 0 1 2544 -1 0 2335
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4637
timestamp 0
transform 0 1 2544 -1 0 2334
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4636
timestamp 0
transform 0 1 2544 -1 0 2333
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4635
timestamp 0
transform 0 1 2544 -1 0 2332
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4634
timestamp 0
transform 0 1 2544 -1 0 2331
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4633
timestamp 0
transform 0 1 2544 -1 0 2330
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4632
timestamp 0
transform 0 1 2544 -1 0 2329
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4631
timestamp 0
transform 0 1 2544 -1 0 2328
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4630
timestamp 0
transform 0 1 2544 -1 0 2327
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4629
timestamp 0
transform 0 1 2544 -1 0 2326
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4628
timestamp 0
transform 0 1 2544 -1 0 2325
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4627
timestamp 0
transform 0 1 2544 -1 0 2324
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4626
timestamp 0
transform 0 1 2544 -1 0 2323
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4625
timestamp 0
transform 0 1 2544 -1 0 2322
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4624
timestamp 0
transform 0 1 2544 -1 0 2321
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4623
timestamp 0
transform 0 1 2544 -1 0 2320
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4622
timestamp 0
transform 0 1 2544 -1 0 2319
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4621
timestamp 0
transform 0 1 2544 -1 0 2318
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4620
timestamp 0
transform 0 1 2544 -1 0 2317
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4619
timestamp 0
transform 0 1 2544 -1 0 2316
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4618
timestamp 0
transform 0 1 2544 -1 0 2315
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4617
timestamp 0
transform 0 1 2544 -1 0 2314
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4616
timestamp 0
transform 0 1 2544 -1 0 2313
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4615
timestamp 0
transform 0 1 2544 -1 0 2312
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4614
timestamp 0
transform 0 1 2544 -1 0 2311
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4613
timestamp 0
transform 0 1 2544 -1 0 2310
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4612
timestamp 0
transform 0 1 2544 -1 0 2309
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4611
timestamp 0
transform 0 1 2544 -1 0 2308
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4610
timestamp 0
transform 0 1 2544 -1 0 2307
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4609
timestamp 0
transform 0 1 2544 -1 0 2306
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4608
timestamp 0
transform 0 1 2544 -1 0 2305
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4607
timestamp 0
transform 0 1 2544 -1 0 2304
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4606
timestamp 0
transform 0 1 2544 -1 0 2303
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4605
timestamp 0
transform 0 1 2544 -1 0 2302
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4604
timestamp 0
transform 0 1 2544 -1 0 2301
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4603
timestamp 0
transform 0 1 2544 -1 0 2300
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4602
timestamp 0
transform 0 1 2544 -1 0 2299
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4601
timestamp 0
transform 0 1 2544 -1 0 2298
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4600
timestamp 0
transform 0 1 2544 -1 0 2297
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4599
timestamp 0
transform 0 1 2544 -1 0 2296
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4598
timestamp 0
transform 0 1 2544 -1 0 2295
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4597
timestamp 0
transform 0 1 2544 -1 0 2294
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4596
timestamp 0
transform 0 1 2544 -1 0 2293
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4595
timestamp 0
transform 0 1 2544 -1 0 2292
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4594
timestamp 0
transform 0 1 2544 -1 0 2291
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4593
timestamp 0
transform 0 1 2544 -1 0 2290
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4592
timestamp 0
transform 0 1 2544 -1 0 2289
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4591
timestamp 0
transform 0 1 2544 -1 0 2288
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4590
timestamp 0
transform 0 1 2544 -1 0 2287
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4589
timestamp 0
transform 0 1 2544 -1 0 2286
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4588
timestamp 0
transform 0 1 2544 -1 0 2285
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4587
timestamp 0
transform 0 1 2544 -1 0 2284
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4586
timestamp 0
transform 0 1 2544 -1 0 2283
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4585
timestamp 0
transform 0 1 2544 -1 0 2282
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4584
timestamp 0
transform 0 1 2544 -1 0 2281
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4583
timestamp 0
transform 0 1 2544 -1 0 2280
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4582
timestamp 0
transform 0 1 2544 -1 0 2279
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4581
timestamp 0
transform 0 1 2544 -1 0 2278
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4580
timestamp 0
transform 0 1 2544 -1 0 2277
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4579
timestamp 0
transform 0 1 2544 -1 0 2276
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4578
timestamp 0
transform 0 1 2544 -1 0 2275
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4577
timestamp 0
transform 0 1 2544 -1 0 2274
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4576
timestamp 0
transform 0 1 2544 -1 0 2273
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4575
timestamp 0
transform 0 1 2544 -1 0 2272
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4574
timestamp 0
transform 0 1 2544 -1 0 2271
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4573
timestamp 0
transform 0 1 2544 -1 0 2270
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4572
timestamp 0
transform 0 1 2544 -1 0 2269
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4571
timestamp 0
transform 0 1 2544 -1 0 2268
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4570
timestamp 0
transform 0 1 2544 -1 0 2267
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4569
timestamp 0
transform 0 1 2544 -1 0 2266
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4568
timestamp 0
transform 0 1 2544 -1 0 2265
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4567
timestamp 0
transform 0 1 2544 -1 0 2264
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4566
timestamp 0
transform 0 1 2544 -1 0 2263
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4565
timestamp 0
transform 0 1 2544 -1 0 2262
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4564
timestamp 0
transform 0 1 2544 -1 0 2261
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4563
timestamp 0
transform 0 1 2544 -1 0 2260
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4562
timestamp 0
transform 0 1 2544 -1 0 2259
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4561
timestamp 0
transform 0 1 2544 -1 0 2258
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4560
timestamp 0
transform 0 1 2544 -1 0 2257
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4559
timestamp 0
transform 0 1 2544 -1 0 2256
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4558
timestamp 0
transform 0 1 2544 -1 0 2255
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4557
timestamp 0
transform 0 1 2544 -1 0 2254
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4556
timestamp 0
transform 0 1 2544 -1 0 2253
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4555
timestamp 0
transform 0 1 2544 -1 0 2252
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4554
timestamp 0
transform 0 1 2544 -1 0 2251
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4553
timestamp 0
transform 0 1 2544 -1 0 2250
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4552
timestamp 0
transform 0 1 2544 -1 0 2249
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4551
timestamp 0
transform 0 1 2544 -1 0 2248
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4550
timestamp 0
transform 0 1 2544 -1 0 2247
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4549
timestamp 0
transform 0 1 2544 -1 0 2246
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4548
timestamp 0
transform 0 1 2544 -1 0 2245
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4547
timestamp 0
transform 0 1 2544 -1 0 2244
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4546
timestamp 0
transform 0 1 2544 -1 0 2243
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4545
timestamp 0
transform 0 1 2544 -1 0 2242
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4544
timestamp 0
transform 0 1 2544 -1 0 2241
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4543
timestamp 0
transform 0 1 2544 -1 0 2240
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4542
timestamp 0
transform 0 1 2544 -1 0 2239
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4541
timestamp 0
transform 0 1 2544 -1 0 2238
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4540
timestamp 0
transform 0 1 2544 -1 0 2237
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4539
timestamp 0
transform 0 1 2544 -1 0 2236
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4538
timestamp 0
transform 0 1 2544 -1 0 2235
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4537
timestamp 0
transform 0 1 2544 -1 0 2234
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4536
timestamp 0
transform 0 1 2544 -1 0 2233
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4535
timestamp 0
transform 0 1 2544 -1 0 2232
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4534
timestamp 0
transform 0 1 2544 -1 0 2231
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4533
timestamp 0
transform 0 1 2544 -1 0 2230
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4532
timestamp 0
transform 0 1 2544 -1 0 2229
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4531
timestamp 0
transform 0 1 2544 -1 0 2228
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4530
timestamp 0
transform 0 1 2544 -1 0 2227
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4529
timestamp 0
transform 0 1 2544 -1 0 2226
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4528
timestamp 0
transform 0 1 2544 -1 0 2225
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4527
timestamp 0
transform 0 1 2544 -1 0 2224
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4526
timestamp 0
transform 0 1 2544 -1 0 2223
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4525
timestamp 0
transform 0 1 2544 -1 0 2222
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4524
timestamp 0
transform 0 1 2544 -1 0 2221
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4523
timestamp 0
transform 0 1 2544 -1 0 2220
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4522
timestamp 0
transform 0 1 2544 -1 0 2219
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4521
timestamp 0
transform 0 1 2544 -1 0 2218
box 0 0 1 1
use s8iom0_gpiov2_pad  gpio_pad[0]
timestamp 0
transform 0 1 2544 -1 0 2217
box 0 0 1 1
use s8iom0s8_top_gpio_ovtv2  ser_rx_pad
timestamp 0
transform 0 -1 200 1 0 2155
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3151
timestamp 0
transform 0 -1 198 1 0 2154
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3150
timestamp 0
transform 0 -1 198 1 0 2153
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3149
timestamp 0
transform 0 -1 198 1 0 2152
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3148
timestamp 0
transform 0 -1 198 1 0 2151
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3147
timestamp 0
transform 0 -1 198 1 0 2150
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3146
timestamp 0
transform 0 -1 198 1 0 2149
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3145
timestamp 0
transform 0 -1 198 1 0 2148
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3144
timestamp 0
transform 0 -1 198 1 0 2147
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3143
timestamp 0
transform 0 -1 198 1 0 2146
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3142
timestamp 0
transform 0 -1 198 1 0 2145
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3141
timestamp 0
transform 0 -1 198 1 0 2144
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3140
timestamp 0
transform 0 -1 198 1 0 2143
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3139
timestamp 0
transform 0 -1 198 1 0 2142
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3138
timestamp 0
transform 0 -1 198 1 0 2141
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3137
timestamp 0
transform 0 -1 198 1 0 2140
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3136
timestamp 0
transform 0 -1 198 1 0 2139
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3135
timestamp 0
transform 0 -1 198 1 0 2138
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3134
timestamp 0
transform 0 -1 198 1 0 2137
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3133
timestamp 0
transform 0 -1 198 1 0 2136
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3132
timestamp 0
transform 0 -1 198 1 0 2135
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3131
timestamp 0
transform 0 -1 198 1 0 2134
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3130
timestamp 0
transform 0 -1 198 1 0 2133
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3129
timestamp 0
transform 0 -1 198 1 0 2132
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3128
timestamp 0
transform 0 -1 198 1 0 2131
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3127
timestamp 0
transform 0 -1 198 1 0 2130
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3126
timestamp 0
transform 0 -1 198 1 0 2129
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3125
timestamp 0
transform 0 -1 198 1 0 2128
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3124
timestamp 0
transform 0 -1 198 1 0 2127
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3123
timestamp 0
transform 0 -1 198 1 0 2126
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3122
timestamp 0
transform 0 -1 198 1 0 2125
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3121
timestamp 0
transform 0 -1 198 1 0 2124
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3120
timestamp 0
transform 0 -1 198 1 0 2123
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3119
timestamp 0
transform 0 -1 198 1 0 2122
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3118
timestamp 0
transform 0 -1 198 1 0 2121
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3117
timestamp 0
transform 0 -1 198 1 0 2120
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3116
timestamp 0
transform 0 -1 198 1 0 2119
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3115
timestamp 0
transform 0 -1 198 1 0 2118
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3114
timestamp 0
transform 0 -1 198 1 0 2117
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3113
timestamp 0
transform 0 -1 198 1 0 2116
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3112
timestamp 0
transform 0 -1 198 1 0 2115
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3111
timestamp 0
transform 0 -1 198 1 0 2114
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3110
timestamp 0
transform 0 -1 198 1 0 2113
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3109
timestamp 0
transform 0 -1 198 1 0 2112
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3108
timestamp 0
transform 0 -1 198 1 0 2111
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3107
timestamp 0
transform 0 -1 198 1 0 2110
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3106
timestamp 0
transform 0 -1 198 1 0 2109
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3105
timestamp 0
transform 0 -1 198 1 0 2108
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3104
timestamp 0
transform 0 -1 198 1 0 2107
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3103
timestamp 0
transform 0 -1 198 1 0 2106
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3102
timestamp 0
transform 0 -1 198 1 0 2105
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3101
timestamp 0
transform 0 -1 198 1 0 2104
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3100
timestamp 0
transform 0 -1 198 1 0 2103
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3099
timestamp 0
transform 0 -1 198 1 0 2102
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3098
timestamp 0
transform 0 -1 198 1 0 2101
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3097
timestamp 0
transform 0 -1 198 1 0 2100
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3096
timestamp 0
transform 0 -1 198 1 0 2099
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3095
timestamp 0
transform 0 -1 198 1 0 2098
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4519
timestamp 0
transform 0 1 2544 -1 0 2137
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4518
timestamp 0
transform 0 1 2544 -1 0 2136
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4517
timestamp 0
transform 0 1 2544 -1 0 2135
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4516
timestamp 0
transform 0 1 2544 -1 0 2134
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4515
timestamp 0
transform 0 1 2544 -1 0 2133
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4514
timestamp 0
transform 0 1 2544 -1 0 2132
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4513
timestamp 0
transform 0 1 2544 -1 0 2131
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4512
timestamp 0
transform 0 1 2544 -1 0 2130
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4511
timestamp 0
transform 0 1 2544 -1 0 2129
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4510
timestamp 0
transform 0 1 2544 -1 0 2128
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4509
timestamp 0
transform 0 1 2544 -1 0 2127
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4508
timestamp 0
transform 0 1 2544 -1 0 2126
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4507
timestamp 0
transform 0 1 2544 -1 0 2125
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4506
timestamp 0
transform 0 1 2544 -1 0 2124
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4505
timestamp 0
transform 0 1 2544 -1 0 2123
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4504
timestamp 0
transform 0 1 2544 -1 0 2122
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4503
timestamp 0
transform 0 1 2544 -1 0 2121
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4502
timestamp 0
transform 0 1 2544 -1 0 2120
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4501
timestamp 0
transform 0 1 2544 -1 0 2119
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4500
timestamp 0
transform 0 1 2544 -1 0 2118
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4499
timestamp 0
transform 0 1 2544 -1 0 2117
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4498
timestamp 0
transform 0 1 2544 -1 0 2116
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4497
timestamp 0
transform 0 1 2544 -1 0 2115
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4496
timestamp 0
transform 0 1 2544 -1 0 2114
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4495
timestamp 0
transform 0 1 2544 -1 0 2113
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4494
timestamp 0
transform 0 1 2544 -1 0 2112
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4493
timestamp 0
transform 0 1 2544 -1 0 2111
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4492
timestamp 0
transform 0 1 2544 -1 0 2110
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4491
timestamp 0
transform 0 1 2544 -1 0 2109
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4490
timestamp 0
transform 0 1 2544 -1 0 2108
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4489
timestamp 0
transform 0 1 2544 -1 0 2107
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4488
timestamp 0
transform 0 1 2544 -1 0 2106
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4487
timestamp 0
transform 0 1 2544 -1 0 2105
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4486
timestamp 0
transform 0 1 2544 -1 0 2104
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4485
timestamp 0
transform 0 1 2544 -1 0 2103
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4484
timestamp 0
transform 0 1 2544 -1 0 2102
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4483
timestamp 0
transform 0 1 2544 -1 0 2101
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4482
timestamp 0
transform 0 1 2544 -1 0 2100
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4481
timestamp 0
transform 0 1 2544 -1 0 2099
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4480
timestamp 0
transform 0 1 2544 -1 0 2098
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4479
timestamp 0
transform 0 1 2544 -1 0 2097
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4478
timestamp 0
transform 0 1 2544 -1 0 2096
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4477
timestamp 0
transform 0 1 2544 -1 0 2095
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4476
timestamp 0
transform 0 1 2544 -1 0 2094
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4475
timestamp 0
transform 0 1 2544 -1 0 2093
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4474
timestamp 0
transform 0 1 2544 -1 0 2092
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4473
timestamp 0
transform 0 1 2544 -1 0 2091
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4472
timestamp 0
transform 0 1 2544 -1 0 2090
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4471
timestamp 0
transform 0 1 2544 -1 0 2089
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4470
timestamp 0
transform 0 1 2544 -1 0 2088
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4469
timestamp 0
transform 0 1 2544 -1 0 2087
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4468
timestamp 0
transform 0 1 2544 -1 0 2086
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4467
timestamp 0
transform 0 1 2544 -1 0 2085
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4466
timestamp 0
transform 0 1 2544 -1 0 2084
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4465
timestamp 0
transform 0 1 2544 -1 0 2083
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4464
timestamp 0
transform 0 1 2544 -1 0 2082
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4463
timestamp 0
transform 0 1 2544 -1 0 2081
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4462
timestamp 0
transform 0 1 2544 -1 0 2080
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4461
timestamp 0
transform 0 1 2544 -1 0 2079
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4460
timestamp 0
transform 0 1 2544 -1 0 2078
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4459
timestamp 0
transform 0 1 2544 -1 0 2077
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4458
timestamp 0
transform 0 1 2544 -1 0 2076
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4457
timestamp 0
transform 0 1 2544 -1 0 2075
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4456
timestamp 0
transform 0 1 2544 -1 0 2074
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4455
timestamp 0
transform 0 1 2544 -1 0 2073
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4454
timestamp 0
transform 0 1 2544 -1 0 2072
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4453
timestamp 0
transform 0 1 2544 -1 0 2071
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4452
timestamp 0
transform 0 1 2544 -1 0 2070
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4451
timestamp 0
transform 0 1 2544 -1 0 2069
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4450
timestamp 0
transform 0 1 2544 -1 0 2068
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4449
timestamp 0
transform 0 1 2544 -1 0 2067
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4448
timestamp 0
transform 0 1 2544 -1 0 2066
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4447
timestamp 0
transform 0 1 2544 -1 0 2065
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4446
timestamp 0
transform 0 1 2544 -1 0 2064
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4445
timestamp 0
transform 0 1 2544 -1 0 2063
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4444
timestamp 0
transform 0 1 2544 -1 0 2062
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4443
timestamp 0
transform 0 1 2544 -1 0 2061
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4442
timestamp 0
transform 0 1 2544 -1 0 2060
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4441
timestamp 0
transform 0 1 2544 -1 0 2059
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4440
timestamp 0
transform 0 1 2544 -1 0 2058
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4439
timestamp 0
transform 0 1 2544 -1 0 2057
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4438
timestamp 0
transform 0 1 2544 -1 0 2056
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4437
timestamp 0
transform 0 1 2544 -1 0 2055
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4436
timestamp 0
transform 0 1 2544 -1 0 2054
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4435
timestamp 0
transform 0 1 2544 -1 0 2053
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4434
timestamp 0
transform 0 1 2544 -1 0 2052
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4433
timestamp 0
transform 0 1 2544 -1 0 2051
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4432
timestamp 0
transform 0 1 2544 -1 0 2050
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4431
timestamp 0
transform 0 1 2544 -1 0 2049
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4430
timestamp 0
transform 0 1 2544 -1 0 2048
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4429
timestamp 0
transform 0 1 2544 -1 0 2047
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4428
timestamp 0
transform 0 1 2544 -1 0 2046
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4427
timestamp 0
transform 0 1 2544 -1 0 2045
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4426
timestamp 0
transform 0 1 2544 -1 0 2044
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4425
timestamp 0
transform 0 1 2544 -1 0 2043
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4424
timestamp 0
transform 0 1 2544 -1 0 2042
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4423
timestamp 0
transform 0 1 2544 -1 0 2041
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4422
timestamp 0
transform 0 1 2544 -1 0 2040
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4421
timestamp 0
transform 0 1 2544 -1 0 2039
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4420
timestamp 0
transform 0 1 2544 -1 0 2038
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4419
timestamp 0
transform 0 1 2544 -1 0 2037
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4418
timestamp 0
transform 0 1 2544 -1 0 2036
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4417
timestamp 0
transform 0 1 2544 -1 0 2035
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4416
timestamp 0
transform 0 1 2544 -1 0 2034
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4415
timestamp 0
transform 0 1 2544 -1 0 2033
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4414
timestamp 0
transform 0 1 2544 -1 0 2032
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4413
timestamp 0
transform 0 1 2544 -1 0 2031
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4412
timestamp 0
transform 0 1 2544 -1 0 2030
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4411
timestamp 0
transform 0 1 2544 -1 0 2029
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4410
timestamp 0
transform 0 1 2544 -1 0 2028
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4409
timestamp 0
transform 0 1 2544 -1 0 2027
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4408
timestamp 0
transform 0 1 2544 -1 0 2026
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4407
timestamp 0
transform 0 1 2544 -1 0 2025
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4406
timestamp 0
transform 0 1 2544 -1 0 2024
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4405
timestamp 0
transform 0 1 2544 -1 0 2023
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4404
timestamp 0
transform 0 1 2544 -1 0 2022
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4403
timestamp 0
transform 0 1 2544 -1 0 2021
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4402
timestamp 0
transform 0 1 2544 -1 0 2020
box 0 0 1 1
use s8iom0_gpiov2_pad  flash_io3_pad
timestamp 0
transform 0 -1 198 1 0 2018
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3093
timestamp 0
transform 0 -1 198 1 0 2017
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3092
timestamp 0
transform 0 -1 198 1 0 2016
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3091
timestamp 0
transform 0 -1 198 1 0 2015
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3090
timestamp 0
transform 0 -1 198 1 0 2014
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3089
timestamp 0
transform 0 -1 198 1 0 2013
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3088
timestamp 0
transform 0 -1 198 1 0 2012
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4401
timestamp 0
transform 0 1 2544 -1 0 2019
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4400
timestamp 0
transform 0 1 2544 -1 0 2018
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4399
timestamp 0
transform 0 1 2544 -1 0 2017
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4398
timestamp 0
transform 0 1 2544 -1 0 2016
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4397
timestamp 0
transform 0 1 2544 -1 0 2015
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4396
timestamp 0
transform 0 1 2544 -1 0 2014
box 0 0 1 1
use s8iom0_gpiov2_pad  gpio_pad[1]
timestamp 0
transform 0 1 2544 -1 0 2013
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3087
timestamp 0
transform 0 -1 198 1 0 2011
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3086
timestamp 0
transform 0 -1 198 1 0 2010
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3085
timestamp 0
transform 0 -1 198 1 0 2009
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3084
timestamp 0
transform 0 -1 198 1 0 2008
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3083
timestamp 0
transform 0 -1 198 1 0 2007
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3082
timestamp 0
transform 0 -1 198 1 0 2006
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3081
timestamp 0
transform 0 -1 198 1 0 2005
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3080
timestamp 0
transform 0 -1 198 1 0 2004
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3079
timestamp 0
transform 0 -1 198 1 0 2003
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3078
timestamp 0
transform 0 -1 198 1 0 2002
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3077
timestamp 0
transform 0 -1 198 1 0 2001
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3076
timestamp 0
transform 0 -1 198 1 0 2000
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3075
timestamp 0
transform 0 -1 198 1 0 1999
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3074
timestamp 0
transform 0 -1 198 1 0 1998
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3073
timestamp 0
transform 0 -1 198 1 0 1997
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3072
timestamp 0
transform 0 -1 198 1 0 1996
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3071
timestamp 0
transform 0 -1 198 1 0 1995
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3070
timestamp 0
transform 0 -1 198 1 0 1994
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3069
timestamp 0
transform 0 -1 198 1 0 1993
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3068
timestamp 0
transform 0 -1 198 1 0 1992
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3067
timestamp 0
transform 0 -1 198 1 0 1991
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3066
timestamp 0
transform 0 -1 198 1 0 1990
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3065
timestamp 0
transform 0 -1 198 1 0 1989
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3064
timestamp 0
transform 0 -1 198 1 0 1988
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3063
timestamp 0
transform 0 -1 198 1 0 1987
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3062
timestamp 0
transform 0 -1 198 1 0 1986
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3061
timestamp 0
transform 0 -1 198 1 0 1985
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3060
timestamp 0
transform 0 -1 198 1 0 1984
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3059
timestamp 0
transform 0 -1 198 1 0 1983
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3058
timestamp 0
transform 0 -1 198 1 0 1982
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3057
timestamp 0
transform 0 -1 198 1 0 1981
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3056
timestamp 0
transform 0 -1 198 1 0 1980
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3055
timestamp 0
transform 0 -1 198 1 0 1979
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3054
timestamp 0
transform 0 -1 198 1 0 1978
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3053
timestamp 0
transform 0 -1 198 1 0 1977
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3052
timestamp 0
transform 0 -1 198 1 0 1976
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3051
timestamp 0
transform 0 -1 198 1 0 1975
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3050
timestamp 0
transform 0 -1 198 1 0 1974
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3049
timestamp 0
transform 0 -1 198 1 0 1973
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3048
timestamp 0
transform 0 -1 198 1 0 1972
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3047
timestamp 0
transform 0 -1 198 1 0 1971
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3046
timestamp 0
transform 0 -1 198 1 0 1970
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3045
timestamp 0
transform 0 -1 198 1 0 1969
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3044
timestamp 0
transform 0 -1 198 1 0 1968
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3043
timestamp 0
transform 0 -1 198 1 0 1967
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3042
timestamp 0
transform 0 -1 198 1 0 1966
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3041
timestamp 0
transform 0 -1 198 1 0 1965
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3040
timestamp 0
transform 0 -1 198 1 0 1964
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3039
timestamp 0
transform 0 -1 198 1 0 1963
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3038
timestamp 0
transform 0 -1 198 1 0 1962
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3037
timestamp 0
transform 0 -1 198 1 0 1961
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4394
timestamp 0
transform 0 1 2544 -1 0 1933
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4393
timestamp 0
transform 0 1 2544 -1 0 1932
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4392
timestamp 0
transform 0 1 2544 -1 0 1931
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4391
timestamp 0
transform 0 1 2544 -1 0 1930
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4390
timestamp 0
transform 0 1 2544 -1 0 1929
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4389
timestamp 0
transform 0 1 2544 -1 0 1928
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4388
timestamp 0
transform 0 1 2544 -1 0 1927
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4387
timestamp 0
transform 0 1 2544 -1 0 1926
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4386
timestamp 0
transform 0 1 2544 -1 0 1925
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4385
timestamp 0
transform 0 1 2544 -1 0 1924
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4384
timestamp 0
transform 0 1 2544 -1 0 1923
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4383
timestamp 0
transform 0 1 2544 -1 0 1922
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4382
timestamp 0
transform 0 1 2544 -1 0 1921
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4381
timestamp 0
transform 0 1 2544 -1 0 1920
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4380
timestamp 0
transform 0 1 2544 -1 0 1919
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4379
timestamp 0
transform 0 1 2544 -1 0 1918
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4378
timestamp 0
transform 0 1 2544 -1 0 1917
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4377
timestamp 0
transform 0 1 2544 -1 0 1916
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4376
timestamp 0
transform 0 1 2544 -1 0 1915
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4375
timestamp 0
transform 0 1 2544 -1 0 1914
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4374
timestamp 0
transform 0 1 2544 -1 0 1913
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4373
timestamp 0
transform 0 1 2544 -1 0 1912
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4372
timestamp 0
transform 0 1 2544 -1 0 1911
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4371
timestamp 0
transform 0 1 2544 -1 0 1910
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4370
timestamp 0
transform 0 1 2544 -1 0 1909
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4369
timestamp 0
transform 0 1 2544 -1 0 1908
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4368
timestamp 0
transform 0 1 2544 -1 0 1907
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4367
timestamp 0
transform 0 1 2544 -1 0 1906
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4366
timestamp 0
transform 0 1 2544 -1 0 1905
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4365
timestamp 0
transform 0 1 2544 -1 0 1904
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4364
timestamp 0
transform 0 1 2544 -1 0 1903
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4363
timestamp 0
transform 0 1 2544 -1 0 1902
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4362
timestamp 0
transform 0 1 2544 -1 0 1901
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4361
timestamp 0
transform 0 1 2544 -1 0 1900
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4360
timestamp 0
transform 0 1 2544 -1 0 1899
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4359
timestamp 0
transform 0 1 2544 -1 0 1898
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4358
timestamp 0
transform 0 1 2544 -1 0 1897
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4357
timestamp 0
transform 0 1 2544 -1 0 1896
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4356
timestamp 0
transform 0 1 2544 -1 0 1895
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4355
timestamp 0
transform 0 1 2544 -1 0 1894
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4354
timestamp 0
transform 0 1 2544 -1 0 1893
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4353
timestamp 0
transform 0 1 2544 -1 0 1892
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4352
timestamp 0
transform 0 1 2544 -1 0 1891
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4351
timestamp 0
transform 0 1 2544 -1 0 1890
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4350
timestamp 0
transform 0 1 2544 -1 0 1889
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4349
timestamp 0
transform 0 1 2544 -1 0 1888
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4348
timestamp 0
transform 0 1 2544 -1 0 1887
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4347
timestamp 0
transform 0 1 2544 -1 0 1886
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4346
timestamp 0
transform 0 1 2544 -1 0 1885
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4345
timestamp 0
transform 0 1 2544 -1 0 1884
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4344
timestamp 0
transform 0 1 2544 -1 0 1883
box 0 0 1 1
use s8iom0_gpiov2_pad  flash_io2_pad
timestamp 0
transform 0 -1 198 1 0 1881
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3035
timestamp 0
transform 0 -1 198 1 0 1880
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3034
timestamp 0
transform 0 -1 198 1 0 1879
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3033
timestamp 0
transform 0 -1 198 1 0 1878
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3032
timestamp 0
transform 0 -1 198 1 0 1877
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3031
timestamp 0
transform 0 -1 198 1 0 1876
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3030
timestamp 0
transform 0 -1 198 1 0 1875
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3029
timestamp 0
transform 0 -1 198 1 0 1874
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3028
timestamp 0
transform 0 -1 198 1 0 1873
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3027
timestamp 0
transform 0 -1 198 1 0 1872
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3026
timestamp 0
transform 0 -1 198 1 0 1871
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3025
timestamp 0
transform 0 -1 198 1 0 1870
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3024
timestamp 0
transform 0 -1 198 1 0 1869
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3023
timestamp 0
transform 0 -1 198 1 0 1868
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3022
timestamp 0
transform 0 -1 198 1 0 1867
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3021
timestamp 0
transform 0 -1 198 1 0 1866
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3020
timestamp 0
transform 0 -1 198 1 0 1865
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3019
timestamp 0
transform 0 -1 198 1 0 1864
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3018
timestamp 0
transform 0 -1 198 1 0 1863
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3017
timestamp 0
transform 0 -1 198 1 0 1862
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3016
timestamp 0
transform 0 -1 198 1 0 1861
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3015
timestamp 0
transform 0 -1 198 1 0 1860
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3014
timestamp 0
transform 0 -1 198 1 0 1859
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3013
timestamp 0
transform 0 -1 198 1 0 1858
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3012
timestamp 0
transform 0 -1 198 1 0 1857
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3011
timestamp 0
transform 0 -1 198 1 0 1856
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3010
timestamp 0
transform 0 -1 198 1 0 1855
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3009
timestamp 0
transform 0 -1 198 1 0 1854
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3008
timestamp 0
transform 0 -1 198 1 0 1853
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3007
timestamp 0
transform 0 -1 198 1 0 1852
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3006
timestamp 0
transform 0 -1 198 1 0 1851
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3005
timestamp 0
transform 0 -1 198 1 0 1850
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3004
timestamp 0
transform 0 -1 198 1 0 1849
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3003
timestamp 0
transform 0 -1 198 1 0 1848
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3002
timestamp 0
transform 0 -1 198 1 0 1847
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3001
timestamp 0
transform 0 -1 198 1 0 1846
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3000
timestamp 0
transform 0 -1 198 1 0 1845
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2999
timestamp 0
transform 0 -1 198 1 0 1844
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2998
timestamp 0
transform 0 -1 198 1 0 1843
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2997
timestamp 0
transform 0 -1 198 1 0 1842
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2996
timestamp 0
transform 0 -1 198 1 0 1841
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2995
timestamp 0
transform 0 -1 198 1 0 1840
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2994
timestamp 0
transform 0 -1 198 1 0 1839
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2993
timestamp 0
transform 0 -1 198 1 0 1838
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2992
timestamp 0
transform 0 -1 198 1 0 1837
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2991
timestamp 0
transform 0 -1 198 1 0 1836
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2990
timestamp 0
transform 0 -1 198 1 0 1835
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2989
timestamp 0
transform 0 -1 198 1 0 1834
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2988
timestamp 0
transform 0 -1 198 1 0 1833
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2987
timestamp 0
transform 0 -1 198 1 0 1832
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2986
timestamp 0
transform 0 -1 198 1 0 1831
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2985
timestamp 0
transform 0 -1 198 1 0 1830
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2984
timestamp 0
transform 0 -1 198 1 0 1829
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2983
timestamp 0
transform 0 -1 198 1 0 1828
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2982
timestamp 0
transform 0 -1 198 1 0 1827
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2981
timestamp 0
transform 0 -1 198 1 0 1826
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2980
timestamp 0
transform 0 -1 198 1 0 1825
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2979
timestamp 0
transform 0 -1 198 1 0 1824
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4343
timestamp 0
transform 0 1 2544 -1 0 1882
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4342
timestamp 0
transform 0 1 2544 -1 0 1881
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4341
timestamp 0
transform 0 1 2544 -1 0 1880
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4340
timestamp 0
transform 0 1 2544 -1 0 1879
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4339
timestamp 0
transform 0 1 2544 -1 0 1878
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4338
timestamp 0
transform 0 1 2544 -1 0 1877
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4337
timestamp 0
transform 0 1 2544 -1 0 1876
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4336
timestamp 0
transform 0 1 2544 -1 0 1875
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4335
timestamp 0
transform 0 1 2544 -1 0 1874
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4334
timestamp 0
transform 0 1 2544 -1 0 1873
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4333
timestamp 0
transform 0 1 2544 -1 0 1872
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4332
timestamp 0
transform 0 1 2544 -1 0 1871
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4331
timestamp 0
transform 0 1 2544 -1 0 1870
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4330
timestamp 0
transform 0 1 2544 -1 0 1869
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4329
timestamp 0
transform 0 1 2544 -1 0 1868
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4328
timestamp 0
transform 0 1 2544 -1 0 1867
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4327
timestamp 0
transform 0 1 2544 -1 0 1866
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4326
timestamp 0
transform 0 1 2544 -1 0 1865
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4325
timestamp 0
transform 0 1 2544 -1 0 1864
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4324
timestamp 0
transform 0 1 2544 -1 0 1863
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4323
timestamp 0
transform 0 1 2544 -1 0 1862
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4322
timestamp 0
transform 0 1 2544 -1 0 1861
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4321
timestamp 0
transform 0 1 2544 -1 0 1860
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4320
timestamp 0
transform 0 1 2544 -1 0 1859
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4319
timestamp 0
transform 0 1 2544 -1 0 1858
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4318
timestamp 0
transform 0 1 2544 -1 0 1857
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4317
timestamp 0
transform 0 1 2544 -1 0 1856
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4316
timestamp 0
transform 0 1 2544 -1 0 1855
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4315
timestamp 0
transform 0 1 2544 -1 0 1854
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4314
timestamp 0
transform 0 1 2544 -1 0 1853
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4313
timestamp 0
transform 0 1 2544 -1 0 1852
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4312
timestamp 0
transform 0 1 2544 -1 0 1851
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4311
timestamp 0
transform 0 1 2544 -1 0 1850
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4310
timestamp 0
transform 0 1 2544 -1 0 1849
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4309
timestamp 0
transform 0 1 2544 -1 0 1848
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4308
timestamp 0
transform 0 1 2544 -1 0 1847
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4307
timestamp 0
transform 0 1 2544 -1 0 1846
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4306
timestamp 0
transform 0 1 2544 -1 0 1845
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4305
timestamp 0
transform 0 1 2544 -1 0 1844
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4304
timestamp 0
transform 0 1 2544 -1 0 1843
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4303
timestamp 0
transform 0 1 2544 -1 0 1842
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4302
timestamp 0
transform 0 1 2544 -1 0 1841
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4301
timestamp 0
transform 0 1 2544 -1 0 1840
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4300
timestamp 0
transform 0 1 2544 -1 0 1839
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4299
timestamp 0
transform 0 1 2544 -1 0 1838
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4298
timestamp 0
transform 0 1 2544 -1 0 1837
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4297
timestamp 0
transform 0 1 2544 -1 0 1836
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4296
timestamp 0
transform 0 1 2544 -1 0 1835
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4295
timestamp 0
transform 0 1 2544 -1 0 1834
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4294
timestamp 0
transform 0 1 2544 -1 0 1833
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4293
timestamp 0
transform 0 1 2544 -1 0 1832
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4292
timestamp 0
transform 0 1 2544 -1 0 1831
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4291
timestamp 0
transform 0 1 2544 -1 0 1830
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4290
timestamp 0
transform 0 1 2544 -1 0 1829
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4289
timestamp 0
transform 0 1 2544 -1 0 1828
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4288
timestamp 0
transform 0 1 2544 -1 0 1827
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4287
timestamp 0
transform 0 1 2544 -1 0 1826
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4286
timestamp 0
transform 0 1 2544 -1 0 1825
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4285
timestamp 0
transform 0 1 2544 -1 0 1824
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4284
timestamp 0
transform 0 1 2544 -1 0 1823
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4283
timestamp 0
transform 0 1 2544 -1 0 1822
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4282
timestamp 0
transform 0 1 2544 -1 0 1821
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4281
timestamp 0
transform 0 1 2544 -1 0 1820
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4280
timestamp 0
transform 0 1 2544 -1 0 1819
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4279
timestamp 0
transform 0 1 2544 -1 0 1818
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4278
timestamp 0
transform 0 1 2544 -1 0 1817
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4277
timestamp 0
transform 0 1 2544 -1 0 1816
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4276
timestamp 0
transform 0 1 2544 -1 0 1815
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4275
timestamp 0
transform 0 1 2544 -1 0 1814
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4274
timestamp 0
transform 0 1 2544 -1 0 1813
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4273
timestamp 0
transform 0 1 2544 -1 0 1812
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4272
timestamp 0
transform 0 1 2544 -1 0 1811
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4271
timestamp 0
transform 0 1 2544 -1 0 1810
box 0 0 1 1
use s8iom0_gpiov2_pad  gpio_pad[2]
timestamp 0
transform 0 1 2544 -1 0 1809
box 0 0 1 1
use s8iom0_gpiov2_pad  flash_io1_pad
timestamp 0
transform 0 -1 198 1 0 1744
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2977
timestamp 0
transform 0 -1 198 1 0 1743
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2976
timestamp 0
transform 0 -1 198 1 0 1742
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2975
timestamp 0
transform 0 -1 198 1 0 1741
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2974
timestamp 0
transform 0 -1 198 1 0 1740
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2973
timestamp 0
transform 0 -1 198 1 0 1739
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2972
timestamp 0
transform 0 -1 198 1 0 1738
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2971
timestamp 0
transform 0 -1 198 1 0 1737
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2970
timestamp 0
transform 0 -1 198 1 0 1736
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2969
timestamp 0
transform 0 -1 198 1 0 1735
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2968
timestamp 0
transform 0 -1 198 1 0 1734
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2967
timestamp 0
transform 0 -1 198 1 0 1733
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2966
timestamp 0
transform 0 -1 198 1 0 1732
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2965
timestamp 0
transform 0 -1 198 1 0 1731
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2964
timestamp 0
transform 0 -1 198 1 0 1730
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2963
timestamp 0
transform 0 -1 198 1 0 1729
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2962
timestamp 0
transform 0 -1 198 1 0 1728
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2961
timestamp 0
transform 0 -1 198 1 0 1727
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2960
timestamp 0
transform 0 -1 198 1 0 1726
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2959
timestamp 0
transform 0 -1 198 1 0 1725
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2958
timestamp 0
transform 0 -1 198 1 0 1724
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2957
timestamp 0
transform 0 -1 198 1 0 1723
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2956
timestamp 0
transform 0 -1 198 1 0 1722
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2955
timestamp 0
transform 0 -1 198 1 0 1721
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2954
timestamp 0
transform 0 -1 198 1 0 1720
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2953
timestamp 0
transform 0 -1 198 1 0 1719
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2952
timestamp 0
transform 0 -1 198 1 0 1718
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2951
timestamp 0
transform 0 -1 198 1 0 1717
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2950
timestamp 0
transform 0 -1 198 1 0 1716
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2949
timestamp 0
transform 0 -1 198 1 0 1715
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2948
timestamp 0
transform 0 -1 198 1 0 1714
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2947
timestamp 0
transform 0 -1 198 1 0 1713
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2946
timestamp 0
transform 0 -1 198 1 0 1712
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2945
timestamp 0
transform 0 -1 198 1 0 1711
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2944
timestamp 0
transform 0 -1 198 1 0 1710
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2943
timestamp 0
transform 0 -1 198 1 0 1709
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2942
timestamp 0
transform 0 -1 198 1 0 1708
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2941
timestamp 0
transform 0 -1 198 1 0 1707
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2940
timestamp 0
transform 0 -1 198 1 0 1706
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2939
timestamp 0
transform 0 -1 198 1 0 1705
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2938
timestamp 0
transform 0 -1 198 1 0 1704
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2937
timestamp 0
transform 0 -1 198 1 0 1703
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2936
timestamp 0
transform 0 -1 198 1 0 1702
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2935
timestamp 0
transform 0 -1 198 1 0 1701
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2934
timestamp 0
transform 0 -1 198 1 0 1700
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2933
timestamp 0
transform 0 -1 198 1 0 1699
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2932
timestamp 0
transform 0 -1 198 1 0 1698
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2931
timestamp 0
transform 0 -1 198 1 0 1697
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2930
timestamp 0
transform 0 -1 198 1 0 1696
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2929
timestamp 0
transform 0 -1 198 1 0 1695
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2928
timestamp 0
transform 0 -1 198 1 0 1694
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2927
timestamp 0
transform 0 -1 198 1 0 1693
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2926
timestamp 0
transform 0 -1 198 1 0 1692
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2925
timestamp 0
transform 0 -1 198 1 0 1691
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2924
timestamp 0
transform 0 -1 198 1 0 1690
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2923
timestamp 0
transform 0 -1 198 1 0 1689
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2922
timestamp 0
transform 0 -1 198 1 0 1688
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2921
timestamp 0
transform 0 -1 198 1 0 1687
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4269
timestamp 0
transform 0 1 2544 -1 0 1729
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4268
timestamp 0
transform 0 1 2544 -1 0 1728
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4267
timestamp 0
transform 0 1 2544 -1 0 1727
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4266
timestamp 0
transform 0 1 2544 -1 0 1726
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4265
timestamp 0
transform 0 1 2544 -1 0 1725
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4264
timestamp 0
transform 0 1 2544 -1 0 1724
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4263
timestamp 0
transform 0 1 2544 -1 0 1723
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4262
timestamp 0
transform 0 1 2544 -1 0 1722
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4261
timestamp 0
transform 0 1 2544 -1 0 1721
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4260
timestamp 0
transform 0 1 2544 -1 0 1720
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4259
timestamp 0
transform 0 1 2544 -1 0 1719
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4258
timestamp 0
transform 0 1 2544 -1 0 1718
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4257
timestamp 0
transform 0 1 2544 -1 0 1717
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4256
timestamp 0
transform 0 1 2544 -1 0 1716
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4255
timestamp 0
transform 0 1 2544 -1 0 1715
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4254
timestamp 0
transform 0 1 2544 -1 0 1714
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4253
timestamp 0
transform 0 1 2544 -1 0 1713
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4252
timestamp 0
transform 0 1 2544 -1 0 1712
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4251
timestamp 0
transform 0 1 2544 -1 0 1711
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4250
timestamp 0
transform 0 1 2544 -1 0 1710
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4249
timestamp 0
transform 0 1 2544 -1 0 1709
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4248
timestamp 0
transform 0 1 2544 -1 0 1708
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4247
timestamp 0
transform 0 1 2544 -1 0 1707
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4246
timestamp 0
transform 0 1 2544 -1 0 1706
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4245
timestamp 0
transform 0 1 2544 -1 0 1705
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4244
timestamp 0
transform 0 1 2544 -1 0 1704
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4243
timestamp 0
transform 0 1 2544 -1 0 1703
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4242
timestamp 0
transform 0 1 2544 -1 0 1702
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4241
timestamp 0
transform 0 1 2544 -1 0 1701
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4240
timestamp 0
transform 0 1 2544 -1 0 1700
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4239
timestamp 0
transform 0 1 2544 -1 0 1699
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4238
timestamp 0
transform 0 1 2544 -1 0 1698
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4237
timestamp 0
transform 0 1 2544 -1 0 1697
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4236
timestamp 0
transform 0 1 2544 -1 0 1696
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4235
timestamp 0
transform 0 1 2544 -1 0 1695
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4234
timestamp 0
transform 0 1 2544 -1 0 1694
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4233
timestamp 0
transform 0 1 2544 -1 0 1693
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4232
timestamp 0
transform 0 1 2544 -1 0 1692
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4231
timestamp 0
transform 0 1 2544 -1 0 1691
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4230
timestamp 0
transform 0 1 2544 -1 0 1690
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4229
timestamp 0
transform 0 1 2544 -1 0 1689
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4228
timestamp 0
transform 0 1 2544 -1 0 1688
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4227
timestamp 0
transform 0 1 2544 -1 0 1687
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4226
timestamp 0
transform 0 1 2544 -1 0 1686
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4225
timestamp 0
transform 0 1 2544 -1 0 1685
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4224
timestamp 0
transform 0 1 2544 -1 0 1684
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4223
timestamp 0
transform 0 1 2544 -1 0 1683
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4222
timestamp 0
transform 0 1 2544 -1 0 1682
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4221
timestamp 0
transform 0 1 2544 -1 0 1681
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4220
timestamp 0
transform 0 1 2544 -1 0 1680
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4219
timestamp 0
transform 0 1 2544 -1 0 1679
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4218
timestamp 0
transform 0 1 2544 -1 0 1678
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4217
timestamp 0
transform 0 1 2544 -1 0 1677
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4216
timestamp 0
transform 0 1 2544 -1 0 1676
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4215
timestamp 0
transform 0 1 2544 -1 0 1675
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4214
timestamp 0
transform 0 1 2544 -1 0 1674
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4213
timestamp 0
transform 0 1 2544 -1 0 1673
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4212
timestamp 0
transform 0 1 2544 -1 0 1672
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4211
timestamp 0
transform 0 1 2544 -1 0 1671
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4210
timestamp 0
transform 0 1 2544 -1 0 1670
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4209
timestamp 0
transform 0 1 2544 -1 0 1669
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4208
timestamp 0
transform 0 1 2544 -1 0 1668
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4207
timestamp 0
transform 0 1 2544 -1 0 1667
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4206
timestamp 0
transform 0 1 2544 -1 0 1666
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4205
timestamp 0
transform 0 1 2544 -1 0 1665
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4204
timestamp 0
transform 0 1 2544 -1 0 1664
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4203
timestamp 0
transform 0 1 2544 -1 0 1663
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4202
timestamp 0
transform 0 1 2544 -1 0 1662
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4201
timestamp 0
transform 0 1 2544 -1 0 1661
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4200
timestamp 0
transform 0 1 2544 -1 0 1660
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4199
timestamp 0
transform 0 1 2544 -1 0 1659
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4198
timestamp 0
transform 0 1 2544 -1 0 1658
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4197
timestamp 0
transform 0 1 2544 -1 0 1657
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4196
timestamp 0
transform 0 1 2544 -1 0 1656
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4195
timestamp 0
transform 0 1 2544 -1 0 1655
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4194
timestamp 0
transform 0 1 2544 -1 0 1654
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4193
timestamp 0
transform 0 1 2544 -1 0 1653
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4192
timestamp 0
transform 0 1 2544 -1 0 1652
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4191
timestamp 0
transform 0 1 2544 -1 0 1651
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4190
timestamp 0
transform 0 1 2544 -1 0 1650
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4189
timestamp 0
transform 0 1 2544 -1 0 1649
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4188
timestamp 0
transform 0 1 2544 -1 0 1648
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4187
timestamp 0
transform 0 1 2544 -1 0 1647
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4186
timestamp 0
transform 0 1 2544 -1 0 1646
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4185
timestamp 0
transform 0 1 2544 -1 0 1645
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4184
timestamp 0
transform 0 1 2544 -1 0 1644
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4183
timestamp 0
transform 0 1 2544 -1 0 1643
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4182
timestamp 0
transform 0 1 2544 -1 0 1642
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4181
timestamp 0
transform 0 1 2544 -1 0 1641
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4180
timestamp 0
transform 0 1 2544 -1 0 1640
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4179
timestamp 0
transform 0 1 2544 -1 0 1639
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4178
timestamp 0
transform 0 1 2544 -1 0 1638
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4177
timestamp 0
transform 0 1 2544 -1 0 1637
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4176
timestamp 0
transform 0 1 2544 -1 0 1636
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4175
timestamp 0
transform 0 1 2544 -1 0 1635
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4174
timestamp 0
transform 0 1 2544 -1 0 1634
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4173
timestamp 0
transform 0 1 2544 -1 0 1633
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4172
timestamp 0
transform 0 1 2544 -1 0 1632
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4171
timestamp 0
transform 0 1 2544 -1 0 1631
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4170
timestamp 0
transform 0 1 2544 -1 0 1630
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4169
timestamp 0
transform 0 1 2544 -1 0 1629
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4168
timestamp 0
transform 0 1 2544 -1 0 1628
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4167
timestamp 0
transform 0 1 2544 -1 0 1627
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4166
timestamp 0
transform 0 1 2544 -1 0 1626
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4165
timestamp 0
transform 0 1 2544 -1 0 1625
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4164
timestamp 0
transform 0 1 2544 -1 0 1624
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4163
timestamp 0
transform 0 1 2544 -1 0 1623
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4162
timestamp 0
transform 0 1 2544 -1 0 1622
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4161
timestamp 0
transform 0 1 2544 -1 0 1621
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4160
timestamp 0
transform 0 1 2544 -1 0 1620
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4159
timestamp 0
transform 0 1 2544 -1 0 1619
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4158
timestamp 0
transform 0 1 2544 -1 0 1618
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4157
timestamp 0
transform 0 1 2544 -1 0 1617
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4156
timestamp 0
transform 0 1 2544 -1 0 1616
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4155
timestamp 0
transform 0 1 2544 -1 0 1615
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4154
timestamp 0
transform 0 1 2544 -1 0 1614
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4153
timestamp 0
transform 0 1 2544 -1 0 1613
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4152
timestamp 0
transform 0 1 2544 -1 0 1612
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4151
timestamp 0
transform 0 1 2544 -1 0 1611
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4150
timestamp 0
transform 0 1 2544 -1 0 1610
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4149
timestamp 0
transform 0 1 2544 -1 0 1609
box 0 0 1 1
use s8iom0_gpiov2_pad  flash_io0_pad
timestamp 0
transform 0 -1 198 1 0 1607
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2919
timestamp 0
transform 0 -1 198 1 0 1606
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2918
timestamp 0
transform 0 -1 198 1 0 1605
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2917
timestamp 0
transform 0 -1 198 1 0 1604
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2916
timestamp 0
transform 0 -1 198 1 0 1603
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4148
timestamp 0
transform 0 1 2544 -1 0 1608
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4147
timestamp 0
transform 0 1 2544 -1 0 1607
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4146
timestamp 0
transform 0 1 2544 -1 0 1606
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4145
timestamp 0
transform 0 1 2544 -1 0 1605
box 0 0 1 1
use s8iom0_gpiov2_pad  gpio_pad[3]
timestamp 0
transform 0 1 2544 -1 0 1604
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2915
timestamp 0
transform 0 -1 198 1 0 1602
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2914
timestamp 0
transform 0 -1 198 1 0 1601
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2913
timestamp 0
transform 0 -1 198 1 0 1600
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2912
timestamp 0
transform 0 -1 198 1 0 1599
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2911
timestamp 0
transform 0 -1 198 1 0 1598
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2910
timestamp 0
transform 0 -1 198 1 0 1597
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2909
timestamp 0
transform 0 -1 198 1 0 1596
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2908
timestamp 0
transform 0 -1 198 1 0 1595
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2907
timestamp 0
transform 0 -1 198 1 0 1594
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2906
timestamp 0
transform 0 -1 198 1 0 1593
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2905
timestamp 0
transform 0 -1 198 1 0 1592
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2904
timestamp 0
transform 0 -1 198 1 0 1591
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2903
timestamp 0
transform 0 -1 198 1 0 1590
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2902
timestamp 0
transform 0 -1 198 1 0 1589
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2901
timestamp 0
transform 0 -1 198 1 0 1588
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2900
timestamp 0
transform 0 -1 198 1 0 1587
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2899
timestamp 0
transform 0 -1 198 1 0 1586
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2898
timestamp 0
transform 0 -1 198 1 0 1585
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2897
timestamp 0
transform 0 -1 198 1 0 1584
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2896
timestamp 0
transform 0 -1 198 1 0 1583
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2895
timestamp 0
transform 0 -1 198 1 0 1582
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2894
timestamp 0
transform 0 -1 198 1 0 1581
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2893
timestamp 0
transform 0 -1 198 1 0 1580
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2892
timestamp 0
transform 0 -1 198 1 0 1579
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2891
timestamp 0
transform 0 -1 198 1 0 1578
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2890
timestamp 0
transform 0 -1 198 1 0 1577
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2889
timestamp 0
transform 0 -1 198 1 0 1576
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2888
timestamp 0
transform 0 -1 198 1 0 1575
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2887
timestamp 0
transform 0 -1 198 1 0 1574
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2886
timestamp 0
transform 0 -1 198 1 0 1573
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2885
timestamp 0
transform 0 -1 198 1 0 1572
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2884
timestamp 0
transform 0 -1 198 1 0 1571
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2883
timestamp 0
transform 0 -1 198 1 0 1570
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2882
timestamp 0
transform 0 -1 198 1 0 1569
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2881
timestamp 0
transform 0 -1 198 1 0 1568
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2880
timestamp 0
transform 0 -1 198 1 0 1567
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2879
timestamp 0
transform 0 -1 198 1 0 1566
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2878
timestamp 0
transform 0 -1 198 1 0 1565
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2877
timestamp 0
transform 0 -1 198 1 0 1564
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2876
timestamp 0
transform 0 -1 198 1 0 1563
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2875
timestamp 0
transform 0 -1 198 1 0 1562
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2874
timestamp 0
transform 0 -1 198 1 0 1561
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2873
timestamp 0
transform 0 -1 198 1 0 1560
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2872
timestamp 0
transform 0 -1 198 1 0 1559
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2871
timestamp 0
transform 0 -1 198 1 0 1558
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2870
timestamp 0
transform 0 -1 198 1 0 1557
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2869
timestamp 0
transform 0 -1 198 1 0 1556
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2868
timestamp 0
transform 0 -1 198 1 0 1555
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2867
timestamp 0
transform 0 -1 198 1 0 1554
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2866
timestamp 0
transform 0 -1 198 1 0 1553
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2865
timestamp 0
transform 0 -1 198 1 0 1552
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2864
timestamp 0
transform 0 -1 198 1 0 1551
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2863
timestamp 0
transform 0 -1 198 1 0 1550
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4143
timestamp 0
transform 0 1 2544 -1 0 1524
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4142
timestamp 0
transform 0 1 2544 -1 0 1523
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4141
timestamp 0
transform 0 1 2544 -1 0 1522
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4140
timestamp 0
transform 0 1 2544 -1 0 1521
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4139
timestamp 0
transform 0 1 2544 -1 0 1520
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4138
timestamp 0
transform 0 1 2544 -1 0 1519
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4137
timestamp 0
transform 0 1 2544 -1 0 1518
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4136
timestamp 0
transform 0 1 2544 -1 0 1517
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4135
timestamp 0
transform 0 1 2544 -1 0 1516
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4134
timestamp 0
transform 0 1 2544 -1 0 1515
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4133
timestamp 0
transform 0 1 2544 -1 0 1514
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4132
timestamp 0
transform 0 1 2544 -1 0 1513
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4131
timestamp 0
transform 0 1 2544 -1 0 1512
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4130
timestamp 0
transform 0 1 2544 -1 0 1511
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4129
timestamp 0
transform 0 1 2544 -1 0 1510
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4128
timestamp 0
transform 0 1 2544 -1 0 1509
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4127
timestamp 0
transform 0 1 2544 -1 0 1508
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4126
timestamp 0
transform 0 1 2544 -1 0 1507
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4125
timestamp 0
transform 0 1 2544 -1 0 1506
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4124
timestamp 0
transform 0 1 2544 -1 0 1505
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4123
timestamp 0
transform 0 1 2544 -1 0 1504
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4122
timestamp 0
transform 0 1 2544 -1 0 1503
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4121
timestamp 0
transform 0 1 2544 -1 0 1502
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4120
timestamp 0
transform 0 1 2544 -1 0 1501
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4119
timestamp 0
transform 0 1 2544 -1 0 1500
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4118
timestamp 0
transform 0 1 2544 -1 0 1499
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4117
timestamp 0
transform 0 1 2544 -1 0 1498
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4116
timestamp 0
transform 0 1 2544 -1 0 1497
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4115
timestamp 0
transform 0 1 2544 -1 0 1496
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4114
timestamp 0
transform 0 1 2544 -1 0 1495
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4113
timestamp 0
transform 0 1 2544 -1 0 1494
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4112
timestamp 0
transform 0 1 2544 -1 0 1493
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4111
timestamp 0
transform 0 1 2544 -1 0 1492
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4110
timestamp 0
transform 0 1 2544 -1 0 1491
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4109
timestamp 0
transform 0 1 2544 -1 0 1490
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4108
timestamp 0
transform 0 1 2544 -1 0 1489
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4107
timestamp 0
transform 0 1 2544 -1 0 1488
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4106
timestamp 0
transform 0 1 2544 -1 0 1487
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4105
timestamp 0
transform 0 1 2544 -1 0 1486
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4104
timestamp 0
transform 0 1 2544 -1 0 1485
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4103
timestamp 0
transform 0 1 2544 -1 0 1484
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4102
timestamp 0
transform 0 1 2544 -1 0 1483
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4101
timestamp 0
transform 0 1 2544 -1 0 1482
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4100
timestamp 0
transform 0 1 2544 -1 0 1481
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4099
timestamp 0
transform 0 1 2544 -1 0 1480
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4098
timestamp 0
transform 0 1 2544 -1 0 1479
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4097
timestamp 0
transform 0 1 2544 -1 0 1478
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4096
timestamp 0
transform 0 1 2544 -1 0 1477
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4095
timestamp 0
transform 0 1 2544 -1 0 1476
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4094
timestamp 0
transform 0 1 2544 -1 0 1475
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4093
timestamp 0
transform 0 1 2544 -1 0 1474
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4092
timestamp 0
transform 0 1 2544 -1 0 1473
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4091
timestamp 0
transform 0 1 2544 -1 0 1472
box 0 0 1 1
use s8iom0_gpiov2_pad  flash_clk_pad
timestamp 0
transform 0 -1 198 1 0 1470
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2861
timestamp 0
transform 0 -1 198 1 0 1469
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2860
timestamp 0
transform 0 -1 198 1 0 1468
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2859
timestamp 0
transform 0 -1 198 1 0 1467
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2858
timestamp 0
transform 0 -1 198 1 0 1466
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2857
timestamp 0
transform 0 -1 198 1 0 1465
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2856
timestamp 0
transform 0 -1 198 1 0 1464
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2855
timestamp 0
transform 0 -1 198 1 0 1463
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2854
timestamp 0
transform 0 -1 198 1 0 1462
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2853
timestamp 0
transform 0 -1 198 1 0 1461
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2852
timestamp 0
transform 0 -1 198 1 0 1460
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2851
timestamp 0
transform 0 -1 198 1 0 1459
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2850
timestamp 0
transform 0 -1 198 1 0 1458
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2849
timestamp 0
transform 0 -1 198 1 0 1457
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2848
timestamp 0
transform 0 -1 198 1 0 1456
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2847
timestamp 0
transform 0 -1 198 1 0 1455
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2846
timestamp 0
transform 0 -1 198 1 0 1454
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2845
timestamp 0
transform 0 -1 198 1 0 1453
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2844
timestamp 0
transform 0 -1 198 1 0 1452
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2843
timestamp 0
transform 0 -1 198 1 0 1451
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2842
timestamp 0
transform 0 -1 198 1 0 1450
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2841
timestamp 0
transform 0 -1 198 1 0 1449
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2840
timestamp 0
transform 0 -1 198 1 0 1448
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2839
timestamp 0
transform 0 -1 198 1 0 1447
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2838
timestamp 0
transform 0 -1 198 1 0 1446
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2837
timestamp 0
transform 0 -1 198 1 0 1445
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2836
timestamp 0
transform 0 -1 198 1 0 1444
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2835
timestamp 0
transform 0 -1 198 1 0 1443
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2834
timestamp 0
transform 0 -1 198 1 0 1442
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2833
timestamp 0
transform 0 -1 198 1 0 1441
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2832
timestamp 0
transform 0 -1 198 1 0 1440
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2831
timestamp 0
transform 0 -1 198 1 0 1439
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2830
timestamp 0
transform 0 -1 198 1 0 1438
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2829
timestamp 0
transform 0 -1 198 1 0 1437
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2828
timestamp 0
transform 0 -1 198 1 0 1436
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2827
timestamp 0
transform 0 -1 198 1 0 1435
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2826
timestamp 0
transform 0 -1 198 1 0 1434
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2825
timestamp 0
transform 0 -1 198 1 0 1433
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2824
timestamp 0
transform 0 -1 198 1 0 1432
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2823
timestamp 0
transform 0 -1 198 1 0 1431
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2822
timestamp 0
transform 0 -1 198 1 0 1430
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2821
timestamp 0
transform 0 -1 198 1 0 1429
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2820
timestamp 0
transform 0 -1 198 1 0 1428
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2819
timestamp 0
transform 0 -1 198 1 0 1427
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2818
timestamp 0
transform 0 -1 198 1 0 1426
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2817
timestamp 0
transform 0 -1 198 1 0 1425
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2816
timestamp 0
transform 0 -1 198 1 0 1424
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2815
timestamp 0
transform 0 -1 198 1 0 1423
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2814
timestamp 0
transform 0 -1 198 1 0 1422
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2813
timestamp 0
transform 0 -1 198 1 0 1421
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2812
timestamp 0
transform 0 -1 198 1 0 1420
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2811
timestamp 0
transform 0 -1 198 1 0 1419
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2810
timestamp 0
transform 0 -1 198 1 0 1418
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2809
timestamp 0
transform 0 -1 198 1 0 1417
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2808
timestamp 0
transform 0 -1 198 1 0 1416
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2807
timestamp 0
transform 0 -1 198 1 0 1415
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2806
timestamp 0
transform 0 -1 198 1 0 1414
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2805
timestamp 0
transform 0 -1 198 1 0 1413
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4090
timestamp 0
transform 0 1 2544 -1 0 1471
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4089
timestamp 0
transform 0 1 2544 -1 0 1470
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4088
timestamp 0
transform 0 1 2544 -1 0 1469
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4087
timestamp 0
transform 0 1 2544 -1 0 1468
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4086
timestamp 0
transform 0 1 2544 -1 0 1467
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4085
timestamp 0
transform 0 1 2544 -1 0 1466
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4084
timestamp 0
transform 0 1 2544 -1 0 1465
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4083
timestamp 0
transform 0 1 2544 -1 0 1464
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4082
timestamp 0
transform 0 1 2544 -1 0 1463
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4081
timestamp 0
transform 0 1 2544 -1 0 1462
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4080
timestamp 0
transform 0 1 2544 -1 0 1461
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4079
timestamp 0
transform 0 1 2544 -1 0 1460
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4078
timestamp 0
transform 0 1 2544 -1 0 1459
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4077
timestamp 0
transform 0 1 2544 -1 0 1458
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4076
timestamp 0
transform 0 1 2544 -1 0 1457
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4075
timestamp 0
transform 0 1 2544 -1 0 1456
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4074
timestamp 0
transform 0 1 2544 -1 0 1455
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4073
timestamp 0
transform 0 1 2544 -1 0 1454
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4072
timestamp 0
transform 0 1 2544 -1 0 1453
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4071
timestamp 0
transform 0 1 2544 -1 0 1452
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4070
timestamp 0
transform 0 1 2544 -1 0 1451
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4069
timestamp 0
transform 0 1 2544 -1 0 1450
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4068
timestamp 0
transform 0 1 2544 -1 0 1449
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4067
timestamp 0
transform 0 1 2544 -1 0 1448
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4066
timestamp 0
transform 0 1 2544 -1 0 1447
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4065
timestamp 0
transform 0 1 2544 -1 0 1446
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4064
timestamp 0
transform 0 1 2544 -1 0 1445
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4063
timestamp 0
transform 0 1 2544 -1 0 1444
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4062
timestamp 0
transform 0 1 2544 -1 0 1443
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4061
timestamp 0
transform 0 1 2544 -1 0 1442
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4060
timestamp 0
transform 0 1 2544 -1 0 1441
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4059
timestamp 0
transform 0 1 2544 -1 0 1440
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4058
timestamp 0
transform 0 1 2544 -1 0 1439
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4057
timestamp 0
transform 0 1 2544 -1 0 1438
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4056
timestamp 0
transform 0 1 2544 -1 0 1437
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4055
timestamp 0
transform 0 1 2544 -1 0 1436
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4054
timestamp 0
transform 0 1 2544 -1 0 1435
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4053
timestamp 0
transform 0 1 2544 -1 0 1434
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4052
timestamp 0
transform 0 1 2544 -1 0 1433
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4051
timestamp 0
transform 0 1 2544 -1 0 1432
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4050
timestamp 0
transform 0 1 2544 -1 0 1431
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4049
timestamp 0
transform 0 1 2544 -1 0 1430
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4048
timestamp 0
transform 0 1 2544 -1 0 1429
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4047
timestamp 0
transform 0 1 2544 -1 0 1428
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4046
timestamp 0
transform 0 1 2544 -1 0 1427
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4045
timestamp 0
transform 0 1 2544 -1 0 1426
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4044
timestamp 0
transform 0 1 2544 -1 0 1425
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4043
timestamp 0
transform 0 1 2544 -1 0 1424
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4042
timestamp 0
transform 0 1 2544 -1 0 1423
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4041
timestamp 0
transform 0 1 2544 -1 0 1422
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4040
timestamp 0
transform 0 1 2544 -1 0 1421
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4039
timestamp 0
transform 0 1 2544 -1 0 1420
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4038
timestamp 0
transform 0 1 2544 -1 0 1419
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4037
timestamp 0
transform 0 1 2544 -1 0 1418
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4036
timestamp 0
transform 0 1 2544 -1 0 1417
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4035
timestamp 0
transform 0 1 2544 -1 0 1416
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4034
timestamp 0
transform 0 1 2544 -1 0 1415
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4033
timestamp 0
transform 0 1 2544 -1 0 1414
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4032
timestamp 0
transform 0 1 2544 -1 0 1413
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4031
timestamp 0
transform 0 1 2544 -1 0 1412
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4030
timestamp 0
transform 0 1 2544 -1 0 1411
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4029
timestamp 0
transform 0 1 2544 -1 0 1410
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4028
timestamp 0
transform 0 1 2544 -1 0 1409
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4027
timestamp 0
transform 0 1 2544 -1 0 1408
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4026
timestamp 0
transform 0 1 2544 -1 0 1407
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4025
timestamp 0
transform 0 1 2544 -1 0 1406
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4024
timestamp 0
transform 0 1 2544 -1 0 1405
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4023
timestamp 0
transform 0 1 2544 -1 0 1404
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4022
timestamp 0
transform 0 1 2544 -1 0 1403
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4021
timestamp 0
transform 0 1 2544 -1 0 1402
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4020
timestamp 0
transform 0 1 2544 -1 0 1401
box 0 0 1 1
use s8iom0_gpiov2_pad  gpio_pad[4]
timestamp 0
transform 0 1 2544 -1 0 1400
box 0 0 1 1
use s8iom0_gpiov2_pad  xclk_pad
timestamp 0
transform 0 -1 198 1 0 1333
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2803
timestamp 0
transform 0 -1 198 1 0 1332
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2802
timestamp 0
transform 0 -1 198 1 0 1331
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2801
timestamp 0
transform 0 -1 198 1 0 1330
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2800
timestamp 0
transform 0 -1 198 1 0 1329
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2799
timestamp 0
transform 0 -1 198 1 0 1328
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2798
timestamp 0
transform 0 -1 198 1 0 1327
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2797
timestamp 0
transform 0 -1 198 1 0 1326
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2796
timestamp 0
transform 0 -1 198 1 0 1325
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2795
timestamp 0
transform 0 -1 198 1 0 1324
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2794
timestamp 0
transform 0 -1 198 1 0 1323
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2793
timestamp 0
transform 0 -1 198 1 0 1322
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2792
timestamp 0
transform 0 -1 198 1 0 1321
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2791
timestamp 0
transform 0 -1 198 1 0 1320
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2790
timestamp 0
transform 0 -1 198 1 0 1319
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2789
timestamp 0
transform 0 -1 198 1 0 1318
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2788
timestamp 0
transform 0 -1 198 1 0 1317
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2787
timestamp 0
transform 0 -1 198 1 0 1316
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2786
timestamp 0
transform 0 -1 198 1 0 1315
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2785
timestamp 0
transform 0 -1 198 1 0 1314
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2784
timestamp 0
transform 0 -1 198 1 0 1313
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2783
timestamp 0
transform 0 -1 198 1 0 1312
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2782
timestamp 0
transform 0 -1 198 1 0 1311
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2781
timestamp 0
transform 0 -1 198 1 0 1310
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2780
timestamp 0
transform 0 -1 198 1 0 1309
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2779
timestamp 0
transform 0 -1 198 1 0 1308
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2778
timestamp 0
transform 0 -1 198 1 0 1307
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2777
timestamp 0
transform 0 -1 198 1 0 1306
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2776
timestamp 0
transform 0 -1 198 1 0 1305
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2775
timestamp 0
transform 0 -1 198 1 0 1304
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2774
timestamp 0
transform 0 -1 198 1 0 1303
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2773
timestamp 0
transform 0 -1 198 1 0 1302
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2772
timestamp 0
transform 0 -1 198 1 0 1301
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2771
timestamp 0
transform 0 -1 198 1 0 1300
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2770
timestamp 0
transform 0 -1 198 1 0 1299
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2769
timestamp 0
transform 0 -1 198 1 0 1298
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2768
timestamp 0
transform 0 -1 198 1 0 1297
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2767
timestamp 0
transform 0 -1 198 1 0 1296
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2766
timestamp 0
transform 0 -1 198 1 0 1295
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2765
timestamp 0
transform 0 -1 198 1 0 1294
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2764
timestamp 0
transform 0 -1 198 1 0 1293
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2763
timestamp 0
transform 0 -1 198 1 0 1292
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2762
timestamp 0
transform 0 -1 198 1 0 1291
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2761
timestamp 0
transform 0 -1 198 1 0 1290
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2760
timestamp 0
transform 0 -1 198 1 0 1289
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2759
timestamp 0
transform 0 -1 198 1 0 1288
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2758
timestamp 0
transform 0 -1 198 1 0 1287
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2757
timestamp 0
transform 0 -1 198 1 0 1286
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2756
timestamp 0
transform 0 -1 198 1 0 1285
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2755
timestamp 0
transform 0 -1 198 1 0 1284
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2754
timestamp 0
transform 0 -1 198 1 0 1283
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2753
timestamp 0
transform 0 -1 198 1 0 1282
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2752
timestamp 0
transform 0 -1 198 1 0 1281
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2751
timestamp 0
transform 0 -1 198 1 0 1280
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2750
timestamp 0
transform 0 -1 198 1 0 1279
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2749
timestamp 0
transform 0 -1 198 1 0 1278
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2748
timestamp 0
transform 0 -1 198 1 0 1277
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2747
timestamp 0
transform 0 -1 198 1 0 1276
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2746
timestamp 0
transform 0 -1 198 1 0 1275
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4018
timestamp 0
transform 0 1 2544 -1 0 1320
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4017
timestamp 0
transform 0 1 2544 -1 0 1319
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4016
timestamp 0
transform 0 1 2544 -1 0 1318
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4015
timestamp 0
transform 0 1 2544 -1 0 1317
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4014
timestamp 0
transform 0 1 2544 -1 0 1316
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4013
timestamp 0
transform 0 1 2544 -1 0 1315
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4012
timestamp 0
transform 0 1 2544 -1 0 1314
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4011
timestamp 0
transform 0 1 2544 -1 0 1313
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4010
timestamp 0
transform 0 1 2544 -1 0 1312
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4009
timestamp 0
transform 0 1 2544 -1 0 1311
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4008
timestamp 0
transform 0 1 2544 -1 0 1310
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4007
timestamp 0
transform 0 1 2544 -1 0 1309
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4006
timestamp 0
transform 0 1 2544 -1 0 1308
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4005
timestamp 0
transform 0 1 2544 -1 0 1307
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4004
timestamp 0
transform 0 1 2544 -1 0 1306
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4003
timestamp 0
transform 0 1 2544 -1 0 1305
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4002
timestamp 0
transform 0 1 2544 -1 0 1304
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4001
timestamp 0
transform 0 1 2544 -1 0 1303
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_4000
timestamp 0
transform 0 1 2544 -1 0 1302
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3999
timestamp 0
transform 0 1 2544 -1 0 1301
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3998
timestamp 0
transform 0 1 2544 -1 0 1300
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3997
timestamp 0
transform 0 1 2544 -1 0 1299
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3996
timestamp 0
transform 0 1 2544 -1 0 1298
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3995
timestamp 0
transform 0 1 2544 -1 0 1297
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3994
timestamp 0
transform 0 1 2544 -1 0 1296
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3993
timestamp 0
transform 0 1 2544 -1 0 1295
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3992
timestamp 0
transform 0 1 2544 -1 0 1294
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3991
timestamp 0
transform 0 1 2544 -1 0 1293
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3990
timestamp 0
transform 0 1 2544 -1 0 1292
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3989
timestamp 0
transform 0 1 2544 -1 0 1291
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3988
timestamp 0
transform 0 1 2544 -1 0 1290
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3987
timestamp 0
transform 0 1 2544 -1 0 1289
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3986
timestamp 0
transform 0 1 2544 -1 0 1288
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3985
timestamp 0
transform 0 1 2544 -1 0 1287
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3984
timestamp 0
transform 0 1 2544 -1 0 1286
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3983
timestamp 0
transform 0 1 2544 -1 0 1285
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3982
timestamp 0
transform 0 1 2544 -1 0 1284
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3981
timestamp 0
transform 0 1 2544 -1 0 1283
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3980
timestamp 0
transform 0 1 2544 -1 0 1282
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3979
timestamp 0
transform 0 1 2544 -1 0 1281
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3978
timestamp 0
transform 0 1 2544 -1 0 1280
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3977
timestamp 0
transform 0 1 2544 -1 0 1279
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3976
timestamp 0
transform 0 1 2544 -1 0 1278
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3975
timestamp 0
transform 0 1 2544 -1 0 1277
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3974
timestamp 0
transform 0 1 2544 -1 0 1276
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3973
timestamp 0
transform 0 1 2544 -1 0 1275
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3972
timestamp 0
transform 0 1 2544 -1 0 1274
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3971
timestamp 0
transform 0 1 2544 -1 0 1273
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3970
timestamp 0
transform 0 1 2544 -1 0 1272
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3969
timestamp 0
transform 0 1 2544 -1 0 1271
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3968
timestamp 0
transform 0 1 2544 -1 0 1270
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3967
timestamp 0
transform 0 1 2544 -1 0 1269
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3966
timestamp 0
transform 0 1 2544 -1 0 1268
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3965
timestamp 0
transform 0 1 2544 -1 0 1267
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3964
timestamp 0
transform 0 1 2544 -1 0 1266
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3963
timestamp 0
transform 0 1 2544 -1 0 1265
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3962
timestamp 0
transform 0 1 2544 -1 0 1264
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3961
timestamp 0
transform 0 1 2544 -1 0 1263
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3960
timestamp 0
transform 0 1 2544 -1 0 1262
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3959
timestamp 0
transform 0 1 2544 -1 0 1261
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3958
timestamp 0
transform 0 1 2544 -1 0 1260
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3957
timestamp 0
transform 0 1 2544 -1 0 1259
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3956
timestamp 0
transform 0 1 2544 -1 0 1258
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3955
timestamp 0
transform 0 1 2544 -1 0 1257
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3954
timestamp 0
transform 0 1 2544 -1 0 1256
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3953
timestamp 0
transform 0 1 2544 -1 0 1255
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3952
timestamp 0
transform 0 1 2544 -1 0 1254
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3951
timestamp 0
transform 0 1 2544 -1 0 1253
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3950
timestamp 0
transform 0 1 2544 -1 0 1252
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3949
timestamp 0
transform 0 1 2544 -1 0 1251
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3948
timestamp 0
transform 0 1 2544 -1 0 1250
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3947
timestamp 0
transform 0 1 2544 -1 0 1249
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3946
timestamp 0
transform 0 1 2544 -1 0 1248
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3945
timestamp 0
transform 0 1 2544 -1 0 1247
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3944
timestamp 0
transform 0 1 2544 -1 0 1246
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3943
timestamp 0
transform 0 1 2544 -1 0 1245
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3942
timestamp 0
transform 0 1 2544 -1 0 1244
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3941
timestamp 0
transform 0 1 2544 -1 0 1243
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3940
timestamp 0
transform 0 1 2544 -1 0 1242
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3939
timestamp 0
transform 0 1 2544 -1 0 1241
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3938
timestamp 0
transform 0 1 2544 -1 0 1240
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3937
timestamp 0
transform 0 1 2544 -1 0 1239
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3936
timestamp 0
transform 0 1 2544 -1 0 1238
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3935
timestamp 0
transform 0 1 2544 -1 0 1237
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3934
timestamp 0
transform 0 1 2544 -1 0 1236
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3933
timestamp 0
transform 0 1 2544 -1 0 1235
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3932
timestamp 0
transform 0 1 2544 -1 0 1234
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3931
timestamp 0
transform 0 1 2544 -1 0 1233
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3930
timestamp 0
transform 0 1 2544 -1 0 1232
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3929
timestamp 0
transform 0 1 2544 -1 0 1231
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3928
timestamp 0
transform 0 1 2544 -1 0 1230
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3927
timestamp 0
transform 0 1 2544 -1 0 1229
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3926
timestamp 0
transform 0 1 2544 -1 0 1228
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3925
timestamp 0
transform 0 1 2544 -1 0 1227
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3924
timestamp 0
transform 0 1 2544 -1 0 1226
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3923
timestamp 0
transform 0 1 2544 -1 0 1225
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3922
timestamp 0
transform 0 1 2544 -1 0 1224
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3921
timestamp 0
transform 0 1 2544 -1 0 1223
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3920
timestamp 0
transform 0 1 2544 -1 0 1222
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3919
timestamp 0
transform 0 1 2544 -1 0 1221
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3918
timestamp 0
transform 0 1 2544 -1 0 1220
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3917
timestamp 0
transform 0 1 2544 -1 0 1219
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3916
timestamp 0
transform 0 1 2544 -1 0 1218
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3915
timestamp 0
transform 0 1 2544 -1 0 1217
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3914
timestamp 0
transform 0 1 2544 -1 0 1216
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3913
timestamp 0
transform 0 1 2544 -1 0 1215
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3912
timestamp 0
transform 0 1 2544 -1 0 1214
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3911
timestamp 0
transform 0 1 2544 -1 0 1213
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3910
timestamp 0
transform 0 1 2544 -1 0 1212
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3909
timestamp 0
transform 0 1 2544 -1 0 1211
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3908
timestamp 0
transform 0 1 2544 -1 0 1210
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3907
timestamp 0
transform 0 1 2544 -1 0 1209
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3906
timestamp 0
transform 0 1 2544 -1 0 1208
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3905
timestamp 0
transform 0 1 2544 -1 0 1207
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3904
timestamp 0
transform 0 1 2544 -1 0 1206
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3903
timestamp 0
transform 0 1 2544 -1 0 1205
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3902
timestamp 0
transform 0 1 2544 -1 0 1204
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3901
timestamp 0
transform 0 1 2544 -1 0 1203
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3900
timestamp 0
transform 0 1 2544 -1 0 1202
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3899
timestamp 0
transform 0 1 2544 -1 0 1201
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3898
timestamp 0
transform 0 1 2544 -1 0 1200
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3897
timestamp 0
transform 0 1 2544 -1 0 1199
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3896
timestamp 0
transform 0 1 2544 -1 0 1198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3895
timestamp 0
transform 0 1 2544 -1 0 1197
box 0 0 1 1
use s8iom0_gpiov2_pad  SCK_pad
timestamp 0
transform 0 -1 198 1 0 1195
box 0 0 1 1
use s8iom0_vssd_lvc_pad  vssdlclamp
timestamp 0
transform 0 1 2544 -1 0 1196
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2744
timestamp 0
transform 0 -1 198 1 0 1194
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2743
timestamp 0
transform 0 -1 198 1 0 1193
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2742
timestamp 0
transform 0 -1 198 1 0 1192
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2741
timestamp 0
transform 0 -1 198 1 0 1191
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2740
timestamp 0
transform 0 -1 198 1 0 1190
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2739
timestamp 0
transform 0 -1 198 1 0 1189
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2738
timestamp 0
transform 0 -1 198 1 0 1188
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2737
timestamp 0
transform 0 -1 198 1 0 1187
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2736
timestamp 0
transform 0 -1 198 1 0 1186
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2735
timestamp 0
transform 0 -1 198 1 0 1185
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2734
timestamp 0
transform 0 -1 198 1 0 1184
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2733
timestamp 0
transform 0 -1 198 1 0 1183
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2732
timestamp 0
transform 0 -1 198 1 0 1182
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2731
timestamp 0
transform 0 -1 198 1 0 1181
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2730
timestamp 0
transform 0 -1 198 1 0 1180
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2729
timestamp 0
transform 0 -1 198 1 0 1179
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2728
timestamp 0
transform 0 -1 198 1 0 1178
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2727
timestamp 0
transform 0 -1 198 1 0 1177
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2726
timestamp 0
transform 0 -1 198 1 0 1176
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2725
timestamp 0
transform 0 -1 198 1 0 1175
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2724
timestamp 0
transform 0 -1 198 1 0 1174
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2723
timestamp 0
transform 0 -1 198 1 0 1173
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2722
timestamp 0
transform 0 -1 198 1 0 1172
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2721
timestamp 0
transform 0 -1 198 1 0 1171
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2720
timestamp 0
transform 0 -1 198 1 0 1170
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2719
timestamp 0
transform 0 -1 198 1 0 1169
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2718
timestamp 0
transform 0 -1 198 1 0 1168
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2717
timestamp 0
transform 0 -1 198 1 0 1167
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2716
timestamp 0
transform 0 -1 198 1 0 1166
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2715
timestamp 0
transform 0 -1 198 1 0 1165
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2714
timestamp 0
transform 0 -1 198 1 0 1164
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2713
timestamp 0
transform 0 -1 198 1 0 1163
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2712
timestamp 0
transform 0 -1 198 1 0 1162
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2711
timestamp 0
transform 0 -1 198 1 0 1161
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2710
timestamp 0
transform 0 -1 198 1 0 1160
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2709
timestamp 0
transform 0 -1 198 1 0 1159
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2708
timestamp 0
transform 0 -1 198 1 0 1158
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2707
timestamp 0
transform 0 -1 198 1 0 1157
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2706
timestamp 0
transform 0 -1 198 1 0 1156
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2705
timestamp 0
transform 0 -1 198 1 0 1155
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2704
timestamp 0
transform 0 -1 198 1 0 1154
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2703
timestamp 0
transform 0 -1 198 1 0 1153
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2702
timestamp 0
transform 0 -1 198 1 0 1152
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2701
timestamp 0
transform 0 -1 198 1 0 1151
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2700
timestamp 0
transform 0 -1 198 1 0 1150
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2699
timestamp 0
transform 0 -1 198 1 0 1149
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2698
timestamp 0
transform 0 -1 198 1 0 1148
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2697
timestamp 0
transform 0 -1 198 1 0 1147
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2696
timestamp 0
transform 0 -1 198 1 0 1146
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2695
timestamp 0
transform 0 -1 198 1 0 1145
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2694
timestamp 0
transform 0 -1 198 1 0 1144
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2693
timestamp 0
transform 0 -1 198 1 0 1143
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2692
timestamp 0
transform 0 -1 198 1 0 1142
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2691
timestamp 0
transform 0 -1 198 1 0 1141
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2690
timestamp 0
transform 0 -1 198 1 0 1140
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2689
timestamp 0
transform 0 -1 198 1 0 1139
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2688
timestamp 0
transform 0 -1 198 1 0 1138
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3893
timestamp 0
transform 0 1 2544 -1 0 1121
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3892
timestamp 0
transform 0 1 2544 -1 0 1120
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3891
timestamp 0
transform 0 1 2544 -1 0 1119
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3890
timestamp 0
transform 0 1 2544 -1 0 1118
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3889
timestamp 0
transform 0 1 2544 -1 0 1117
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3888
timestamp 0
transform 0 1 2544 -1 0 1116
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3887
timestamp 0
transform 0 1 2544 -1 0 1115
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3886
timestamp 0
transform 0 1 2544 -1 0 1114
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3885
timestamp 0
transform 0 1 2544 -1 0 1113
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3884
timestamp 0
transform 0 1 2544 -1 0 1112
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3883
timestamp 0
transform 0 1 2544 -1 0 1111
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3882
timestamp 0
transform 0 1 2544 -1 0 1110
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3881
timestamp 0
transform 0 1 2544 -1 0 1109
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3880
timestamp 0
transform 0 1 2544 -1 0 1108
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3879
timestamp 0
transform 0 1 2544 -1 0 1107
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3878
timestamp 0
transform 0 1 2544 -1 0 1106
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3877
timestamp 0
transform 0 1 2544 -1 0 1105
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3876
timestamp 0
transform 0 1 2544 -1 0 1104
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3875
timestamp 0
transform 0 1 2544 -1 0 1103
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3874
timestamp 0
transform 0 1 2544 -1 0 1102
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3873
timestamp 0
transform 0 1 2544 -1 0 1101
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3872
timestamp 0
transform 0 1 2544 -1 0 1100
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3871
timestamp 0
transform 0 1 2544 -1 0 1099
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3870
timestamp 0
transform 0 1 2544 -1 0 1098
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3869
timestamp 0
transform 0 1 2544 -1 0 1097
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3868
timestamp 0
transform 0 1 2544 -1 0 1096
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3867
timestamp 0
transform 0 1 2544 -1 0 1095
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3866
timestamp 0
transform 0 1 2544 -1 0 1094
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3865
timestamp 0
transform 0 1 2544 -1 0 1093
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3864
timestamp 0
transform 0 1 2544 -1 0 1092
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3863
timestamp 0
transform 0 1 2544 -1 0 1091
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3862
timestamp 0
transform 0 1 2544 -1 0 1090
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3861
timestamp 0
transform 0 1 2544 -1 0 1089
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3860
timestamp 0
transform 0 1 2544 -1 0 1088
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3859
timestamp 0
transform 0 1 2544 -1 0 1087
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3858
timestamp 0
transform 0 1 2544 -1 0 1086
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3857
timestamp 0
transform 0 1 2544 -1 0 1085
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3856
timestamp 0
transform 0 1 2544 -1 0 1084
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3855
timestamp 0
transform 0 1 2544 -1 0 1083
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3854
timestamp 0
transform 0 1 2544 -1 0 1082
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3853
timestamp 0
transform 0 1 2544 -1 0 1081
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3852
timestamp 0
transform 0 1 2544 -1 0 1080
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3851
timestamp 0
transform 0 1 2544 -1 0 1079
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3850
timestamp 0
transform 0 1 2544 -1 0 1078
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3849
timestamp 0
transform 0 1 2544 -1 0 1077
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3848
timestamp 0
transform 0 1 2544 -1 0 1076
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3847
timestamp 0
transform 0 1 2544 -1 0 1075
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3846
timestamp 0
transform 0 1 2544 -1 0 1074
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3845
timestamp 0
transform 0 1 2544 -1 0 1073
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3844
timestamp 0
transform 0 1 2544 -1 0 1072
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3843
timestamp 0
transform 0 1 2544 -1 0 1071
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3842
timestamp 0
transform 0 1 2544 -1 0 1070
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3841
timestamp 0
transform 0 1 2544 -1 0 1069
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3840
timestamp 0
transform 0 1 2544 -1 0 1068
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3839
timestamp 0
transform 0 1 2544 -1 0 1067
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3838
timestamp 0
transform 0 1 2544 -1 0 1066
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3837
timestamp 0
transform 0 1 2544 -1 0 1065
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3836
timestamp 0
transform 0 1 2544 -1 0 1064
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3835
timestamp 0
transform 0 1 2544 -1 0 1063
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3834
timestamp 0
transform 0 1 2544 -1 0 1062
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3833
timestamp 0
transform 0 1 2544 -1 0 1061
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3832
timestamp 0
transform 0 1 2544 -1 0 1060
box 0 0 1 1
use s8iom0_gpiov2_pad  CSB_pad
timestamp 0
transform 0 -1 198 1 0 1058
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2686
timestamp 0
transform 0 -1 198 1 0 1057
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2685
timestamp 0
transform 0 -1 198 1 0 1056
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2684
timestamp 0
transform 0 -1 198 1 0 1055
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2683
timestamp 0
transform 0 -1 198 1 0 1054
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2682
timestamp 0
transform 0 -1 198 1 0 1053
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2681
timestamp 0
transform 0 -1 198 1 0 1052
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2680
timestamp 0
transform 0 -1 198 1 0 1051
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2679
timestamp 0
transform 0 -1 198 1 0 1050
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2678
timestamp 0
transform 0 -1 198 1 0 1049
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2677
timestamp 0
transform 0 -1 198 1 0 1048
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2676
timestamp 0
transform 0 -1 198 1 0 1047
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2675
timestamp 0
transform 0 -1 198 1 0 1046
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2674
timestamp 0
transform 0 -1 198 1 0 1045
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2673
timestamp 0
transform 0 -1 198 1 0 1044
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2672
timestamp 0
transform 0 -1 198 1 0 1043
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2671
timestamp 0
transform 0 -1 198 1 0 1042
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2670
timestamp 0
transform 0 -1 198 1 0 1041
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2669
timestamp 0
transform 0 -1 198 1 0 1040
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2668
timestamp 0
transform 0 -1 198 1 0 1039
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2667
timestamp 0
transform 0 -1 198 1 0 1038
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2666
timestamp 0
transform 0 -1 198 1 0 1037
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2665
timestamp 0
transform 0 -1 198 1 0 1036
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2664
timestamp 0
transform 0 -1 198 1 0 1035
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2663
timestamp 0
transform 0 -1 198 1 0 1034
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2662
timestamp 0
transform 0 -1 198 1 0 1033
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2661
timestamp 0
transform 0 -1 198 1 0 1032
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2660
timestamp 0
transform 0 -1 198 1 0 1031
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2659
timestamp 0
transform 0 -1 198 1 0 1030
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2658
timestamp 0
transform 0 -1 198 1 0 1029
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2657
timestamp 0
transform 0 -1 198 1 0 1028
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2656
timestamp 0
transform 0 -1 198 1 0 1027
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2655
timestamp 0
transform 0 -1 198 1 0 1026
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2654
timestamp 0
transform 0 -1 198 1 0 1025
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2653
timestamp 0
transform 0 -1 198 1 0 1024
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2652
timestamp 0
transform 0 -1 198 1 0 1023
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2651
timestamp 0
transform 0 -1 198 1 0 1022
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2650
timestamp 0
transform 0 -1 198 1 0 1021
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2649
timestamp 0
transform 0 -1 198 1 0 1020
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2648
timestamp 0
transform 0 -1 198 1 0 1019
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2647
timestamp 0
transform 0 -1 198 1 0 1018
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2646
timestamp 0
transform 0 -1 198 1 0 1017
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2645
timestamp 0
transform 0 -1 198 1 0 1016
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2644
timestamp 0
transform 0 -1 198 1 0 1015
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2643
timestamp 0
transform 0 -1 198 1 0 1014
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2642
timestamp 0
transform 0 -1 198 1 0 1013
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2641
timestamp 0
transform 0 -1 198 1 0 1012
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2640
timestamp 0
transform 0 -1 198 1 0 1011
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2639
timestamp 0
transform 0 -1 198 1 0 1010
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2638
timestamp 0
transform 0 -1 198 1 0 1009
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2637
timestamp 0
transform 0 -1 198 1 0 1008
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2636
timestamp 0
transform 0 -1 198 1 0 1007
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2635
timestamp 0
transform 0 -1 198 1 0 1006
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2634
timestamp 0
transform 0 -1 198 1 0 1005
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2633
timestamp 0
transform 0 -1 198 1 0 1004
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2632
timestamp 0
transform 0 -1 198 1 0 1003
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2631
timestamp 0
transform 0 -1 198 1 0 1002
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2630
timestamp 0
transform 0 -1 198 1 0 1001
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3831
timestamp 0
transform 0 1 2544 -1 0 1059
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3830
timestamp 0
transform 0 1 2544 -1 0 1058
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3829
timestamp 0
transform 0 1 2544 -1 0 1057
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3828
timestamp 0
transform 0 1 2544 -1 0 1056
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3827
timestamp 0
transform 0 1 2544 -1 0 1055
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3826
timestamp 0
transform 0 1 2544 -1 0 1054
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3825
timestamp 0
transform 0 1 2544 -1 0 1053
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3824
timestamp 0
transform 0 1 2544 -1 0 1052
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3823
timestamp 0
transform 0 1 2544 -1 0 1051
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3822
timestamp 0
transform 0 1 2544 -1 0 1050
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3821
timestamp 0
transform 0 1 2544 -1 0 1049
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3820
timestamp 0
transform 0 1 2544 -1 0 1048
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3819
timestamp 0
transform 0 1 2544 -1 0 1047
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3818
timestamp 0
transform 0 1 2544 -1 0 1046
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3817
timestamp 0
transform 0 1 2544 -1 0 1045
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3816
timestamp 0
transform 0 1 2544 -1 0 1044
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3815
timestamp 0
transform 0 1 2544 -1 0 1043
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3814
timestamp 0
transform 0 1 2544 -1 0 1042
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3813
timestamp 0
transform 0 1 2544 -1 0 1041
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3812
timestamp 0
transform 0 1 2544 -1 0 1040
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3811
timestamp 0
transform 0 1 2544 -1 0 1039
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3810
timestamp 0
transform 0 1 2544 -1 0 1038
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3809
timestamp 0
transform 0 1 2544 -1 0 1037
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3808
timestamp 0
transform 0 1 2544 -1 0 1036
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3807
timestamp 0
transform 0 1 2544 -1 0 1035
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3806
timestamp 0
transform 0 1 2544 -1 0 1034
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3805
timestamp 0
transform 0 1 2544 -1 0 1033
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3804
timestamp 0
transform 0 1 2544 -1 0 1032
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3803
timestamp 0
transform 0 1 2544 -1 0 1031
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3802
timestamp 0
transform 0 1 2544 -1 0 1030
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3801
timestamp 0
transform 0 1 2544 -1 0 1029
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3800
timestamp 0
transform 0 1 2544 -1 0 1028
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3799
timestamp 0
transform 0 1 2544 -1 0 1027
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3798
timestamp 0
transform 0 1 2544 -1 0 1026
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3797
timestamp 0
transform 0 1 2544 -1 0 1025
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3796
timestamp 0
transform 0 1 2544 -1 0 1024
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3795
timestamp 0
transform 0 1 2544 -1 0 1023
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3794
timestamp 0
transform 0 1 2544 -1 0 1022
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3793
timestamp 0
transform 0 1 2544 -1 0 1021
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3792
timestamp 0
transform 0 1 2544 -1 0 1020
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3791
timestamp 0
transform 0 1 2544 -1 0 1019
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3790
timestamp 0
transform 0 1 2544 -1 0 1018
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3789
timestamp 0
transform 0 1 2544 -1 0 1017
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3788
timestamp 0
transform 0 1 2544 -1 0 1016
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3787
timestamp 0
transform 0 1 2544 -1 0 1015
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3786
timestamp 0
transform 0 1 2544 -1 0 1014
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3785
timestamp 0
transform 0 1 2544 -1 0 1013
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3784
timestamp 0
transform 0 1 2544 -1 0 1012
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3783
timestamp 0
transform 0 1 2544 -1 0 1011
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3782
timestamp 0
transform 0 1 2544 -1 0 1010
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3781
timestamp 0
transform 0 1 2544 -1 0 1009
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3780
timestamp 0
transform 0 1 2544 -1 0 1008
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3779
timestamp 0
transform 0 1 2544 -1 0 1007
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3778
timestamp 0
transform 0 1 2544 -1 0 1006
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3777
timestamp 0
transform 0 1 2544 -1 0 1005
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3776
timestamp 0
transform 0 1 2544 -1 0 1004
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3775
timestamp 0
transform 0 1 2544 -1 0 1003
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3774
timestamp 0
transform 0 1 2544 -1 0 1002
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3773
timestamp 0
transform 0 1 2544 -1 0 1001
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3772
timestamp 0
transform 0 1 2544 -1 0 1000
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3771
timestamp 0
transform 0 1 2544 -1 0 999
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3770
timestamp 0
transform 0 1 2544 -1 0 998
box 0 0 1 1
use s8iom0_vssa_hvc_pad  vsshclamp[3]
timestamp 0
transform 0 1 2544 -1 0 997
box 0 0 1 1
use s8iom0s8_top_xres4v2  RSTB_pad
timestamp 0
transform 0 -1 200 1 0 926
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2628
timestamp 0
transform 0 -1 198 1 0 925
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2627
timestamp 0
transform 0 -1 198 1 0 924
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2626
timestamp 0
transform 0 -1 198 1 0 923
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2625
timestamp 0
transform 0 -1 198 1 0 922
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2624
timestamp 0
transform 0 -1 198 1 0 921
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2623
timestamp 0
transform 0 -1 198 1 0 920
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2622
timestamp 0
transform 0 -1 198 1 0 919
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2621
timestamp 0
transform 0 -1 198 1 0 918
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2620
timestamp 0
transform 0 -1 198 1 0 917
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2619
timestamp 0
transform 0 -1 198 1 0 916
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2618
timestamp 0
transform 0 -1 198 1 0 915
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2617
timestamp 0
transform 0 -1 198 1 0 914
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2616
timestamp 0
transform 0 -1 198 1 0 913
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2615
timestamp 0
transform 0 -1 198 1 0 912
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2614
timestamp 0
transform 0 -1 198 1 0 911
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2613
timestamp 0
transform 0 -1 198 1 0 910
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2612
timestamp 0
transform 0 -1 198 1 0 909
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2611
timestamp 0
transform 0 -1 198 1 0 908
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2610
timestamp 0
transform 0 -1 198 1 0 907
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2609
timestamp 0
transform 0 -1 198 1 0 906
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2608
timestamp 0
transform 0 -1 198 1 0 905
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2607
timestamp 0
transform 0 -1 198 1 0 904
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2606
timestamp 0
transform 0 -1 198 1 0 903
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2605
timestamp 0
transform 0 -1 198 1 0 902
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2604
timestamp 0
transform 0 -1 198 1 0 901
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2603
timestamp 0
transform 0 -1 198 1 0 900
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2602
timestamp 0
transform 0 -1 198 1 0 899
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2601
timestamp 0
transform 0 -1 198 1 0 898
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2600
timestamp 0
transform 0 -1 198 1 0 897
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2599
timestamp 0
transform 0 -1 198 1 0 896
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2598
timestamp 0
transform 0 -1 198 1 0 895
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2597
timestamp 0
transform 0 -1 198 1 0 894
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2596
timestamp 0
transform 0 -1 198 1 0 893
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2595
timestamp 0
transform 0 -1 198 1 0 892
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2594
timestamp 0
transform 0 -1 198 1 0 891
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2593
timestamp 0
transform 0 -1 198 1 0 890
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2592
timestamp 0
transform 0 -1 198 1 0 889
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2591
timestamp 0
transform 0 -1 198 1 0 888
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2590
timestamp 0
transform 0 -1 198 1 0 887
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2589
timestamp 0
transform 0 -1 198 1 0 886
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2588
timestamp 0
transform 0 -1 198 1 0 885
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2587
timestamp 0
transform 0 -1 198 1 0 884
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2586
timestamp 0
transform 0 -1 198 1 0 883
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2585
timestamp 0
transform 0 -1 198 1 0 882
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2584
timestamp 0
transform 0 -1 198 1 0 881
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2583
timestamp 0
transform 0 -1 198 1 0 880
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2582
timestamp 0
transform 0 -1 198 1 0 879
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2581
timestamp 0
transform 0 -1 198 1 0 878
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2580
timestamp 0
transform 0 -1 198 1 0 877
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2579
timestamp 0
transform 0 -1 198 1 0 876
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2578
timestamp 0
transform 0 -1 198 1 0 875
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2577
timestamp 0
transform 0 -1 198 1 0 874
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2576
timestamp 0
transform 0 -1 198 1 0 873
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2575
timestamp 0
transform 0 -1 198 1 0 872
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2574
timestamp 0
transform 0 -1 198 1 0 871
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2573
timestamp 0
transform 0 -1 198 1 0 870
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2572
timestamp 0
transform 0 -1 198 1 0 869
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3768
timestamp 0
transform 0 1 2544 -1 0 922
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3767
timestamp 0
transform 0 1 2544 -1 0 921
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3766
timestamp 0
transform 0 1 2544 -1 0 920
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3765
timestamp 0
transform 0 1 2544 -1 0 919
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3764
timestamp 0
transform 0 1 2544 -1 0 918
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3763
timestamp 0
transform 0 1 2544 -1 0 917
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3762
timestamp 0
transform 0 1 2544 -1 0 916
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3761
timestamp 0
transform 0 1 2544 -1 0 915
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3760
timestamp 0
transform 0 1 2544 -1 0 914
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3759
timestamp 0
transform 0 1 2544 -1 0 913
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3758
timestamp 0
transform 0 1 2544 -1 0 912
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3757
timestamp 0
transform 0 1 2544 -1 0 911
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3756
timestamp 0
transform 0 1 2544 -1 0 910
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3755
timestamp 0
transform 0 1 2544 -1 0 909
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3754
timestamp 0
transform 0 1 2544 -1 0 908
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3753
timestamp 0
transform 0 1 2544 -1 0 907
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3752
timestamp 0
transform 0 1 2544 -1 0 906
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3751
timestamp 0
transform 0 1 2544 -1 0 905
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3750
timestamp 0
transform 0 1 2544 -1 0 904
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3749
timestamp 0
transform 0 1 2544 -1 0 903
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3748
timestamp 0
transform 0 1 2544 -1 0 902
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3747
timestamp 0
transform 0 1 2544 -1 0 901
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3746
timestamp 0
transform 0 1 2544 -1 0 900
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3745
timestamp 0
transform 0 1 2544 -1 0 899
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3744
timestamp 0
transform 0 1 2544 -1 0 898
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3743
timestamp 0
transform 0 1 2544 -1 0 897
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3742
timestamp 0
transform 0 1 2544 -1 0 896
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3741
timestamp 0
transform 0 1 2544 -1 0 895
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3740
timestamp 0
transform 0 1 2544 -1 0 894
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3739
timestamp 0
transform 0 1 2544 -1 0 893
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3738
timestamp 0
transform 0 1 2544 -1 0 892
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3737
timestamp 0
transform 0 1 2544 -1 0 891
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3736
timestamp 0
transform 0 1 2544 -1 0 890
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3735
timestamp 0
transform 0 1 2544 -1 0 889
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3734
timestamp 0
transform 0 1 2544 -1 0 888
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3733
timestamp 0
transform 0 1 2544 -1 0 887
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3732
timestamp 0
transform 0 1 2544 -1 0 886
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3731
timestamp 0
transform 0 1 2544 -1 0 885
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3730
timestamp 0
transform 0 1 2544 -1 0 884
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3729
timestamp 0
transform 0 1 2544 -1 0 883
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3728
timestamp 0
transform 0 1 2544 -1 0 882
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3727
timestamp 0
transform 0 1 2544 -1 0 881
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3726
timestamp 0
transform 0 1 2544 -1 0 880
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3725
timestamp 0
transform 0 1 2544 -1 0 879
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3724
timestamp 0
transform 0 1 2544 -1 0 878
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3723
timestamp 0
transform 0 1 2544 -1 0 877
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3722
timestamp 0
transform 0 1 2544 -1 0 876
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3721
timestamp 0
transform 0 1 2544 -1 0 875
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3720
timestamp 0
transform 0 1 2544 -1 0 874
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3719
timestamp 0
transform 0 1 2544 -1 0 873
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3718
timestamp 0
transform 0 1 2544 -1 0 872
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3717
timestamp 0
transform 0 1 2544 -1 0 871
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3716
timestamp 0
transform 0 1 2544 -1 0 870
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3715
timestamp 0
transform 0 1 2544 -1 0 869
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3714
timestamp 0
transform 0 1 2544 -1 0 868
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3713
timestamp 0
transform 0 1 2544 -1 0 867
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3712
timestamp 0
transform 0 1 2544 -1 0 866
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3711
timestamp 0
transform 0 1 2544 -1 0 865
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3710
timestamp 0
transform 0 1 2544 -1 0 864
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3709
timestamp 0
transform 0 1 2544 -1 0 863
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3708
timestamp 0
transform 0 1 2544 -1 0 862
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3707
timestamp 0
transform 0 1 2544 -1 0 861
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3706
timestamp 0
transform 0 1 2544 -1 0 860
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3705
timestamp 0
transform 0 1 2544 -1 0 859
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3704
timestamp 0
transform 0 1 2544 -1 0 858
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3703
timestamp 0
transform 0 1 2544 -1 0 857
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3702
timestamp 0
transform 0 1 2544 -1 0 856
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3701
timestamp 0
transform 0 1 2544 -1 0 855
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3700
timestamp 0
transform 0 1 2544 -1 0 854
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3699
timestamp 0
transform 0 1 2544 -1 0 853
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3698
timestamp 0
transform 0 1 2544 -1 0 852
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3697
timestamp 0
transform 0 1 2544 -1 0 851
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3696
timestamp 0
transform 0 1 2544 -1 0 850
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3695
timestamp 0
transform 0 1 2544 -1 0 849
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3694
timestamp 0
transform 0 1 2544 -1 0 848
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3693
timestamp 0
transform 0 1 2544 -1 0 847
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3692
timestamp 0
transform 0 1 2544 -1 0 846
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3691
timestamp 0
transform 0 1 2544 -1 0 845
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3690
timestamp 0
transform 0 1 2544 -1 0 844
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3689
timestamp 0
transform 0 1 2544 -1 0 843
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3688
timestamp 0
transform 0 1 2544 -1 0 842
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3687
timestamp 0
transform 0 1 2544 -1 0 841
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3686
timestamp 0
transform 0 1 2544 -1 0 840
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3685
timestamp 0
transform 0 1 2544 -1 0 839
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3684
timestamp 0
transform 0 1 2544 -1 0 838
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3683
timestamp 0
transform 0 1 2544 -1 0 837
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3682
timestamp 0
transform 0 1 2544 -1 0 836
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3681
timestamp 0
transform 0 1 2544 -1 0 835
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3680
timestamp 0
transform 0 1 2544 -1 0 834
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3679
timestamp 0
transform 0 1 2544 -1 0 833
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3678
timestamp 0
transform 0 1 2544 -1 0 832
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3677
timestamp 0
transform 0 1 2544 -1 0 831
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3676
timestamp 0
transform 0 1 2544 -1 0 830
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3675
timestamp 0
transform 0 1 2544 -1 0 829
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3674
timestamp 0
transform 0 1 2544 -1 0 828
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3673
timestamp 0
transform 0 1 2544 -1 0 827
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3672
timestamp 0
transform 0 1 2544 -1 0 826
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3671
timestamp 0
transform 0 1 2544 -1 0 825
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3670
timestamp 0
transform 0 1 2544 -1 0 824
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3669
timestamp 0
transform 0 1 2544 -1 0 823
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3668
timestamp 0
transform 0 1 2544 -1 0 822
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3667
timestamp 0
transform 0 1 2544 -1 0 821
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3666
timestamp 0
transform 0 1 2544 -1 0 820
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3665
timestamp 0
transform 0 1 2544 -1 0 819
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3664
timestamp 0
transform 0 1 2544 -1 0 818
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3663
timestamp 0
transform 0 1 2544 -1 0 817
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3662
timestamp 0
transform 0 1 2544 -1 0 816
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3661
timestamp 0
transform 0 1 2544 -1 0 815
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3660
timestamp 0
transform 0 1 2544 -1 0 814
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3659
timestamp 0
transform 0 1 2544 -1 0 813
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3658
timestamp 0
transform 0 1 2544 -1 0 812
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3657
timestamp 0
transform 0 1 2544 -1 0 811
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3656
timestamp 0
transform 0 1 2544 -1 0 810
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3655
timestamp 0
transform 0 1 2544 -1 0 809
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3654
timestamp 0
transform 0 1 2544 -1 0 808
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3653
timestamp 0
transform 0 1 2544 -1 0 807
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3652
timestamp 0
transform 0 1 2544 -1 0 806
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3651
timestamp 0
transform 0 1 2544 -1 0 805
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3650
timestamp 0
transform 0 1 2544 -1 0 804
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3649
timestamp 0
transform 0 1 2544 -1 0 803
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3648
timestamp 0
transform 0 1 2544 -1 0 802
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3647
timestamp 0
transform 0 1 2544 -1 0 801
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3646
timestamp 0
transform 0 1 2544 -1 0 800
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3645
timestamp 0
transform 0 1 2544 -1 0 799
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3644
timestamp 0
transform 0 1 2544 -1 0 798
box 0 0 1 1
use s8iom0_vccd_hvc_pad  vdd1v8hclamp[1]
timestamp 0
transform 0 1 2544 -1 0 797
box 0 0 1 1
use s8iom0_gpiov2_pad  comp_inp_pad
timestamp 0
transform 0 -1 198 1 0 789
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2570
timestamp 0
transform 0 -1 198 1 0 788
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2569
timestamp 0
transform 0 -1 198 1 0 787
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2568
timestamp 0
transform 0 -1 198 1 0 786
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2567
timestamp 0
transform 0 -1 198 1 0 785
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2566
timestamp 0
transform 0 -1 198 1 0 784
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2565
timestamp 0
transform 0 -1 198 1 0 783
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2564
timestamp 0
transform 0 -1 198 1 0 782
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2563
timestamp 0
transform 0 -1 198 1 0 781
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2562
timestamp 0
transform 0 -1 198 1 0 780
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2561
timestamp 0
transform 0 -1 198 1 0 779
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2560
timestamp 0
transform 0 -1 198 1 0 778
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2559
timestamp 0
transform 0 -1 198 1 0 777
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2558
timestamp 0
transform 0 -1 198 1 0 776
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2557
timestamp 0
transform 0 -1 198 1 0 775
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2556
timestamp 0
transform 0 -1 198 1 0 774
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2555
timestamp 0
transform 0 -1 198 1 0 773
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2554
timestamp 0
transform 0 -1 198 1 0 772
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2553
timestamp 0
transform 0 -1 198 1 0 771
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2552
timestamp 0
transform 0 -1 198 1 0 770
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2551
timestamp 0
transform 0 -1 198 1 0 769
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2550
timestamp 0
transform 0 -1 198 1 0 768
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2549
timestamp 0
transform 0 -1 198 1 0 767
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2548
timestamp 0
transform 0 -1 198 1 0 766
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2547
timestamp 0
transform 0 -1 198 1 0 765
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2546
timestamp 0
transform 0 -1 198 1 0 764
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2545
timestamp 0
transform 0 -1 198 1 0 763
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2544
timestamp 0
transform 0 -1 198 1 0 762
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2543
timestamp 0
transform 0 -1 198 1 0 761
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2542
timestamp 0
transform 0 -1 198 1 0 760
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2541
timestamp 0
transform 0 -1 198 1 0 759
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2540
timestamp 0
transform 0 -1 198 1 0 758
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2539
timestamp 0
transform 0 -1 198 1 0 757
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2538
timestamp 0
transform 0 -1 198 1 0 756
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2537
timestamp 0
transform 0 -1 198 1 0 755
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2536
timestamp 0
transform 0 -1 198 1 0 754
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2535
timestamp 0
transform 0 -1 198 1 0 753
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2534
timestamp 0
transform 0 -1 198 1 0 752
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2533
timestamp 0
transform 0 -1 198 1 0 751
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2532
timestamp 0
transform 0 -1 198 1 0 750
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2531
timestamp 0
transform 0 -1 198 1 0 749
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2530
timestamp 0
transform 0 -1 198 1 0 748
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2529
timestamp 0
transform 0 -1 198 1 0 747
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2528
timestamp 0
transform 0 -1 198 1 0 746
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2527
timestamp 0
transform 0 -1 198 1 0 745
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2526
timestamp 0
transform 0 -1 198 1 0 744
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2525
timestamp 0
transform 0 -1 198 1 0 743
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2524
timestamp 0
transform 0 -1 198 1 0 742
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2523
timestamp 0
transform 0 -1 198 1 0 741
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2522
timestamp 0
transform 0 -1 198 1 0 740
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2521
timestamp 0
transform 0 -1 198 1 0 739
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2520
timestamp 0
transform 0 -1 198 1 0 738
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2519
timestamp 0
transform 0 -1 198 1 0 737
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2518
timestamp 0
transform 0 -1 198 1 0 736
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2517
timestamp 0
transform 0 -1 198 1 0 735
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2516
timestamp 0
transform 0 -1 198 1 0 734
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2515
timestamp 0
transform 0 -1 198 1 0 733
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2514
timestamp 0
transform 0 -1 198 1 0 732
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3642
timestamp 0
transform 0 1 2544 -1 0 722
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3641
timestamp 0
transform 0 1 2544 -1 0 721
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3640
timestamp 0
transform 0 1 2544 -1 0 720
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3639
timestamp 0
transform 0 1 2544 -1 0 719
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3638
timestamp 0
transform 0 1 2544 -1 0 718
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3637
timestamp 0
transform 0 1 2544 -1 0 717
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3636
timestamp 0
transform 0 1 2544 -1 0 716
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3635
timestamp 0
transform 0 1 2544 -1 0 715
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3634
timestamp 0
transform 0 1 2544 -1 0 714
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3633
timestamp 0
transform 0 1 2544 -1 0 713
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3632
timestamp 0
transform 0 1 2544 -1 0 712
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3631
timestamp 0
transform 0 1 2544 -1 0 711
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3630
timestamp 0
transform 0 1 2544 -1 0 710
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3629
timestamp 0
transform 0 1 2544 -1 0 709
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3628
timestamp 0
transform 0 1 2544 -1 0 708
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3627
timestamp 0
transform 0 1 2544 -1 0 707
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3626
timestamp 0
transform 0 1 2544 -1 0 706
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3625
timestamp 0
transform 0 1 2544 -1 0 705
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3624
timestamp 0
transform 0 1 2544 -1 0 704
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3623
timestamp 0
transform 0 1 2544 -1 0 703
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3622
timestamp 0
transform 0 1 2544 -1 0 702
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3621
timestamp 0
transform 0 1 2544 -1 0 701
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3620
timestamp 0
transform 0 1 2544 -1 0 700
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3619
timestamp 0
transform 0 1 2544 -1 0 699
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3618
timestamp 0
transform 0 1 2544 -1 0 698
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3617
timestamp 0
transform 0 1 2544 -1 0 697
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3616
timestamp 0
transform 0 1 2544 -1 0 696
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3615
timestamp 0
transform 0 1 2544 -1 0 695
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3614
timestamp 0
transform 0 1 2544 -1 0 694
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3613
timestamp 0
transform 0 1 2544 -1 0 693
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3612
timestamp 0
transform 0 1 2544 -1 0 692
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3611
timestamp 0
transform 0 1 2544 -1 0 691
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3610
timestamp 0
transform 0 1 2544 -1 0 690
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3609
timestamp 0
transform 0 1 2544 -1 0 689
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3608
timestamp 0
transform 0 1 2544 -1 0 688
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3607
timestamp 0
transform 0 1 2544 -1 0 687
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3606
timestamp 0
transform 0 1 2544 -1 0 686
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3605
timestamp 0
transform 0 1 2544 -1 0 685
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3604
timestamp 0
transform 0 1 2544 -1 0 684
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3603
timestamp 0
transform 0 1 2544 -1 0 683
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3602
timestamp 0
transform 0 1 2544 -1 0 682
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3601
timestamp 0
transform 0 1 2544 -1 0 681
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3600
timestamp 0
transform 0 1 2544 -1 0 680
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3599
timestamp 0
transform 0 1 2544 -1 0 679
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3598
timestamp 0
transform 0 1 2544 -1 0 678
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3597
timestamp 0
transform 0 1 2544 -1 0 677
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3596
timestamp 0
transform 0 1 2544 -1 0 676
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3595
timestamp 0
transform 0 1 2544 -1 0 675
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3594
timestamp 0
transform 0 1 2544 -1 0 674
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3593
timestamp 0
transform 0 1 2544 -1 0 673
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3592
timestamp 0
transform 0 1 2544 -1 0 672
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3591
timestamp 0
transform 0 1 2544 -1 0 671
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3590
timestamp 0
transform 0 1 2544 -1 0 670
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3589
timestamp 0
transform 0 1 2544 -1 0 669
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3588
timestamp 0
transform 0 1 2544 -1 0 668
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3587
timestamp 0
transform 0 1 2544 -1 0 667
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3586
timestamp 0
transform 0 1 2544 -1 0 666
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3585
timestamp 0
transform 0 1 2544 -1 0 665
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3584
timestamp 0
transform 0 1 2544 -1 0 664
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3583
timestamp 0
transform 0 1 2544 -1 0 663
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3582
timestamp 0
transform 0 1 2544 -1 0 662
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3581
timestamp 0
transform 0 1 2544 -1 0 661
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3580
timestamp 0
transform 0 1 2544 -1 0 660
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3579
timestamp 0
transform 0 1 2544 -1 0 659
box 0 0 1 1
use s8iom0_vssa_hvc_pad  vsshclamp[2]
timestamp 0
transform 0 -1 198 1 0 657
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2512
timestamp 0
transform 0 -1 198 1 0 656
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2511
timestamp 0
transform 0 -1 198 1 0 655
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2510
timestamp 0
transform 0 -1 198 1 0 654
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2509
timestamp 0
transform 0 -1 198 1 0 653
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2508
timestamp 0
transform 0 -1 198 1 0 652
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2507
timestamp 0
transform 0 -1 198 1 0 651
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2506
timestamp 0
transform 0 -1 198 1 0 650
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2505
timestamp 0
transform 0 -1 198 1 0 649
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2504
timestamp 0
transform 0 -1 198 1 0 648
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2503
timestamp 0
transform 0 -1 198 1 0 647
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2502
timestamp 0
transform 0 -1 198 1 0 646
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2501
timestamp 0
transform 0 -1 198 1 0 645
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2500
timestamp 0
transform 0 -1 198 1 0 644
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2499
timestamp 0
transform 0 -1 198 1 0 643
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2498
timestamp 0
transform 0 -1 198 1 0 642
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2497
timestamp 0
transform 0 -1 198 1 0 641
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2496
timestamp 0
transform 0 -1 198 1 0 640
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2495
timestamp 0
transform 0 -1 198 1 0 639
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2494
timestamp 0
transform 0 -1 198 1 0 638
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2493
timestamp 0
transform 0 -1 198 1 0 637
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2492
timestamp 0
transform 0 -1 198 1 0 636
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2491
timestamp 0
transform 0 -1 198 1 0 635
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2490
timestamp 0
transform 0 -1 198 1 0 634
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2489
timestamp 0
transform 0 -1 198 1 0 633
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2488
timestamp 0
transform 0 -1 198 1 0 632
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2487
timestamp 0
transform 0 -1 198 1 0 631
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2486
timestamp 0
transform 0 -1 198 1 0 630
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2485
timestamp 0
transform 0 -1 198 1 0 629
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2484
timestamp 0
transform 0 -1 198 1 0 628
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2483
timestamp 0
transform 0 -1 198 1 0 627
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2482
timestamp 0
transform 0 -1 198 1 0 626
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2481
timestamp 0
transform 0 -1 198 1 0 625
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2480
timestamp 0
transform 0 -1 198 1 0 624
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2479
timestamp 0
transform 0 -1 198 1 0 623
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2478
timestamp 0
transform 0 -1 198 1 0 622
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2477
timestamp 0
transform 0 -1 198 1 0 621
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2476
timestamp 0
transform 0 -1 198 1 0 620
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2475
timestamp 0
transform 0 -1 198 1 0 619
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2474
timestamp 0
transform 0 -1 198 1 0 618
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2473
timestamp 0
transform 0 -1 198 1 0 617
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2472
timestamp 0
transform 0 -1 198 1 0 616
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2471
timestamp 0
transform 0 -1 198 1 0 615
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2470
timestamp 0
transform 0 -1 198 1 0 614
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2469
timestamp 0
transform 0 -1 198 1 0 613
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2468
timestamp 0
transform 0 -1 198 1 0 612
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2467
timestamp 0
transform 0 -1 198 1 0 611
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2466
timestamp 0
transform 0 -1 198 1 0 610
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2465
timestamp 0
transform 0 -1 198 1 0 609
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2464
timestamp 0
transform 0 -1 198 1 0 608
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2463
timestamp 0
transform 0 -1 198 1 0 607
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2462
timestamp 0
transform 0 -1 198 1 0 606
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2461
timestamp 0
transform 0 -1 198 1 0 605
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2460
timestamp 0
transform 0 -1 198 1 0 604
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2459
timestamp 0
transform 0 -1 198 1 0 603
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2458
timestamp 0
transform 0 -1 198 1 0 602
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2457
timestamp 0
transform 0 -1 198 1 0 601
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2456
timestamp 0
transform 0 -1 198 1 0 600
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3578
timestamp 0
transform 0 1 2544 -1 0 658
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3577
timestamp 0
transform 0 1 2544 -1 0 657
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3576
timestamp 0
transform 0 1 2544 -1 0 656
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3575
timestamp 0
transform 0 1 2544 -1 0 655
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3574
timestamp 0
transform 0 1 2544 -1 0 654
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3573
timestamp 0
transform 0 1 2544 -1 0 653
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3572
timestamp 0
transform 0 1 2544 -1 0 652
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3571
timestamp 0
transform 0 1 2544 -1 0 651
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3570
timestamp 0
transform 0 1 2544 -1 0 650
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3569
timestamp 0
transform 0 1 2544 -1 0 649
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3568
timestamp 0
transform 0 1 2544 -1 0 648
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3567
timestamp 0
transform 0 1 2544 -1 0 647
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3566
timestamp 0
transform 0 1 2544 -1 0 646
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3565
timestamp 0
transform 0 1 2544 -1 0 645
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3564
timestamp 0
transform 0 1 2544 -1 0 644
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3563
timestamp 0
transform 0 1 2544 -1 0 643
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3562
timestamp 0
transform 0 1 2544 -1 0 642
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3561
timestamp 0
transform 0 1 2544 -1 0 641
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3560
timestamp 0
transform 0 1 2544 -1 0 640
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3559
timestamp 0
transform 0 1 2544 -1 0 639
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3558
timestamp 0
transform 0 1 2544 -1 0 638
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3557
timestamp 0
transform 0 1 2544 -1 0 637
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3556
timestamp 0
transform 0 1 2544 -1 0 636
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3555
timestamp 0
transform 0 1 2544 -1 0 635
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3554
timestamp 0
transform 0 1 2544 -1 0 634
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3553
timestamp 0
transform 0 1 2544 -1 0 633
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3552
timestamp 0
transform 0 1 2544 -1 0 632
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3551
timestamp 0
transform 0 1 2544 -1 0 631
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3550
timestamp 0
transform 0 1 2544 -1 0 630
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3549
timestamp 0
transform 0 1 2544 -1 0 629
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3548
timestamp 0
transform 0 1 2544 -1 0 628
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3547
timestamp 0
transform 0 1 2544 -1 0 627
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3546
timestamp 0
transform 0 1 2544 -1 0 626
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3545
timestamp 0
transform 0 1 2544 -1 0 625
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3544
timestamp 0
transform 0 1 2544 -1 0 624
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3543
timestamp 0
transform 0 1 2544 -1 0 623
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3542
timestamp 0
transform 0 1 2544 -1 0 622
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3541
timestamp 0
transform 0 1 2544 -1 0 621
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3540
timestamp 0
transform 0 1 2544 -1 0 620
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3539
timestamp 0
transform 0 1 2544 -1 0 619
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3538
timestamp 0
transform 0 1 2544 -1 0 618
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3537
timestamp 0
transform 0 1 2544 -1 0 617
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3536
timestamp 0
transform 0 1 2544 -1 0 616
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3535
timestamp 0
transform 0 1 2544 -1 0 615
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3534
timestamp 0
transform 0 1 2544 -1 0 614
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3533
timestamp 0
transform 0 1 2544 -1 0 613
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3532
timestamp 0
transform 0 1 2544 -1 0 612
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3531
timestamp 0
transform 0 1 2544 -1 0 611
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3530
timestamp 0
transform 0 1 2544 -1 0 610
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3529
timestamp 0
transform 0 1 2544 -1 0 609
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3528
timestamp 0
transform 0 1 2544 -1 0 608
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3527
timestamp 0
transform 0 1 2544 -1 0 607
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3526
timestamp 0
transform 0 1 2544 -1 0 606
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3525
timestamp 0
transform 0 1 2544 -1 0 605
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3524
timestamp 0
transform 0 1 2544 -1 0 604
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3523
timestamp 0
transform 0 1 2544 -1 0 603
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3522
timestamp 0
transform 0 1 2544 -1 0 602
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3521
timestamp 0
transform 0 1 2544 -1 0 601
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3520
timestamp 0
transform 0 1 2544 -1 0 600
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3519
timestamp 0
transform 0 1 2544 -1 0 599
box 0 0 1 1
use s8iom0_vdda_lvc_pad  vdd3v3lclamp[1]
timestamp 0
transform 0 1 2544 -1 0 598
box 0 0 1 1
use s8iom0_vccd_lvc_pad  vdd1v8lclamp[1]
timestamp 0
transform 0 -1 198 1 0 525
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2454
timestamp 0
transform 0 -1 198 1 0 524
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2453
timestamp 0
transform 0 -1 198 1 0 523
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2452
timestamp 0
transform 0 -1 198 1 0 522
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2451
timestamp 0
transform 0 -1 198 1 0 521
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2450
timestamp 0
transform 0 -1 198 1 0 520
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2449
timestamp 0
transform 0 -1 198 1 0 519
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2448
timestamp 0
transform 0 -1 198 1 0 518
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2447
timestamp 0
transform 0 -1 198 1 0 517
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2446
timestamp 0
transform 0 -1 198 1 0 516
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2445
timestamp 0
transform 0 -1 198 1 0 515
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2444
timestamp 0
transform 0 -1 198 1 0 514
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2443
timestamp 0
transform 0 -1 198 1 0 513
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2442
timestamp 0
transform 0 -1 198 1 0 512
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2441
timestamp 0
transform 0 -1 198 1 0 511
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2440
timestamp 0
transform 0 -1 198 1 0 510
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2439
timestamp 0
transform 0 -1 198 1 0 509
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2438
timestamp 0
transform 0 -1 198 1 0 508
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2437
timestamp 0
transform 0 -1 198 1 0 507
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2436
timestamp 0
transform 0 -1 198 1 0 506
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2435
timestamp 0
transform 0 -1 198 1 0 505
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2434
timestamp 0
transform 0 -1 198 1 0 504
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2433
timestamp 0
transform 0 -1 198 1 0 503
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2432
timestamp 0
transform 0 -1 198 1 0 502
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2431
timestamp 0
transform 0 -1 198 1 0 501
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2430
timestamp 0
transform 0 -1 198 1 0 500
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2429
timestamp 0
transform 0 -1 198 1 0 499
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2428
timestamp 0
transform 0 -1 198 1 0 498
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2427
timestamp 0
transform 0 -1 198 1 0 497
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2426
timestamp 0
transform 0 -1 198 1 0 496
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2425
timestamp 0
transform 0 -1 198 1 0 495
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2424
timestamp 0
transform 0 -1 198 1 0 494
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2423
timestamp 0
transform 0 -1 198 1 0 493
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2422
timestamp 0
transform 0 -1 198 1 0 492
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2421
timestamp 0
transform 0 -1 198 1 0 491
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2420
timestamp 0
transform 0 -1 198 1 0 490
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2419
timestamp 0
transform 0 -1 198 1 0 489
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2418
timestamp 0
transform 0 -1 198 1 0 488
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2417
timestamp 0
transform 0 -1 198 1 0 487
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2416
timestamp 0
transform 0 -1 198 1 0 486
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2415
timestamp 0
transform 0 -1 198 1 0 485
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2414
timestamp 0
transform 0 -1 198 1 0 484
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2413
timestamp 0
transform 0 -1 198 1 0 483
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2412
timestamp 0
transform 0 -1 198 1 0 482
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2411
timestamp 0
transform 0 -1 198 1 0 481
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2410
timestamp 0
transform 0 -1 198 1 0 480
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2409
timestamp 0
transform 0 -1 198 1 0 479
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2408
timestamp 0
transform 0 -1 198 1 0 478
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2407
timestamp 0
transform 0 -1 198 1 0 477
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2406
timestamp 0
transform 0 -1 198 1 0 476
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2405
timestamp 0
transform 0 -1 198 1 0 475
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2404
timestamp 0
transform 0 -1 198 1 0 474
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2403
timestamp 0
transform 0 -1 198 1 0 473
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2402
timestamp 0
transform 0 -1 198 1 0 472
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2401
timestamp 0
transform 0 -1 198 1 0 471
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2400
timestamp 0
transform 0 -1 198 1 0 470
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2399
timestamp 0
transform 0 -1 198 1 0 469
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2398
timestamp 0
transform 0 -1 198 1 0 468
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3517
timestamp 0
transform 0 1 2544 -1 0 523
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3516
timestamp 0
transform 0 1 2544 -1 0 522
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3515
timestamp 0
transform 0 1 2544 -1 0 521
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3514
timestamp 0
transform 0 1 2544 -1 0 520
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3513
timestamp 0
transform 0 1 2544 -1 0 519
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3512
timestamp 0
transform 0 1 2544 -1 0 518
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3511
timestamp 0
transform 0 1 2544 -1 0 517
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3510
timestamp 0
transform 0 1 2544 -1 0 516
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3509
timestamp 0
transform 0 1 2544 -1 0 515
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3508
timestamp 0
transform 0 1 2544 -1 0 514
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3507
timestamp 0
transform 0 1 2544 -1 0 513
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3506
timestamp 0
transform 0 1 2544 -1 0 512
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3505
timestamp 0
transform 0 1 2544 -1 0 511
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3504
timestamp 0
transform 0 1 2544 -1 0 510
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3503
timestamp 0
transform 0 1 2544 -1 0 509
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3502
timestamp 0
transform 0 1 2544 -1 0 508
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3501
timestamp 0
transform 0 1 2544 -1 0 507
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3500
timestamp 0
transform 0 1 2544 -1 0 506
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3499
timestamp 0
transform 0 1 2544 -1 0 505
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3498
timestamp 0
transform 0 1 2544 -1 0 504
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3497
timestamp 0
transform 0 1 2544 -1 0 503
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3496
timestamp 0
transform 0 1 2544 -1 0 502
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3495
timestamp 0
transform 0 1 2544 -1 0 501
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3494
timestamp 0
transform 0 1 2544 -1 0 500
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3493
timestamp 0
transform 0 1 2544 -1 0 499
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3492
timestamp 0
transform 0 1 2544 -1 0 498
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3491
timestamp 0
transform 0 1 2544 -1 0 497
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3490
timestamp 0
transform 0 1 2544 -1 0 496
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3489
timestamp 0
transform 0 1 2544 -1 0 495
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3488
timestamp 0
transform 0 1 2544 -1 0 494
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3487
timestamp 0
transform 0 1 2544 -1 0 493
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3486
timestamp 0
transform 0 1 2544 -1 0 492
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3485
timestamp 0
transform 0 1 2544 -1 0 491
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3484
timestamp 0
transform 0 1 2544 -1 0 490
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3483
timestamp 0
transform 0 1 2544 -1 0 489
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3482
timestamp 0
transform 0 1 2544 -1 0 488
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3481
timestamp 0
transform 0 1 2544 -1 0 487
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3480
timestamp 0
transform 0 1 2544 -1 0 486
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3479
timestamp 0
transform 0 1 2544 -1 0 485
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3478
timestamp 0
transform 0 1 2544 -1 0 484
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3477
timestamp 0
transform 0 1 2544 -1 0 483
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3476
timestamp 0
transform 0 1 2544 -1 0 482
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3475
timestamp 0
transform 0 1 2544 -1 0 481
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3474
timestamp 0
transform 0 1 2544 -1 0 480
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3473
timestamp 0
transform 0 1 2544 -1 0 479
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3472
timestamp 0
transform 0 1 2544 -1 0 478
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3471
timestamp 0
transform 0 1 2544 -1 0 477
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3470
timestamp 0
transform 0 1 2544 -1 0 476
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3469
timestamp 0
transform 0 1 2544 -1 0 475
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3468
timestamp 0
transform 0 1 2544 -1 0 474
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3467
timestamp 0
transform 0 1 2544 -1 0 473
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3466
timestamp 0
transform 0 1 2544 -1 0 472
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3465
timestamp 0
transform 0 1 2544 -1 0 471
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3464
timestamp 0
transform 0 1 2544 -1 0 470
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3463
timestamp 0
transform 0 1 2544 -1 0 469
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3462
timestamp 0
transform 0 1 2544 -1 0 468
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3461
timestamp 0
transform 0 1 2544 -1 0 467
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3460
timestamp 0
transform 0 1 2544 -1 0 466
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3459
timestamp 0
transform 0 1 2544 -1 0 465
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3458
timestamp 0
transform 0 1 2544 -1 0 464
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3457
timestamp 0
transform 0 1 2544 -1 0 463
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3456
timestamp 0
transform 0 1 2544 -1 0 462
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3455
timestamp 0
transform 0 1 2544 -1 0 461
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3454
timestamp 0
transform 0 1 2544 -1 0 460
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3453
timestamp 0
transform 0 1 2544 -1 0 459
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3452
timestamp 0
transform 0 1 2544 -1 0 458
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3451
timestamp 0
transform 0 1 2544 -1 0 457
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3450
timestamp 0
transform 0 1 2544 -1 0 456
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3449
timestamp 0
transform 0 1 2544 -1 0 455
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3448
timestamp 0
transform 0 1 2544 -1 0 454
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3447
timestamp 0
transform 0 1 2544 -1 0 453
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3446
timestamp 0
transform 0 1 2544 -1 0 452
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3445
timestamp 0
transform 0 1 2544 -1 0 451
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3444
timestamp 0
transform 0 1 2544 -1 0 450
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3443
timestamp 0
transform 0 1 2544 -1 0 449
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3442
timestamp 0
transform 0 1 2544 -1 0 448
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3441
timestamp 0
transform 0 1 2544 -1 0 447
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3440
timestamp 0
transform 0 1 2544 -1 0 446
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3439
timestamp 0
transform 0 1 2544 -1 0 445
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3438
timestamp 0
transform 0 1 2544 -1 0 444
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3437
timestamp 0
transform 0 1 2544 -1 0 443
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3436
timestamp 0
transform 0 1 2544 -1 0 442
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3435
timestamp 0
transform 0 1 2544 -1 0 441
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3434
timestamp 0
transform 0 1 2544 -1 0 440
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3433
timestamp 0
transform 0 1 2544 -1 0 439
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3432
timestamp 0
transform 0 1 2544 -1 0 438
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3431
timestamp 0
transform 0 1 2544 -1 0 437
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3430
timestamp 0
transform 0 1 2544 -1 0 436
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3429
timestamp 0
transform 0 1 2544 -1 0 435
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3428
timestamp 0
transform 0 1 2544 -1 0 434
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3427
timestamp 0
transform 0 1 2544 -1 0 433
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3426
timestamp 0
transform 0 1 2544 -1 0 432
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3425
timestamp 0
transform 0 1 2544 -1 0 431
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3424
timestamp 0
transform 0 1 2544 -1 0 430
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3423
timestamp 0
transform 0 1 2544 -1 0 429
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3422
timestamp 0
transform 0 1 2544 -1 0 428
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3421
timestamp 0
transform 0 1 2544 -1 0 427
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3420
timestamp 0
transform 0 1 2544 -1 0 426
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3419
timestamp 0
transform 0 1 2544 -1 0 425
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3418
timestamp 0
transform 0 1 2544 -1 0 424
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3417
timestamp 0
transform 0 1 2544 -1 0 423
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3416
timestamp 0
transform 0 1 2544 -1 0 422
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3415
timestamp 0
transform 0 1 2544 -1 0 421
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3414
timestamp 0
transform 0 1 2544 -1 0 420
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3413
timestamp 0
transform 0 1 2544 -1 0 419
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3412
timestamp 0
transform 0 1 2544 -1 0 418
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3411
timestamp 0
transform 0 1 2544 -1 0 417
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3410
timestamp 0
transform 0 1 2544 -1 0 416
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3409
timestamp 0
transform 0 1 2544 -1 0 415
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3408
timestamp 0
transform 0 1 2544 -1 0 414
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3407
timestamp 0
transform 0 1 2544 -1 0 413
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3406
timestamp 0
transform 0 1 2544 -1 0 412
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3405
timestamp 0
transform 0 1 2544 -1 0 411
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3404
timestamp 0
transform 0 1 2544 -1 0 410
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3403
timestamp 0
transform 0 1 2544 -1 0 409
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3402
timestamp 0
transform 0 1 2544 -1 0 408
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3401
timestamp 0
transform 0 1 2544 -1 0 407
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3400
timestamp 0
transform 0 1 2544 -1 0 406
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3399
timestamp 0
transform 0 1 2544 -1 0 405
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3398
timestamp 0
transform 0 1 2544 -1 0 404
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3397
timestamp 0
transform 0 1 2544 -1 0 403
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3396
timestamp 0
transform 0 1 2544 -1 0 402
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3395
timestamp 0
transform 0 1 2544 -1 0 401
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3394
timestamp 0
transform 0 1 2544 -1 0 400
box 0 0 1 1
use s8iom0_vdda_hvc_pad  vdd3v3hclamp[1]
timestamp 0
transform 0 1 2544 -1 0 399
box 0 0 1 1
use s8iom0_vdda_lvc_pad  vdd3v3lclamp[3]
timestamp 0
transform 0 -1 198 1 0 393
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2396
timestamp 0
transform 0 -1 198 1 0 392
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2395
timestamp 0
transform 0 -1 198 1 0 391
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2394
timestamp 0
transform 0 -1 198 1 0 390
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2393
timestamp 0
transform 0 -1 198 1 0 389
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2392
timestamp 0
transform 0 -1 198 1 0 388
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2391
timestamp 0
transform 0 -1 198 1 0 387
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2390
timestamp 0
transform 0 -1 198 1 0 386
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2389
timestamp 0
transform 0 -1 198 1 0 385
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2388
timestamp 0
transform 0 -1 198 1 0 384
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2387
timestamp 0
transform 0 -1 198 1 0 383
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2386
timestamp 0
transform 0 -1 198 1 0 382
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2385
timestamp 0
transform 0 -1 198 1 0 381
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2384
timestamp 0
transform 0 -1 198 1 0 380
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2383
timestamp 0
transform 0 -1 198 1 0 379
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2382
timestamp 0
transform 0 -1 198 1 0 378
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2381
timestamp 0
transform 0 -1 198 1 0 377
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2380
timestamp 0
transform 0 -1 198 1 0 376
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2379
timestamp 0
transform 0 -1 198 1 0 375
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2378
timestamp 0
transform 0 -1 198 1 0 374
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2377
timestamp 0
transform 0 -1 198 1 0 373
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2376
timestamp 0
transform 0 -1 198 1 0 372
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2375
timestamp 0
transform 0 -1 198 1 0 371
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2374
timestamp 0
transform 0 -1 198 1 0 370
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2373
timestamp 0
transform 0 -1 198 1 0 369
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2372
timestamp 0
transform 0 -1 198 1 0 368
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2371
timestamp 0
transform 0 -1 198 1 0 367
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2370
timestamp 0
transform 0 -1 198 1 0 366
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2369
timestamp 0
transform 0 -1 198 1 0 365
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2368
timestamp 0
transform 0 -1 198 1 0 364
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2367
timestamp 0
transform 0 -1 198 1 0 363
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2366
timestamp 0
transform 0 -1 198 1 0 362
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2365
timestamp 0
transform 0 -1 198 1 0 361
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2364
timestamp 0
transform 0 -1 198 1 0 360
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2363
timestamp 0
transform 0 -1 198 1 0 359
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2362
timestamp 0
transform 0 -1 198 1 0 358
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2361
timestamp 0
transform 0 -1 198 1 0 357
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2360
timestamp 0
transform 0 -1 198 1 0 356
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2359
timestamp 0
transform 0 -1 198 1 0 355
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2358
timestamp 0
transform 0 -1 198 1 0 354
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2357
timestamp 0
transform 0 -1 198 1 0 353
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2356
timestamp 0
transform 0 -1 198 1 0 352
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2355
timestamp 0
transform 0 -1 198 1 0 351
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2354
timestamp 0
transform 0 -1 198 1 0 350
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2353
timestamp 0
transform 0 -1 198 1 0 349
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2352
timestamp 0
transform 0 -1 198 1 0 348
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2351
timestamp 0
transform 0 -1 198 1 0 347
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2350
timestamp 0
transform 0 -1 198 1 0 346
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2349
timestamp 0
transform 0 -1 198 1 0 345
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2348
timestamp 0
transform 0 -1 198 1 0 344
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2347
timestamp 0
transform 0 -1 198 1 0 343
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2346
timestamp 0
transform 0 -1 198 1 0 342
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2345
timestamp 0
transform 0 -1 198 1 0 341
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2344
timestamp 0
transform 0 -1 198 1 0 340
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2343
timestamp 0
transform 0 -1 198 1 0 339
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2342
timestamp 0
transform 0 -1 198 1 0 338
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2341
timestamp 0
transform 0 -1 198 1 0 337
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2340
timestamp 0
transform 0 -1 198 1 0 336
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3392
timestamp 0
transform 0 1 2544 -1 0 324
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3391
timestamp 0
transform 0 1 2544 -1 0 323
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3390
timestamp 0
transform 0 1 2544 -1 0 322
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3389
timestamp 0
transform 0 1 2544 -1 0 321
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3388
timestamp 0
transform 0 1 2544 -1 0 320
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3387
timestamp 0
transform 0 1 2544 -1 0 319
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3386
timestamp 0
transform 0 1 2544 -1 0 318
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3385
timestamp 0
transform 0 1 2544 -1 0 317
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3384
timestamp 0
transform 0 1 2544 -1 0 316
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3383
timestamp 0
transform 0 1 2544 -1 0 315
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3382
timestamp 0
transform 0 1 2544 -1 0 314
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3381
timestamp 0
transform 0 1 2544 -1 0 313
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3380
timestamp 0
transform 0 1 2544 -1 0 312
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3379
timestamp 0
transform 0 1 2544 -1 0 311
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3378
timestamp 0
transform 0 1 2544 -1 0 310
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3377
timestamp 0
transform 0 1 2544 -1 0 309
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3376
timestamp 0
transform 0 1 2544 -1 0 308
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3375
timestamp 0
transform 0 1 2544 -1 0 307
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3374
timestamp 0
transform 0 1 2544 -1 0 306
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3373
timestamp 0
transform 0 1 2544 -1 0 305
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3372
timestamp 0
transform 0 1 2544 -1 0 304
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3371
timestamp 0
transform 0 1 2544 -1 0 303
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3370
timestamp 0
transform 0 1 2544 -1 0 302
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3369
timestamp 0
transform 0 1 2544 -1 0 301
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3368
timestamp 0
transform 0 1 2544 -1 0 300
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3367
timestamp 0
transform 0 1 2544 -1 0 299
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3366
timestamp 0
transform 0 1 2544 -1 0 298
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3365
timestamp 0
transform 0 1 2544 -1 0 297
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3364
timestamp 0
transform 0 1 2544 -1 0 296
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3363
timestamp 0
transform 0 1 2544 -1 0 295
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3362
timestamp 0
transform 0 1 2544 -1 0 294
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3361
timestamp 0
transform 0 1 2544 -1 0 293
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3360
timestamp 0
transform 0 1 2544 -1 0 292
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3359
timestamp 0
transform 0 1 2544 -1 0 291
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3358
timestamp 0
transform 0 1 2544 -1 0 290
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3357
timestamp 0
transform 0 1 2544 -1 0 289
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3356
timestamp 0
transform 0 1 2544 -1 0 288
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3355
timestamp 0
transform 0 1 2544 -1 0 287
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3354
timestamp 0
transform 0 1 2544 -1 0 286
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3353
timestamp 0
transform 0 1 2544 -1 0 285
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3352
timestamp 0
transform 0 1 2544 -1 0 284
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3351
timestamp 0
transform 0 1 2544 -1 0 283
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3350
timestamp 0
transform 0 1 2544 -1 0 282
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3349
timestamp 0
transform 0 1 2544 -1 0 281
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3348
timestamp 0
transform 0 1 2544 -1 0 280
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3347
timestamp 0
transform 0 1 2544 -1 0 279
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3346
timestamp 0
transform 0 1 2544 -1 0 278
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3345
timestamp 0
transform 0 1 2544 -1 0 277
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3344
timestamp 0
transform 0 1 2544 -1 0 276
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3343
timestamp 0
transform 0 1 2544 -1 0 275
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3342
timestamp 0
transform 0 1 2544 -1 0 274
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3341
timestamp 0
transform 0 1 2544 -1 0 273
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3340
timestamp 0
transform 0 1 2544 -1 0 272
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3339
timestamp 0
transform 0 1 2544 -1 0 271
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3338
timestamp 0
transform 0 1 2544 -1 0 270
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3337
timestamp 0
transform 0 1 2544 -1 0 269
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3336
timestamp 0
transform 0 1 2544 -1 0 268
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3335
timestamp 0
transform 0 1 2544 -1 0 267
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3334
timestamp 0
transform 0 1 2544 -1 0 266
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3333
timestamp 0
transform 0 1 2544 -1 0 265
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3332
timestamp 0
transform 0 1 2544 -1 0 264
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3331
timestamp 0
transform 0 1 2544 -1 0 263
box 0 0 1 1
use s8iom0_vdda_hvc_pad  vddiohclamp[1]
timestamp 0
transform 0 -1 198 1 0 261
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2338
timestamp 0
transform 0 -1 198 1 0 260
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2337
timestamp 0
transform 0 -1 198 1 0 259
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2336
timestamp 0
transform 0 -1 198 1 0 258
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2335
timestamp 0
transform 0 -1 198 1 0 257
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2334
timestamp 0
transform 0 -1 198 1 0 256
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2333
timestamp 0
transform 0 -1 198 1 0 255
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2332
timestamp 0
transform 0 -1 198 1 0 254
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2331
timestamp 0
transform 0 -1 198 1 0 253
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2330
timestamp 0
transform 0 -1 198 1 0 252
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2329
timestamp 0
transform 0 -1 198 1 0 251
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2328
timestamp 0
transform 0 -1 198 1 0 250
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2327
timestamp 0
transform 0 -1 198 1 0 249
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2326
timestamp 0
transform 0 -1 198 1 0 248
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2325
timestamp 0
transform 0 -1 198 1 0 247
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2324
timestamp 0
transform 0 -1 198 1 0 246
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2323
timestamp 0
transform 0 -1 198 1 0 245
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2322
timestamp 0
transform 0 -1 198 1 0 244
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2321
timestamp 0
transform 0 -1 198 1 0 243
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2320
timestamp 0
transform 0 -1 198 1 0 242
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2319
timestamp 0
transform 0 -1 198 1 0 241
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2318
timestamp 0
transform 0 -1 198 1 0 240
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2317
timestamp 0
transform 0 -1 198 1 0 239
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2316
timestamp 0
transform 0 -1 198 1 0 238
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2315
timestamp 0
transform 0 -1 198 1 0 237
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2314
timestamp 0
transform 0 -1 198 1 0 236
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2313
timestamp 0
transform 0 -1 198 1 0 235
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2312
timestamp 0
transform 0 -1 198 1 0 234
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2311
timestamp 0
transform 0 -1 198 1 0 233
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2310
timestamp 0
transform 0 -1 198 1 0 232
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2309
timestamp 0
transform 0 -1 198 1 0 231
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2308
timestamp 0
transform 0 -1 198 1 0 230
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2307
timestamp 0
transform 0 -1 198 1 0 229
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2306
timestamp 0
transform 0 -1 198 1 0 228
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2305
timestamp 0
transform 0 -1 198 1 0 227
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2304
timestamp 0
transform 0 -1 198 1 0 226
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2303
timestamp 0
transform 0 -1 198 1 0 225
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2302
timestamp 0
transform 0 -1 198 1 0 224
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2301
timestamp 0
transform 0 -1 198 1 0 223
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2300
timestamp 0
transform 0 -1 198 1 0 222
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2299
timestamp 0
transform 0 -1 198 1 0 221
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2298
timestamp 0
transform 0 -1 198 1 0 220
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2297
timestamp 0
transform 0 -1 198 1 0 219
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2296
timestamp 0
transform 0 -1 198 1 0 218
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2295
timestamp 0
transform 0 -1 198 1 0 217
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2294
timestamp 0
transform 0 -1 198 1 0 216
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2293
timestamp 0
transform 0 -1 198 1 0 215
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2292
timestamp 0
transform 0 -1 198 1 0 214
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2291
timestamp 0
transform 0 -1 198 1 0 213
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2290
timestamp 0
transform 0 -1 198 1 0 212
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2289
timestamp 0
transform 0 -1 198 1 0 211
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2288
timestamp 0
transform 0 -1 198 1 0 210
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2287
timestamp 0
transform 0 -1 198 1 0 209
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2286
timestamp 0
transform 0 -1 198 1 0 208
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2285
timestamp 0
transform 0 -1 198 1 0 207
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2284
timestamp 0
transform 0 -1 198 1 0 206
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2283
timestamp 0
transform 0 -1 198 1 0 205
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2282
timestamp 0
transform 0 -1 198 1 0 204
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3330
timestamp 0
transform 0 1 2544 -1 0 262
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3329
timestamp 0
transform 0 1 2544 -1 0 261
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3328
timestamp 0
transform 0 1 2544 -1 0 260
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3327
timestamp 0
transform 0 1 2544 -1 0 259
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3326
timestamp 0
transform 0 1 2544 -1 0 258
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3325
timestamp 0
transform 0 1 2544 -1 0 257
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3324
timestamp 0
transform 0 1 2544 -1 0 256
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3323
timestamp 0
transform 0 1 2544 -1 0 255
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3322
timestamp 0
transform 0 1 2544 -1 0 254
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3321
timestamp 0
transform 0 1 2544 -1 0 253
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3320
timestamp 0
transform 0 1 2544 -1 0 252
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3319
timestamp 0
transform 0 1 2544 -1 0 251
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3318
timestamp 0
transform 0 1 2544 -1 0 250
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3317
timestamp 0
transform 0 1 2544 -1 0 249
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3316
timestamp 0
transform 0 1 2544 -1 0 248
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3315
timestamp 0
transform 0 1 2544 -1 0 247
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3314
timestamp 0
transform 0 1 2544 -1 0 246
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3313
timestamp 0
transform 0 1 2544 -1 0 245
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3312
timestamp 0
transform 0 1 2544 -1 0 244
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3311
timestamp 0
transform 0 1 2544 -1 0 243
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3310
timestamp 0
transform 0 1 2544 -1 0 242
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3309
timestamp 0
transform 0 1 2544 -1 0 241
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3308
timestamp 0
transform 0 1 2544 -1 0 240
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3307
timestamp 0
transform 0 1 2544 -1 0 239
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3306
timestamp 0
transform 0 1 2544 -1 0 238
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3305
timestamp 0
transform 0 1 2544 -1 0 237
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3304
timestamp 0
transform 0 1 2544 -1 0 236
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3303
timestamp 0
transform 0 1 2544 -1 0 235
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3302
timestamp 0
transform 0 1 2544 -1 0 234
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3301
timestamp 0
transform 0 1 2544 -1 0 233
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3300
timestamp 0
transform 0 1 2544 -1 0 232
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3299
timestamp 0
transform 0 1 2544 -1 0 231
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3298
timestamp 0
transform 0 1 2544 -1 0 230
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3297
timestamp 0
transform 0 1 2544 -1 0 229
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3296
timestamp 0
transform 0 1 2544 -1 0 228
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3295
timestamp 0
transform 0 1 2544 -1 0 227
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3294
timestamp 0
transform 0 1 2544 -1 0 226
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3293
timestamp 0
transform 0 1 2544 -1 0 225
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3292
timestamp 0
transform 0 1 2544 -1 0 224
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3291
timestamp 0
transform 0 1 2544 -1 0 223
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3290
timestamp 0
transform 0 1 2544 -1 0 222
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3289
timestamp 0
transform 0 1 2544 -1 0 221
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3288
timestamp 0
transform 0 1 2544 -1 0 220
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3287
timestamp 0
transform 0 1 2544 -1 0 219
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3286
timestamp 0
transform 0 1 2544 -1 0 218
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3285
timestamp 0
transform 0 1 2544 -1 0 217
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3284
timestamp 0
transform 0 1 2544 -1 0 216
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3283
timestamp 0
transform 0 1 2544 -1 0 215
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3282
timestamp 0
transform 0 1 2544 -1 0 214
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3281
timestamp 0
transform 0 1 2544 -1 0 213
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3280
timestamp 0
transform 0 1 2544 -1 0 212
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3279
timestamp 0
transform 0 1 2544 -1 0 211
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3278
timestamp 0
transform 0 1 2544 -1 0 210
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3277
timestamp 0
transform 0 1 2544 -1 0 209
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3276
timestamp 0
transform 0 1 2544 -1 0 208
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3275
timestamp 0
transform 0 1 2544 -1 0 207
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3274
timestamp 0
transform 0 1 2544 -1 0 206
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3273
timestamp 0
transform 0 1 2544 -1 0 205
box 0 0 1 1
use s8iom0_corner_pad  corner[1]
timestamp 0
transform -1 0 200 0 -1 204
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3272
timestamp 0
transform 0 1 2544 -1 0 204
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3271
timestamp 0
transform 0 1 2544 -1 0 203
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3270
timestamp 0
transform 0 1 2544 -1 0 202
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_3269
timestamp 0
transform 0 1 2544 -1 0 201
box 0 0 1 1
use s8iom0_corner_pad  corner[0]
timestamp 0
transform 0 1 2538 -1 0 200
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1025
timestamp 0
transform -1 0 201 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1026
timestamp 0
transform -1 0 202 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1027
timestamp 0
transform -1 0 203 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1028
timestamp 0
transform -1 0 204 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1029
timestamp 0
transform -1 0 205 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1030
timestamp 0
transform -1 0 206 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1031
timestamp 0
transform -1 0 207 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1032
timestamp 0
transform -1 0 208 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1033
timestamp 0
transform -1 0 209 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1034
timestamp 0
transform -1 0 210 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1035
timestamp 0
transform -1 0 211 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1036
timestamp 0
transform -1 0 212 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1037
timestamp 0
transform -1 0 213 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1038
timestamp 0
transform -1 0 214 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1039
timestamp 0
transform -1 0 215 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1040
timestamp 0
transform -1 0 216 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1041
timestamp 0
transform -1 0 217 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1042
timestamp 0
transform -1 0 218 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1043
timestamp 0
transform -1 0 219 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1044
timestamp 0
transform -1 0 220 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1045
timestamp 0
transform -1 0 221 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1046
timestamp 0
transform -1 0 222 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1047
timestamp 0
transform -1 0 223 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1048
timestamp 0
transform -1 0 224 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1049
timestamp 0
transform -1 0 225 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1050
timestamp 0
transform -1 0 226 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1051
timestamp 0
transform -1 0 227 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1052
timestamp 0
transform -1 0 228 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1053
timestamp 0
transform -1 0 229 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1054
timestamp 0
transform -1 0 230 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1055
timestamp 0
transform -1 0 231 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1056
timestamp 0
transform -1 0 232 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1057
timestamp 0
transform -1 0 233 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1058
timestamp 0
transform -1 0 234 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1059
timestamp 0
transform -1 0 235 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1060
timestamp 0
transform -1 0 236 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1061
timestamp 0
transform -1 0 237 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1062
timestamp 0
transform -1 0 238 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1063
timestamp 0
transform -1 0 239 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1064
timestamp 0
transform -1 0 240 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1065
timestamp 0
transform -1 0 241 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1066
timestamp 0
transform -1 0 242 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1067
timestamp 0
transform -1 0 243 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1068
timestamp 0
transform -1 0 244 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1069
timestamp 0
transform -1 0 245 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1070
timestamp 0
transform -1 0 246 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1071
timestamp 0
transform -1 0 247 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1072
timestamp 0
transform -1 0 248 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1073
timestamp 0
transform -1 0 249 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1074
timestamp 0
transform -1 0 250 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1075
timestamp 0
transform -1 0 251 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1076
timestamp 0
transform -1 0 252 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1077
timestamp 0
transform -1 0 253 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1078
timestamp 0
transform -1 0 254 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1079
timestamp 0
transform -1 0 255 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1080
timestamp 0
transform -1 0 256 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1081
timestamp 0
transform -1 0 257 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1082
timestamp 0
transform -1 0 258 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1083
timestamp 0
transform -1 0 259 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1084
timestamp 0
transform -1 0 260 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1085
timestamp 0
transform -1 0 261 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1086
timestamp 0
transform -1 0 262 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1087
timestamp 0
transform -1 0 263 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1088
timestamp 0
transform -1 0 264 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1089
timestamp 0
transform -1 0 265 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1090
timestamp 0
transform -1 0 266 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1091
timestamp 0
transform -1 0 267 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1092
timestamp 0
transform -1 0 268 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1093
timestamp 0
transform -1 0 269 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1094
timestamp 0
transform -1 0 270 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1095
timestamp 0
transform -1 0 271 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1096
timestamp 0
transform -1 0 272 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1097
timestamp 0
transform -1 0 273 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1098
timestamp 0
transform -1 0 274 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1099
timestamp 0
transform -1 0 275 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1100
timestamp 0
transform -1 0 276 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1101
timestamp 0
transform -1 0 277 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1102
timestamp 0
transform -1 0 278 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1103
timestamp 0
transform -1 0 279 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1104
timestamp 0
transform -1 0 280 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1105
timestamp 0
transform -1 0 281 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1106
timestamp 0
transform -1 0 282 0 -1 198
box 0 0 1 1
use s8iom0_vdda_hvc_pad  vddiohclamp[0]
timestamp 0
transform -1 0 357 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1108
timestamp 0
transform -1 0 358 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1109
timestamp 0
transform -1 0 359 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1110
timestamp 0
transform -1 0 360 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1111
timestamp 0
transform -1 0 361 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1112
timestamp 0
transform -1 0 362 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1113
timestamp 0
transform -1 0 363 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1114
timestamp 0
transform -1 0 364 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1115
timestamp 0
transform -1 0 365 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1116
timestamp 0
transform -1 0 366 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1117
timestamp 0
transform -1 0 367 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1118
timestamp 0
transform -1 0 368 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1119
timestamp 0
transform -1 0 369 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1120
timestamp 0
transform -1 0 370 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1121
timestamp 0
transform -1 0 371 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1122
timestamp 0
transform -1 0 372 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1123
timestamp 0
transform -1 0 373 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1124
timestamp 0
transform -1 0 374 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1125
timestamp 0
transform -1 0 375 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1126
timestamp 0
transform -1 0 376 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1127
timestamp 0
transform -1 0 377 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1128
timestamp 0
transform -1 0 378 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1129
timestamp 0
transform -1 0 379 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1130
timestamp 0
transform -1 0 380 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1131
timestamp 0
transform -1 0 381 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1132
timestamp 0
transform -1 0 382 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1133
timestamp 0
transform -1 0 383 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1134
timestamp 0
transform -1 0 384 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1135
timestamp 0
transform -1 0 385 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1136
timestamp 0
transform -1 0 386 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1137
timestamp 0
transform -1 0 387 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1138
timestamp 0
transform -1 0 388 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1139
timestamp 0
transform -1 0 389 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1140
timestamp 0
transform -1 0 390 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1141
timestamp 0
transform -1 0 391 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1142
timestamp 0
transform -1 0 392 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1143
timestamp 0
transform -1 0 393 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1144
timestamp 0
transform -1 0 394 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1145
timestamp 0
transform -1 0 395 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1146
timestamp 0
transform -1 0 396 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1147
timestamp 0
transform -1 0 397 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1148
timestamp 0
transform -1 0 398 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1149
timestamp 0
transform -1 0 399 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1150
timestamp 0
transform -1 0 400 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1151
timestamp 0
transform -1 0 401 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1152
timestamp 0
transform -1 0 402 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1153
timestamp 0
transform -1 0 403 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1154
timestamp 0
transform -1 0 404 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1155
timestamp 0
transform -1 0 405 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1156
timestamp 0
transform -1 0 406 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1157
timestamp 0
transform -1 0 407 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1158
timestamp 0
transform -1 0 408 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1159
timestamp 0
transform -1 0 409 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1160
timestamp 0
transform -1 0 410 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1161
timestamp 0
transform -1 0 411 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1162
timestamp 0
transform -1 0 412 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1163
timestamp 0
transform -1 0 413 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1164
timestamp 0
transform -1 0 414 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1165
timestamp 0
transform -1 0 415 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1166
timestamp 0
transform -1 0 416 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1167
timestamp 0
transform -1 0 417 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1168
timestamp 0
transform -1 0 418 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1169
timestamp 0
transform -1 0 419 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1170
timestamp 0
transform -1 0 420 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1171
timestamp 0
transform -1 0 421 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1172
timestamp 0
transform -1 0 422 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1173
timestamp 0
transform -1 0 423 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1174
timestamp 0
transform -1 0 424 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1175
timestamp 0
transform -1 0 425 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1176
timestamp 0
transform -1 0 426 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1177
timestamp 0
transform -1 0 427 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1178
timestamp 0
transform -1 0 428 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1179
timestamp 0
transform -1 0 429 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1180
timestamp 0
transform -1 0 430 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1181
timestamp 0
transform -1 0 431 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1182
timestamp 0
transform -1 0 432 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1183
timestamp 0
transform -1 0 433 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1184
timestamp 0
transform -1 0 434 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1185
timestamp 0
transform -1 0 435 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1186
timestamp 0
transform -1 0 436 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1187
timestamp 0
transform -1 0 437 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1188
timestamp 0
transform -1 0 438 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1189
timestamp 0
transform -1 0 439 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1190
timestamp 0
transform -1 0 440 0 -1 198
box 0 0 1 1
use s8iom0_vdda_lvc_pad  vdd3v3lclamp[2]
timestamp 0
transform -1 0 515 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1192
timestamp 0
transform -1 0 516 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1193
timestamp 0
transform -1 0 517 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1194
timestamp 0
transform -1 0 518 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1195
timestamp 0
transform -1 0 519 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1196
timestamp 0
transform -1 0 520 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1197
timestamp 0
transform -1 0 521 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1198
timestamp 0
transform -1 0 522 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1199
timestamp 0
transform -1 0 523 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1200
timestamp 0
transform -1 0 524 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1201
timestamp 0
transform -1 0 525 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1202
timestamp 0
transform -1 0 526 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1203
timestamp 0
transform -1 0 527 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1204
timestamp 0
transform -1 0 528 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1205
timestamp 0
transform -1 0 529 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1206
timestamp 0
transform -1 0 530 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1207
timestamp 0
transform -1 0 531 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1208
timestamp 0
transform -1 0 532 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1209
timestamp 0
transform -1 0 533 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1210
timestamp 0
transform -1 0 534 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1211
timestamp 0
transform -1 0 535 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1212
timestamp 0
transform -1 0 536 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1213
timestamp 0
transform -1 0 537 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1214
timestamp 0
transform -1 0 538 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1215
timestamp 0
transform -1 0 539 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1216
timestamp 0
transform -1 0 540 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1217
timestamp 0
transform -1 0 541 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1218
timestamp 0
transform -1 0 542 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1219
timestamp 0
transform -1 0 543 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1220
timestamp 0
transform -1 0 544 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1221
timestamp 0
transform -1 0 545 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1222
timestamp 0
transform -1 0 546 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1223
timestamp 0
transform -1 0 547 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1224
timestamp 0
transform -1 0 548 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1225
timestamp 0
transform -1 0 549 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1226
timestamp 0
transform -1 0 550 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1227
timestamp 0
transform -1 0 551 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1228
timestamp 0
transform -1 0 552 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1229
timestamp 0
transform -1 0 553 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1230
timestamp 0
transform -1 0 554 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1231
timestamp 0
transform -1 0 555 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1232
timestamp 0
transform -1 0 556 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1233
timestamp 0
transform -1 0 557 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1234
timestamp 0
transform -1 0 558 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1235
timestamp 0
transform -1 0 559 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1236
timestamp 0
transform -1 0 560 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1237
timestamp 0
transform -1 0 561 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1238
timestamp 0
transform -1 0 562 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1239
timestamp 0
transform -1 0 563 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1240
timestamp 0
transform -1 0 564 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1241
timestamp 0
transform -1 0 565 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1242
timestamp 0
transform -1 0 566 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1243
timestamp 0
transform -1 0 567 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1244
timestamp 0
transform -1 0 568 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1245
timestamp 0
transform -1 0 569 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1246
timestamp 0
transform -1 0 570 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1247
timestamp 0
transform -1 0 571 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1248
timestamp 0
transform -1 0 572 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1249
timestamp 0
transform -1 0 573 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1250
timestamp 0
transform -1 0 574 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1251
timestamp 0
transform -1 0 575 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1252
timestamp 0
transform -1 0 576 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1253
timestamp 0
transform -1 0 577 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1254
timestamp 0
transform -1 0 578 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1255
timestamp 0
transform -1 0 579 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1256
timestamp 0
transform -1 0 580 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1257
timestamp 0
transform -1 0 581 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1258
timestamp 0
transform -1 0 582 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1259
timestamp 0
transform -1 0 583 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1260
timestamp 0
transform -1 0 584 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1261
timestamp 0
transform -1 0 585 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1262
timestamp 0
transform -1 0 586 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1263
timestamp 0
transform -1 0 587 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1264
timestamp 0
transform -1 0 588 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1265
timestamp 0
transform -1 0 589 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1266
timestamp 0
transform -1 0 590 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1267
timestamp 0
transform -1 0 591 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1268
timestamp 0
transform -1 0 592 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1269
timestamp 0
transform -1 0 593 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1270
timestamp 0
transform -1 0 594 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1271
timestamp 0
transform -1 0 595 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1272
timestamp 0
transform -1 0 596 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1273
timestamp 0
transform -1 0 597 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1274
timestamp 0
transform -1 0 598 0 -1 198
box 0 0 1 1
use s8iom0_vccd_lvc_pad  vdd1v8lclamp[0]
timestamp 0
transform -1 0 673 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1276
timestamp 0
transform -1 0 674 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1277
timestamp 0
transform -1 0 675 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1278
timestamp 0
transform -1 0 676 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1279
timestamp 0
transform -1 0 677 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1280
timestamp 0
transform -1 0 678 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1281
timestamp 0
transform -1 0 679 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1282
timestamp 0
transform -1 0 680 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1283
timestamp 0
transform -1 0 681 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1284
timestamp 0
transform -1 0 682 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1285
timestamp 0
transform -1 0 683 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1286
timestamp 0
transform -1 0 684 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1287
timestamp 0
transform -1 0 685 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1288
timestamp 0
transform -1 0 686 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1289
timestamp 0
transform -1 0 687 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1290
timestamp 0
transform -1 0 688 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1291
timestamp 0
transform -1 0 689 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1292
timestamp 0
transform -1 0 690 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1293
timestamp 0
transform -1 0 691 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1294
timestamp 0
transform -1 0 692 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1295
timestamp 0
transform -1 0 693 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1296
timestamp 0
transform -1 0 694 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1297
timestamp 0
transform -1 0 695 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1298
timestamp 0
transform -1 0 696 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1299
timestamp 0
transform -1 0 697 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1300
timestamp 0
transform -1 0 698 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1301
timestamp 0
transform -1 0 699 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1302
timestamp 0
transform -1 0 700 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1303
timestamp 0
transform -1 0 701 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1304
timestamp 0
transform -1 0 702 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1305
timestamp 0
transform -1 0 703 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1306
timestamp 0
transform -1 0 704 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1307
timestamp 0
transform -1 0 705 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1308
timestamp 0
transform -1 0 706 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1309
timestamp 0
transform -1 0 707 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1310
timestamp 0
transform -1 0 708 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1311
timestamp 0
transform -1 0 709 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1312
timestamp 0
transform -1 0 710 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1313
timestamp 0
transform -1 0 711 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1314
timestamp 0
transform -1 0 712 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1315
timestamp 0
transform -1 0 713 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1316
timestamp 0
transform -1 0 714 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1317
timestamp 0
transform -1 0 715 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1318
timestamp 0
transform -1 0 716 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1319
timestamp 0
transform -1 0 717 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1320
timestamp 0
transform -1 0 718 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1321
timestamp 0
transform -1 0 719 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1322
timestamp 0
transform -1 0 720 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1323
timestamp 0
transform -1 0 721 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1324
timestamp 0
transform -1 0 722 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1325
timestamp 0
transform -1 0 723 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1326
timestamp 0
transform -1 0 724 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1327
timestamp 0
transform -1 0 725 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1328
timestamp 0
transform -1 0 726 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1329
timestamp 0
transform -1 0 727 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1330
timestamp 0
transform -1 0 728 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1331
timestamp 0
transform -1 0 729 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1332
timestamp 0
transform -1 0 730 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1333
timestamp 0
transform -1 0 731 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1334
timestamp 0
transform -1 0 732 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1335
timestamp 0
transform -1 0 733 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1336
timestamp 0
transform -1 0 734 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1337
timestamp 0
transform -1 0 735 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1338
timestamp 0
transform -1 0 736 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1339
timestamp 0
transform -1 0 737 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1340
timestamp 0
transform -1 0 738 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1341
timestamp 0
transform -1 0 739 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1342
timestamp 0
transform -1 0 740 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1343
timestamp 0
transform -1 0 741 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1344
timestamp 0
transform -1 0 742 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1345
timestamp 0
transform -1 0 743 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1346
timestamp 0
transform -1 0 744 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1347
timestamp 0
transform -1 0 745 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1348
timestamp 0
transform -1 0 746 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1349
timestamp 0
transform -1 0 747 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1350
timestamp 0
transform -1 0 748 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1351
timestamp 0
transform -1 0 749 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1352
timestamp 0
transform -1 0 750 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1353
timestamp 0
transform -1 0 751 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1354
timestamp 0
transform -1 0 752 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1355
timestamp 0
transform -1 0 753 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1356
timestamp 0
transform -1 0 754 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1357
timestamp 0
transform -1 0 755 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1358
timestamp 0
transform -1 0 756 0 -1 198
box 0 0 1 1
use s8iom0_vssa_hvc_pad  vsshclamp[1]
timestamp 0
transform -1 0 831 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1360
timestamp 0
transform -1 0 832 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1361
timestamp 0
transform -1 0 833 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1362
timestamp 0
transform -1 0 834 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1363
timestamp 0
transform -1 0 835 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1364
timestamp 0
transform -1 0 836 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1365
timestamp 0
transform -1 0 837 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1366
timestamp 0
transform -1 0 838 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1367
timestamp 0
transform -1 0 839 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1368
timestamp 0
transform -1 0 840 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1369
timestamp 0
transform -1 0 841 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1370
timestamp 0
transform -1 0 842 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1371
timestamp 0
transform -1 0 843 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1372
timestamp 0
transform -1 0 844 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1373
timestamp 0
transform -1 0 845 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1374
timestamp 0
transform -1 0 846 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1375
timestamp 0
transform -1 0 847 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1376
timestamp 0
transform -1 0 848 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1377
timestamp 0
transform -1 0 849 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1378
timestamp 0
transform -1 0 850 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1379
timestamp 0
transform -1 0 851 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1380
timestamp 0
transform -1 0 852 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1381
timestamp 0
transform -1 0 853 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1382
timestamp 0
transform -1 0 854 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1383
timestamp 0
transform -1 0 855 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1384
timestamp 0
transform -1 0 856 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1385
timestamp 0
transform -1 0 857 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1386
timestamp 0
transform -1 0 858 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1387
timestamp 0
transform -1 0 859 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1388
timestamp 0
transform -1 0 860 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1389
timestamp 0
transform -1 0 861 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1390
timestamp 0
transform -1 0 862 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1391
timestamp 0
transform -1 0 863 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1392
timestamp 0
transform -1 0 864 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1393
timestamp 0
transform -1 0 865 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1394
timestamp 0
transform -1 0 866 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1395
timestamp 0
transform -1 0 867 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1396
timestamp 0
transform -1 0 868 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1397
timestamp 0
transform -1 0 869 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1398
timestamp 0
transform -1 0 870 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1399
timestamp 0
transform -1 0 871 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1400
timestamp 0
transform -1 0 872 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1401
timestamp 0
transform -1 0 873 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1402
timestamp 0
transform -1 0 874 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1403
timestamp 0
transform -1 0 875 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1404
timestamp 0
transform -1 0 876 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1405
timestamp 0
transform -1 0 877 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1406
timestamp 0
transform -1 0 878 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1407
timestamp 0
transform -1 0 879 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1408
timestamp 0
transform -1 0 880 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1409
timestamp 0
transform -1 0 881 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1410
timestamp 0
transform -1 0 882 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1411
timestamp 0
transform -1 0 883 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1412
timestamp 0
transform -1 0 884 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1413
timestamp 0
transform -1 0 885 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1414
timestamp 0
transform -1 0 886 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1415
timestamp 0
transform -1 0 887 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1416
timestamp 0
transform -1 0 888 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1417
timestamp 0
transform -1 0 889 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1418
timestamp 0
transform -1 0 890 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1419
timestamp 0
transform -1 0 891 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1420
timestamp 0
transform -1 0 892 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1421
timestamp 0
transform -1 0 893 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1422
timestamp 0
transform -1 0 894 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1423
timestamp 0
transform -1 0 895 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1424
timestamp 0
transform -1 0 896 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1425
timestamp 0
transform -1 0 897 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1426
timestamp 0
transform -1 0 898 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1427
timestamp 0
transform -1 0 899 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1428
timestamp 0
transform -1 0 900 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1429
timestamp 0
transform -1 0 901 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1430
timestamp 0
transform -1 0 902 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1431
timestamp 0
transform -1 0 903 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1432
timestamp 0
transform -1 0 904 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1433
timestamp 0
transform -1 0 905 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1434
timestamp 0
transform -1 0 906 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1435
timestamp 0
transform -1 0 907 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1436
timestamp 0
transform -1 0 908 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1437
timestamp 0
transform -1 0 909 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1438
timestamp 0
transform -1 0 910 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1439
timestamp 0
transform -1 0 911 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1440
timestamp 0
transform -1 0 912 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1441
timestamp 0
transform -1 0 913 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1442
timestamp 0
transform -1 0 914 0 -1 198
box 0 0 1 1
use s8iom0_vssio_lvc_pad  vssiolclamp
timestamp 0
transform -1 0 989 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1444
timestamp 0
transform -1 0 990 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1445
timestamp 0
transform -1 0 991 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1446
timestamp 0
transform -1 0 992 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1447
timestamp 0
transform -1 0 993 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1448
timestamp 0
transform -1 0 994 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1449
timestamp 0
transform -1 0 995 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1450
timestamp 0
transform -1 0 996 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1451
timestamp 0
transform -1 0 997 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1452
timestamp 0
transform -1 0 998 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1453
timestamp 0
transform -1 0 999 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1454
timestamp 0
transform -1 0 1000 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1455
timestamp 0
transform -1 0 1001 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1456
timestamp 0
transform -1 0 1002 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1457
timestamp 0
transform -1 0 1003 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1458
timestamp 0
transform -1 0 1004 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1459
timestamp 0
transform -1 0 1005 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1460
timestamp 0
transform -1 0 1006 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1461
timestamp 0
transform -1 0 1007 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1462
timestamp 0
transform -1 0 1008 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1463
timestamp 0
transform -1 0 1009 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1464
timestamp 0
transform -1 0 1010 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1465
timestamp 0
transform -1 0 1011 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1466
timestamp 0
transform -1 0 1012 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1467
timestamp 0
transform -1 0 1013 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1468
timestamp 0
transform -1 0 1014 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1469
timestamp 0
transform -1 0 1015 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1470
timestamp 0
transform -1 0 1016 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1471
timestamp 0
transform -1 0 1017 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1472
timestamp 0
transform -1 0 1018 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1473
timestamp 0
transform -1 0 1019 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1474
timestamp 0
transform -1 0 1020 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1475
timestamp 0
transform -1 0 1021 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1476
timestamp 0
transform -1 0 1022 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1477
timestamp 0
transform -1 0 1023 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1478
timestamp 0
transform -1 0 1024 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1479
timestamp 0
transform -1 0 1025 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1480
timestamp 0
transform -1 0 1026 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1481
timestamp 0
transform -1 0 1027 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1482
timestamp 0
transform -1 0 1028 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1483
timestamp 0
transform -1 0 1029 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1484
timestamp 0
transform -1 0 1030 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1485
timestamp 0
transform -1 0 1031 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1486
timestamp 0
transform -1 0 1032 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1487
timestamp 0
transform -1 0 1033 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1488
timestamp 0
transform -1 0 1034 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1489
timestamp 0
transform -1 0 1035 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1490
timestamp 0
transform -1 0 1036 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1491
timestamp 0
transform -1 0 1037 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1492
timestamp 0
transform -1 0 1038 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1493
timestamp 0
transform -1 0 1039 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1494
timestamp 0
transform -1 0 1040 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1495
timestamp 0
transform -1 0 1041 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1496
timestamp 0
transform -1 0 1042 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1497
timestamp 0
transform -1 0 1043 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1498
timestamp 0
transform -1 0 1044 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1499
timestamp 0
transform -1 0 1045 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1500
timestamp 0
transform -1 0 1046 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1501
timestamp 0
transform -1 0 1047 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1502
timestamp 0
transform -1 0 1048 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1503
timestamp 0
transform -1 0 1049 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1504
timestamp 0
transform -1 0 1050 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1505
timestamp 0
transform -1 0 1051 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1506
timestamp 0
transform -1 0 1052 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1507
timestamp 0
transform -1 0 1053 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1508
timestamp 0
transform -1 0 1054 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1509
timestamp 0
transform -1 0 1055 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1510
timestamp 0
transform -1 0 1056 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1511
timestamp 0
transform -1 0 1057 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1512
timestamp 0
transform -1 0 1058 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1513
timestamp 0
transform -1 0 1059 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1514
timestamp 0
transform -1 0 1060 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1515
timestamp 0
transform -1 0 1061 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1516
timestamp 0
transform -1 0 1062 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1517
timestamp 0
transform -1 0 1063 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1518
timestamp 0
transform -1 0 1064 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1519
timestamp 0
transform -1 0 1065 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1520
timestamp 0
transform -1 0 1066 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1521
timestamp 0
transform -1 0 1067 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1522
timestamp 0
transform -1 0 1068 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1523
timestamp 0
transform -1 0 1069 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1524
timestamp 0
transform -1 0 1070 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1525
timestamp 0
transform -1 0 1071 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1526
timestamp 0
transform -1 0 1072 0 -1 198
box 0 0 1 1
use s8iom0_gpiov2_pad  comp_inn_pad
timestamp 0
transform -1 0 1152 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1528
timestamp 0
transform -1 0 1153 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1529
timestamp 0
transform -1 0 1154 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1530
timestamp 0
transform -1 0 1155 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1531
timestamp 0
transform -1 0 1156 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1532
timestamp 0
transform -1 0 1157 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1533
timestamp 0
transform -1 0 1158 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1534
timestamp 0
transform -1 0 1159 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1535
timestamp 0
transform -1 0 1160 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1536
timestamp 0
transform -1 0 1161 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1537
timestamp 0
transform -1 0 1162 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1538
timestamp 0
transform -1 0 1163 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1539
timestamp 0
transform -1 0 1164 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1540
timestamp 0
transform -1 0 1165 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1541
timestamp 0
transform -1 0 1166 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1542
timestamp 0
transform -1 0 1167 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1543
timestamp 0
transform -1 0 1168 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1544
timestamp 0
transform -1 0 1169 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1545
timestamp 0
transform -1 0 1170 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1546
timestamp 0
transform -1 0 1171 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1547
timestamp 0
transform -1 0 1172 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1548
timestamp 0
transform -1 0 1173 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1549
timestamp 0
transform -1 0 1174 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1550
timestamp 0
transform -1 0 1175 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1551
timestamp 0
transform -1 0 1176 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1552
timestamp 0
transform -1 0 1177 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1553
timestamp 0
transform -1 0 1178 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1554
timestamp 0
transform -1 0 1179 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1555
timestamp 0
transform -1 0 1180 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1556
timestamp 0
transform -1 0 1181 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1557
timestamp 0
transform -1 0 1182 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1558
timestamp 0
transform -1 0 1183 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1559
timestamp 0
transform -1 0 1184 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1560
timestamp 0
transform -1 0 1185 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1561
timestamp 0
transform -1 0 1186 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1562
timestamp 0
transform -1 0 1187 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1563
timestamp 0
transform -1 0 1188 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1564
timestamp 0
transform -1 0 1189 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1565
timestamp 0
transform -1 0 1190 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1566
timestamp 0
transform -1 0 1191 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1567
timestamp 0
transform -1 0 1192 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1568
timestamp 0
transform -1 0 1193 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1569
timestamp 0
transform -1 0 1194 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1570
timestamp 0
transform -1 0 1195 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1571
timestamp 0
transform -1 0 1196 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1572
timestamp 0
transform -1 0 1197 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1573
timestamp 0
transform -1 0 1198 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1574
timestamp 0
transform -1 0 1199 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1575
timestamp 0
transform -1 0 1200 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1576
timestamp 0
transform -1 0 1201 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1577
timestamp 0
transform -1 0 1202 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1578
timestamp 0
transform -1 0 1203 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1579
timestamp 0
transform -1 0 1204 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1580
timestamp 0
transform -1 0 1205 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1581
timestamp 0
transform -1 0 1206 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1582
timestamp 0
transform -1 0 1207 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1583
timestamp 0
transform -1 0 1208 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1584
timestamp 0
transform -1 0 1209 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1585
timestamp 0
transform -1 0 1210 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1586
timestamp 0
transform -1 0 1211 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1587
timestamp 0
transform -1 0 1212 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1588
timestamp 0
transform -1 0 1213 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1589
timestamp 0
transform -1 0 1214 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1590
timestamp 0
transform -1 0 1215 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1591
timestamp 0
transform -1 0 1216 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1592
timestamp 0
transform -1 0 1217 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1593
timestamp 0
transform -1 0 1218 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1594
timestamp 0
transform -1 0 1219 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1595
timestamp 0
transform -1 0 1220 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1596
timestamp 0
transform -1 0 1221 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1597
timestamp 0
transform -1 0 1222 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1598
timestamp 0
transform -1 0 1223 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1599
timestamp 0
transform -1 0 1224 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1600
timestamp 0
transform -1 0 1225 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1601
timestamp 0
transform -1 0 1226 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1602
timestamp 0
transform -1 0 1227 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1603
timestamp 0
transform -1 0 1228 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1604
timestamp 0
transform -1 0 1229 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1605
timestamp 0
transform -1 0 1230 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1606
timestamp 0
transform -1 0 1231 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1607
timestamp 0
transform -1 0 1232 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1608
timestamp 0
transform -1 0 1233 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1609
timestamp 0
transform -1 0 1234 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1610
timestamp 0
transform -1 0 1235 0 -1 198
box 0 0 1 1
use s8iom0_gpiov2_pad  adc_low_pad
timestamp 0
transform -1 0 1315 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1612
timestamp 0
transform -1 0 1316 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1613
timestamp 0
transform -1 0 1317 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1614
timestamp 0
transform -1 0 1318 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1615
timestamp 0
transform -1 0 1319 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1616
timestamp 0
transform -1 0 1320 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1617
timestamp 0
transform -1 0 1321 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1618
timestamp 0
transform -1 0 1322 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1619
timestamp 0
transform -1 0 1323 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1620
timestamp 0
transform -1 0 1324 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1621
timestamp 0
transform -1 0 1325 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1622
timestamp 0
transform -1 0 1326 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1623
timestamp 0
transform -1 0 1327 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1624
timestamp 0
transform -1 0 1328 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1625
timestamp 0
transform -1 0 1329 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1626
timestamp 0
transform -1 0 1330 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1627
timestamp 0
transform -1 0 1331 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1628
timestamp 0
transform -1 0 1332 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1629
timestamp 0
transform -1 0 1333 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1630
timestamp 0
transform -1 0 1334 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1631
timestamp 0
transform -1 0 1335 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1632
timestamp 0
transform -1 0 1336 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1633
timestamp 0
transform -1 0 1337 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1634
timestamp 0
transform -1 0 1338 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1635
timestamp 0
transform -1 0 1339 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1636
timestamp 0
transform -1 0 1340 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1637
timestamp 0
transform -1 0 1341 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1638
timestamp 0
transform -1 0 1342 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1639
timestamp 0
transform -1 0 1343 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1640
timestamp 0
transform -1 0 1344 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1641
timestamp 0
transform -1 0 1345 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1642
timestamp 0
transform -1 0 1346 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1643
timestamp 0
transform -1 0 1347 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1644
timestamp 0
transform -1 0 1348 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1645
timestamp 0
transform -1 0 1349 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1646
timestamp 0
transform -1 0 1350 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1647
timestamp 0
transform -1 0 1351 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1648
timestamp 0
transform -1 0 1352 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1649
timestamp 0
transform -1 0 1353 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1650
timestamp 0
transform -1 0 1354 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1651
timestamp 0
transform -1 0 1355 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1652
timestamp 0
transform -1 0 1356 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1653
timestamp 0
transform -1 0 1357 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1654
timestamp 0
transform -1 0 1358 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1655
timestamp 0
transform -1 0 1359 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1656
timestamp 0
transform -1 0 1360 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1657
timestamp 0
transform -1 0 1361 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1658
timestamp 0
transform -1 0 1362 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1659
timestamp 0
transform -1 0 1363 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1660
timestamp 0
transform -1 0 1364 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1661
timestamp 0
transform -1 0 1365 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1662
timestamp 0
transform -1 0 1366 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1663
timestamp 0
transform -1 0 1367 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1664
timestamp 0
transform -1 0 1368 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1665
timestamp 0
transform -1 0 1369 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1666
timestamp 0
transform -1 0 1370 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1667
timestamp 0
transform -1 0 1371 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1668
timestamp 0
transform -1 0 1372 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1669
timestamp 0
transform -1 0 1373 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1670
timestamp 0
transform -1 0 1374 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1671
timestamp 0
transform -1 0 1375 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1672
timestamp 0
transform -1 0 1376 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1673
timestamp 0
transform -1 0 1377 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1674
timestamp 0
transform -1 0 1378 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1675
timestamp 0
transform -1 0 1379 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1676
timestamp 0
transform -1 0 1380 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1677
timestamp 0
transform -1 0 1381 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1678
timestamp 0
transform -1 0 1382 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1679
timestamp 0
transform -1 0 1383 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1680
timestamp 0
transform -1 0 1384 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1681
timestamp 0
transform -1 0 1385 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1682
timestamp 0
transform -1 0 1386 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1683
timestamp 0
transform -1 0 1387 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1684
timestamp 0
transform -1 0 1388 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1685
timestamp 0
transform -1 0 1389 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1686
timestamp 0
transform -1 0 1390 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1687
timestamp 0
transform -1 0 1391 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1688
timestamp 0
transform -1 0 1392 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1689
timestamp 0
transform -1 0 1393 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1690
timestamp 0
transform -1 0 1394 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1691
timestamp 0
transform -1 0 1395 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1692
timestamp 0
transform -1 0 1396 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1693
timestamp 0
transform -1 0 1397 0 -1 198
box 0 0 1 1
use s8iom0_gpiov2_pad  adc_high_pad
timestamp 0
transform -1 0 1477 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1695
timestamp 0
transform -1 0 1478 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1696
timestamp 0
transform -1 0 1479 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1697
timestamp 0
transform -1 0 1480 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1698
timestamp 0
transform -1 0 1481 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1699
timestamp 0
transform -1 0 1482 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1700
timestamp 0
transform -1 0 1483 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1701
timestamp 0
transform -1 0 1484 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1702
timestamp 0
transform -1 0 1485 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1703
timestamp 0
transform -1 0 1486 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1704
timestamp 0
transform -1 0 1487 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1705
timestamp 0
transform -1 0 1488 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1706
timestamp 0
transform -1 0 1489 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1707
timestamp 0
transform -1 0 1490 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1708
timestamp 0
transform -1 0 1491 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1709
timestamp 0
transform -1 0 1492 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1710
timestamp 0
transform -1 0 1493 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1711
timestamp 0
transform -1 0 1494 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1712
timestamp 0
transform -1 0 1495 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1713
timestamp 0
transform -1 0 1496 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1714
timestamp 0
transform -1 0 1497 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1715
timestamp 0
transform -1 0 1498 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1716
timestamp 0
transform -1 0 1499 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1717
timestamp 0
transform -1 0 1500 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1718
timestamp 0
transform -1 0 1501 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1719
timestamp 0
transform -1 0 1502 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1720
timestamp 0
transform -1 0 1503 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1721
timestamp 0
transform -1 0 1504 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1722
timestamp 0
transform -1 0 1505 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1723
timestamp 0
transform -1 0 1506 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1724
timestamp 0
transform -1 0 1507 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1725
timestamp 0
transform -1 0 1508 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1726
timestamp 0
transform -1 0 1509 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1727
timestamp 0
transform -1 0 1510 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1728
timestamp 0
transform -1 0 1511 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1729
timestamp 0
transform -1 0 1512 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1730
timestamp 0
transform -1 0 1513 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1731
timestamp 0
transform -1 0 1514 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1732
timestamp 0
transform -1 0 1515 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1733
timestamp 0
transform -1 0 1516 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1734
timestamp 0
transform -1 0 1517 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1735
timestamp 0
transform -1 0 1518 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1736
timestamp 0
transform -1 0 1519 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1737
timestamp 0
transform -1 0 1520 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1738
timestamp 0
transform -1 0 1521 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1739
timestamp 0
transform -1 0 1522 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1740
timestamp 0
transform -1 0 1523 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1741
timestamp 0
transform -1 0 1524 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1742
timestamp 0
transform -1 0 1525 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1743
timestamp 0
transform -1 0 1526 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1744
timestamp 0
transform -1 0 1527 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1745
timestamp 0
transform -1 0 1528 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1746
timestamp 0
transform -1 0 1529 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1747
timestamp 0
transform -1 0 1530 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1748
timestamp 0
transform -1 0 1531 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1749
timestamp 0
transform -1 0 1532 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1750
timestamp 0
transform -1 0 1533 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1751
timestamp 0
transform -1 0 1534 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1752
timestamp 0
transform -1 0 1535 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1753
timestamp 0
transform -1 0 1536 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1754
timestamp 0
transform -1 0 1537 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1755
timestamp 0
transform -1 0 1538 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1756
timestamp 0
transform -1 0 1539 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1757
timestamp 0
transform -1 0 1540 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1758
timestamp 0
transform -1 0 1541 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1759
timestamp 0
transform -1 0 1542 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1760
timestamp 0
transform -1 0 1543 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1761
timestamp 0
transform -1 0 1544 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1762
timestamp 0
transform -1 0 1545 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1763
timestamp 0
transform -1 0 1546 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1764
timestamp 0
transform -1 0 1547 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1765
timestamp 0
transform -1 0 1548 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1766
timestamp 0
transform -1 0 1549 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1767
timestamp 0
transform -1 0 1550 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1768
timestamp 0
transform -1 0 1551 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1769
timestamp 0
transform -1 0 1552 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1770
timestamp 0
transform -1 0 1553 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1771
timestamp 0
transform -1 0 1554 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1772
timestamp 0
transform -1 0 1555 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1773
timestamp 0
transform -1 0 1556 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1774
timestamp 0
transform -1 0 1557 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1775
timestamp 0
transform -1 0 1558 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1776
timestamp 0
transform -1 0 1559 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1777
timestamp 0
transform -1 0 1560 0 -1 198
box 0 0 1 1
use s8iom0_gpiov2_pad  adc1_in_pad
timestamp 0
transform -1 0 1640 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1779
timestamp 0
transform -1 0 1641 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1780
timestamp 0
transform -1 0 1642 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1781
timestamp 0
transform -1 0 1643 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1782
timestamp 0
transform -1 0 1644 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1783
timestamp 0
transform -1 0 1645 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1784
timestamp 0
transform -1 0 1646 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1785
timestamp 0
transform -1 0 1647 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1786
timestamp 0
transform -1 0 1648 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1787
timestamp 0
transform -1 0 1649 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1788
timestamp 0
transform -1 0 1650 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1789
timestamp 0
transform -1 0 1651 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1790
timestamp 0
transform -1 0 1652 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1791
timestamp 0
transform -1 0 1653 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1792
timestamp 0
transform -1 0 1654 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1793
timestamp 0
transform -1 0 1655 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1794
timestamp 0
transform -1 0 1656 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1795
timestamp 0
transform -1 0 1657 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1796
timestamp 0
transform -1 0 1658 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1797
timestamp 0
transform -1 0 1659 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1798
timestamp 0
transform -1 0 1660 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1799
timestamp 0
transform -1 0 1661 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1800
timestamp 0
transform -1 0 1662 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1801
timestamp 0
transform -1 0 1663 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1802
timestamp 0
transform -1 0 1664 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1803
timestamp 0
transform -1 0 1665 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1804
timestamp 0
transform -1 0 1666 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1805
timestamp 0
transform -1 0 1667 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1806
timestamp 0
transform -1 0 1668 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1807
timestamp 0
transform -1 0 1669 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1808
timestamp 0
transform -1 0 1670 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1809
timestamp 0
transform -1 0 1671 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1810
timestamp 0
transform -1 0 1672 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1811
timestamp 0
transform -1 0 1673 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1812
timestamp 0
transform -1 0 1674 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1813
timestamp 0
transform -1 0 1675 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1814
timestamp 0
transform -1 0 1676 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1815
timestamp 0
transform -1 0 1677 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1816
timestamp 0
transform -1 0 1678 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1817
timestamp 0
transform -1 0 1679 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1818
timestamp 0
transform -1 0 1680 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1819
timestamp 0
transform -1 0 1681 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1820
timestamp 0
transform -1 0 1682 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1821
timestamp 0
transform -1 0 1683 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1822
timestamp 0
transform -1 0 1684 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1823
timestamp 0
transform -1 0 1685 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1824
timestamp 0
transform -1 0 1686 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1825
timestamp 0
transform -1 0 1687 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1826
timestamp 0
transform -1 0 1688 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1827
timestamp 0
transform -1 0 1689 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1828
timestamp 0
transform -1 0 1690 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1829
timestamp 0
transform -1 0 1691 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1830
timestamp 0
transform -1 0 1692 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1831
timestamp 0
transform -1 0 1693 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1832
timestamp 0
transform -1 0 1694 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1833
timestamp 0
transform -1 0 1695 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1834
timestamp 0
transform -1 0 1696 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1835
timestamp 0
transform -1 0 1697 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1836
timestamp 0
transform -1 0 1698 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1837
timestamp 0
transform -1 0 1699 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1838
timestamp 0
transform -1 0 1700 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1839
timestamp 0
transform -1 0 1701 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1840
timestamp 0
transform -1 0 1702 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1841
timestamp 0
transform -1 0 1703 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1842
timestamp 0
transform -1 0 1704 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1843
timestamp 0
transform -1 0 1705 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1844
timestamp 0
transform -1 0 1706 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1845
timestamp 0
transform -1 0 1707 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1846
timestamp 0
transform -1 0 1708 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1847
timestamp 0
transform -1 0 1709 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1848
timestamp 0
transform -1 0 1710 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1849
timestamp 0
transform -1 0 1711 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1850
timestamp 0
transform -1 0 1712 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1851
timestamp 0
transform -1 0 1713 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1852
timestamp 0
transform -1 0 1714 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1853
timestamp 0
transform -1 0 1715 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1854
timestamp 0
transform -1 0 1716 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1855
timestamp 0
transform -1 0 1717 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1856
timestamp 0
transform -1 0 1718 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1857
timestamp 0
transform -1 0 1719 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1858
timestamp 0
transform -1 0 1720 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1859
timestamp 0
transform -1 0 1721 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1860
timestamp 0
transform -1 0 1722 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1861
timestamp 0
transform -1 0 1723 0 -1 198
box 0 0 1 1
use s8iom0_gpiov2_pad  adc0_in_pad
timestamp 0
transform -1 0 1803 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1863
timestamp 0
transform -1 0 1804 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1864
timestamp 0
transform -1 0 1805 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1865
timestamp 0
transform -1 0 1806 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1866
timestamp 0
transform -1 0 1807 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1867
timestamp 0
transform -1 0 1808 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1868
timestamp 0
transform -1 0 1809 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1869
timestamp 0
transform -1 0 1810 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1870
timestamp 0
transform -1 0 1811 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1871
timestamp 0
transform -1 0 1812 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1872
timestamp 0
transform -1 0 1813 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1873
timestamp 0
transform -1 0 1814 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1874
timestamp 0
transform -1 0 1815 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1875
timestamp 0
transform -1 0 1816 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1876
timestamp 0
transform -1 0 1817 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1877
timestamp 0
transform -1 0 1818 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1878
timestamp 0
transform -1 0 1819 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1879
timestamp 0
transform -1 0 1820 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1880
timestamp 0
transform -1 0 1821 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1881
timestamp 0
transform -1 0 1822 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1882
timestamp 0
transform -1 0 1823 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1883
timestamp 0
transform -1 0 1824 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1884
timestamp 0
transform -1 0 1825 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1885
timestamp 0
transform -1 0 1826 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1886
timestamp 0
transform -1 0 1827 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1887
timestamp 0
transform -1 0 1828 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1888
timestamp 0
transform -1 0 1829 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1889
timestamp 0
transform -1 0 1830 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1890
timestamp 0
transform -1 0 1831 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1891
timestamp 0
transform -1 0 1832 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1892
timestamp 0
transform -1 0 1833 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1893
timestamp 0
transform -1 0 1834 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1894
timestamp 0
transform -1 0 1835 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1895
timestamp 0
transform -1 0 1836 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1896
timestamp 0
transform -1 0 1837 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1897
timestamp 0
transform -1 0 1838 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1898
timestamp 0
transform -1 0 1839 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1899
timestamp 0
transform -1 0 1840 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1900
timestamp 0
transform -1 0 1841 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1901
timestamp 0
transform -1 0 1842 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1902
timestamp 0
transform -1 0 1843 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1903
timestamp 0
transform -1 0 1844 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1904
timestamp 0
transform -1 0 1845 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1905
timestamp 0
transform -1 0 1846 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1906
timestamp 0
transform -1 0 1847 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1907
timestamp 0
transform -1 0 1848 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1908
timestamp 0
transform -1 0 1849 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1909
timestamp 0
transform -1 0 1850 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1910
timestamp 0
transform -1 0 1851 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1911
timestamp 0
transform -1 0 1852 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1912
timestamp 0
transform -1 0 1853 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1913
timestamp 0
transform -1 0 1854 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1914
timestamp 0
transform -1 0 1855 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1915
timestamp 0
transform -1 0 1856 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1916
timestamp 0
transform -1 0 1857 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1917
timestamp 0
transform -1 0 1858 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1918
timestamp 0
transform -1 0 1859 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1919
timestamp 0
transform -1 0 1860 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1920
timestamp 0
transform -1 0 1861 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1921
timestamp 0
transform -1 0 1862 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1922
timestamp 0
transform -1 0 1863 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1923
timestamp 0
transform -1 0 1864 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1924
timestamp 0
transform -1 0 1865 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1925
timestamp 0
transform -1 0 1866 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1926
timestamp 0
transform -1 0 1867 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1927
timestamp 0
transform -1 0 1868 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1928
timestamp 0
transform -1 0 1869 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1929
timestamp 0
transform -1 0 1870 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1930
timestamp 0
transform -1 0 1871 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1931
timestamp 0
transform -1 0 1872 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1932
timestamp 0
transform -1 0 1873 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1933
timestamp 0
transform -1 0 1874 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1934
timestamp 0
transform -1 0 1875 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1935
timestamp 0
transform -1 0 1876 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1936
timestamp 0
transform -1 0 1877 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1937
timestamp 0
transform -1 0 1878 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1938
timestamp 0
transform -1 0 1879 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1939
timestamp 0
transform -1 0 1880 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1940
timestamp 0
transform -1 0 1881 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1941
timestamp 0
transform -1 0 1882 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1942
timestamp 0
transform -1 0 1883 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1943
timestamp 0
transform -1 0 1884 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1944
timestamp 0
transform -1 0 1885 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1945
timestamp 0
transform -1 0 1886 0 -1 198
box 0 0 1 1
use s8iom0_gpiov2_pad  xo_pad
timestamp 0
transform -1 0 1966 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1947
timestamp 0
transform -1 0 1967 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1948
timestamp 0
transform -1 0 1968 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1949
timestamp 0
transform -1 0 1969 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1950
timestamp 0
transform -1 0 1970 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1951
timestamp 0
transform -1 0 1971 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1952
timestamp 0
transform -1 0 1972 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1953
timestamp 0
transform -1 0 1973 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1954
timestamp 0
transform -1 0 1974 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1955
timestamp 0
transform -1 0 1975 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1956
timestamp 0
transform -1 0 1976 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1957
timestamp 0
transform -1 0 1977 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1958
timestamp 0
transform -1 0 1978 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1959
timestamp 0
transform -1 0 1979 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1960
timestamp 0
transform -1 0 1980 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1961
timestamp 0
transform -1 0 1981 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1962
timestamp 0
transform -1 0 1982 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1963
timestamp 0
transform -1 0 1983 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1964
timestamp 0
transform -1 0 1984 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1965
timestamp 0
transform -1 0 1985 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1966
timestamp 0
transform -1 0 1986 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1967
timestamp 0
transform -1 0 1987 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1968
timestamp 0
transform -1 0 1988 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1969
timestamp 0
transform -1 0 1989 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1970
timestamp 0
transform -1 0 1990 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1971
timestamp 0
transform -1 0 1991 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1972
timestamp 0
transform -1 0 1992 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1973
timestamp 0
transform -1 0 1993 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1974
timestamp 0
transform -1 0 1994 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1975
timestamp 0
transform -1 0 1995 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1976
timestamp 0
transform -1 0 1996 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1977
timestamp 0
transform -1 0 1997 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1978
timestamp 0
transform -1 0 1998 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1979
timestamp 0
transform -1 0 1999 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1980
timestamp 0
transform -1 0 2000 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1981
timestamp 0
transform -1 0 2001 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1982
timestamp 0
transform -1 0 2002 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1983
timestamp 0
transform -1 0 2003 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1984
timestamp 0
transform -1 0 2004 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1985
timestamp 0
transform -1 0 2005 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1986
timestamp 0
transform -1 0 2006 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1987
timestamp 0
transform -1 0 2007 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1988
timestamp 0
transform -1 0 2008 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1989
timestamp 0
transform -1 0 2009 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1990
timestamp 0
transform -1 0 2010 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1991
timestamp 0
transform -1 0 2011 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1992
timestamp 0
transform -1 0 2012 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1993
timestamp 0
transform -1 0 2013 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1994
timestamp 0
transform -1 0 2014 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1995
timestamp 0
transform -1 0 2015 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1996
timestamp 0
transform -1 0 2016 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1997
timestamp 0
transform -1 0 2017 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1998
timestamp 0
transform -1 0 2018 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_1999
timestamp 0
transform -1 0 2019 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2000
timestamp 0
transform -1 0 2020 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2001
timestamp 0
transform -1 0 2021 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2002
timestamp 0
transform -1 0 2022 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2003
timestamp 0
transform -1 0 2023 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2004
timestamp 0
transform -1 0 2024 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2005
timestamp 0
transform -1 0 2025 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2006
timestamp 0
transform -1 0 2026 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2007
timestamp 0
transform -1 0 2027 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2008
timestamp 0
transform -1 0 2028 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2009
timestamp 0
transform -1 0 2029 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2010
timestamp 0
transform -1 0 2030 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2011
timestamp 0
transform -1 0 2031 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2012
timestamp 0
transform -1 0 2032 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2013
timestamp 0
transform -1 0 2033 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2014
timestamp 0
transform -1 0 2034 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2015
timestamp 0
transform -1 0 2035 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2016
timestamp 0
transform -1 0 2036 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2017
timestamp 0
transform -1 0 2037 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2018
timestamp 0
transform -1 0 2038 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2019
timestamp 0
transform -1 0 2039 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2020
timestamp 0
transform -1 0 2040 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2021
timestamp 0
transform -1 0 2041 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2022
timestamp 0
transform -1 0 2042 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2023
timestamp 0
transform -1 0 2043 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2024
timestamp 0
transform -1 0 2044 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2025
timestamp 0
transform -1 0 2045 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2026
timestamp 0
transform -1 0 2046 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2027
timestamp 0
transform -1 0 2047 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2028
timestamp 0
transform -1 0 2048 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2029
timestamp 0
transform -1 0 2049 0 -1 198
box 0 0 1 1
use s8iom0_gpiov2_pad  xi_pad
timestamp 0
transform -1 0 2129 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2031
timestamp 0
transform -1 0 2130 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2032
timestamp 0
transform -1 0 2131 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2033
timestamp 0
transform -1 0 2132 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2034
timestamp 0
transform -1 0 2133 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2035
timestamp 0
transform -1 0 2134 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2036
timestamp 0
transform -1 0 2135 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2037
timestamp 0
transform -1 0 2136 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2038
timestamp 0
transform -1 0 2137 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2039
timestamp 0
transform -1 0 2138 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2040
timestamp 0
transform -1 0 2139 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2041
timestamp 0
transform -1 0 2140 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2042
timestamp 0
transform -1 0 2141 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2043
timestamp 0
transform -1 0 2142 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2044
timestamp 0
transform -1 0 2143 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2045
timestamp 0
transform -1 0 2144 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2046
timestamp 0
transform -1 0 2145 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2047
timestamp 0
transform -1 0 2146 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2048
timestamp 0
transform -1 0 2147 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2049
timestamp 0
transform -1 0 2148 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2050
timestamp 0
transform -1 0 2149 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2051
timestamp 0
transform -1 0 2150 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2052
timestamp 0
transform -1 0 2151 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2053
timestamp 0
transform -1 0 2152 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2054
timestamp 0
transform -1 0 2153 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2055
timestamp 0
transform -1 0 2154 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2056
timestamp 0
transform -1 0 2155 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2057
timestamp 0
transform -1 0 2156 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2058
timestamp 0
transform -1 0 2157 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2059
timestamp 0
transform -1 0 2158 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2060
timestamp 0
transform -1 0 2159 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2061
timestamp 0
transform -1 0 2160 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2062
timestamp 0
transform -1 0 2161 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2063
timestamp 0
transform -1 0 2162 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2064
timestamp 0
transform -1 0 2163 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2065
timestamp 0
transform -1 0 2164 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2066
timestamp 0
transform -1 0 2165 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2067
timestamp 0
transform -1 0 2166 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2068
timestamp 0
transform -1 0 2167 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2069
timestamp 0
transform -1 0 2168 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2070
timestamp 0
transform -1 0 2169 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2071
timestamp 0
transform -1 0 2170 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2072
timestamp 0
transform -1 0 2171 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2073
timestamp 0
transform -1 0 2172 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2074
timestamp 0
transform -1 0 2173 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2075
timestamp 0
transform -1 0 2174 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2076
timestamp 0
transform -1 0 2175 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2077
timestamp 0
transform -1 0 2176 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2078
timestamp 0
transform -1 0 2177 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2079
timestamp 0
transform -1 0 2178 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2080
timestamp 0
transform -1 0 2179 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2081
timestamp 0
transform -1 0 2180 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2082
timestamp 0
transform -1 0 2181 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2083
timestamp 0
transform -1 0 2182 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2084
timestamp 0
transform -1 0 2183 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2085
timestamp 0
transform -1 0 2184 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2086
timestamp 0
transform -1 0 2185 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2087
timestamp 0
transform -1 0 2186 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2088
timestamp 0
transform -1 0 2187 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2089
timestamp 0
transform -1 0 2188 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2090
timestamp 0
transform -1 0 2189 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2091
timestamp 0
transform -1 0 2190 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2092
timestamp 0
transform -1 0 2191 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2093
timestamp 0
transform -1 0 2192 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2094
timestamp 0
transform -1 0 2193 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2095
timestamp 0
transform -1 0 2194 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2096
timestamp 0
transform -1 0 2195 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2097
timestamp 0
transform -1 0 2196 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2098
timestamp 0
transform -1 0 2197 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2099
timestamp 0
transform -1 0 2198 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2100
timestamp 0
transform -1 0 2199 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2101
timestamp 0
transform -1 0 2200 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2102
timestamp 0
transform -1 0 2201 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2103
timestamp 0
transform -1 0 2202 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2104
timestamp 0
transform -1 0 2203 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2105
timestamp 0
transform -1 0 2204 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2106
timestamp 0
transform -1 0 2205 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2107
timestamp 0
transform -1 0 2206 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2108
timestamp 0
transform -1 0 2207 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2109
timestamp 0
transform -1 0 2208 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2110
timestamp 0
transform -1 0 2209 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2111
timestamp 0
transform -1 0 2210 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2112
timestamp 0
transform -1 0 2211 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2113
timestamp 0
transform -1 0 2212 0 -1 198
box 0 0 1 1
use s8iom0_gpiov2_pad  gpio_pad[10]
timestamp 0
transform -1 0 2292 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2115
timestamp 0
transform -1 0 2293 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2116
timestamp 0
transform -1 0 2294 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2117
timestamp 0
transform -1 0 2295 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2118
timestamp 0
transform -1 0 2296 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2119
timestamp 0
transform -1 0 2297 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2120
timestamp 0
transform -1 0 2298 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2121
timestamp 0
transform -1 0 2299 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2122
timestamp 0
transform -1 0 2300 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2123
timestamp 0
transform -1 0 2301 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2124
timestamp 0
transform -1 0 2302 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2125
timestamp 0
transform -1 0 2303 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2126
timestamp 0
transform -1 0 2304 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2127
timestamp 0
transform -1 0 2305 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2128
timestamp 0
transform -1 0 2306 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2129
timestamp 0
transform -1 0 2307 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2130
timestamp 0
transform -1 0 2308 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2131
timestamp 0
transform -1 0 2309 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2132
timestamp 0
transform -1 0 2310 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2133
timestamp 0
transform -1 0 2311 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2134
timestamp 0
transform -1 0 2312 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2135
timestamp 0
transform -1 0 2313 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2136
timestamp 0
transform -1 0 2314 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2137
timestamp 0
transform -1 0 2315 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2138
timestamp 0
transform -1 0 2316 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2139
timestamp 0
transform -1 0 2317 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2140
timestamp 0
transform -1 0 2318 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2141
timestamp 0
transform -1 0 2319 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2142
timestamp 0
transform -1 0 2320 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2143
timestamp 0
transform -1 0 2321 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2144
timestamp 0
transform -1 0 2322 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2145
timestamp 0
transform -1 0 2323 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2146
timestamp 0
transform -1 0 2324 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2147
timestamp 0
transform -1 0 2325 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2148
timestamp 0
transform -1 0 2326 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2149
timestamp 0
transform -1 0 2327 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2150
timestamp 0
transform -1 0 2328 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2151
timestamp 0
transform -1 0 2329 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2152
timestamp 0
transform -1 0 2330 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2153
timestamp 0
transform -1 0 2331 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2154
timestamp 0
transform -1 0 2332 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2155
timestamp 0
transform -1 0 2333 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2156
timestamp 0
transform -1 0 2334 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2157
timestamp 0
transform -1 0 2335 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2158
timestamp 0
transform -1 0 2336 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2159
timestamp 0
transform -1 0 2337 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2160
timestamp 0
transform -1 0 2338 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2161
timestamp 0
transform -1 0 2339 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2162
timestamp 0
transform -1 0 2340 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2163
timestamp 0
transform -1 0 2341 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2164
timestamp 0
transform -1 0 2342 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2165
timestamp 0
transform -1 0 2343 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2166
timestamp 0
transform -1 0 2344 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2167
timestamp 0
transform -1 0 2345 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2168
timestamp 0
transform -1 0 2346 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2169
timestamp 0
transform -1 0 2347 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2170
timestamp 0
transform -1 0 2348 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2171
timestamp 0
transform -1 0 2349 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2172
timestamp 0
transform -1 0 2350 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2173
timestamp 0
transform -1 0 2351 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2174
timestamp 0
transform -1 0 2352 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2175
timestamp 0
transform -1 0 2353 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2176
timestamp 0
transform -1 0 2354 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2177
timestamp 0
transform -1 0 2355 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2178
timestamp 0
transform -1 0 2356 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2179
timestamp 0
transform -1 0 2357 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2180
timestamp 0
transform -1 0 2358 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2181
timestamp 0
transform -1 0 2359 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2182
timestamp 0
transform -1 0 2360 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2183
timestamp 0
transform -1 0 2361 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2184
timestamp 0
transform -1 0 2362 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2185
timestamp 0
transform -1 0 2363 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2186
timestamp 0
transform -1 0 2364 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2187
timestamp 0
transform -1 0 2365 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2188
timestamp 0
transform -1 0 2366 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2189
timestamp 0
transform -1 0 2367 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2190
timestamp 0
transform -1 0 2368 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2191
timestamp 0
transform -1 0 2369 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2192
timestamp 0
transform -1 0 2370 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2193
timestamp 0
transform -1 0 2371 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2194
timestamp 0
transform -1 0 2372 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2195
timestamp 0
transform -1 0 2373 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2196
timestamp 0
transform -1 0 2374 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2197
timestamp 0
transform -1 0 2375 0 -1 198
box 0 0 1 1
use s8iom0_gpiov2_pad  gpio_pad[9]
timestamp 0
transform -1 0 2455 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2199
timestamp 0
transform -1 0 2456 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2200
timestamp 0
transform -1 0 2457 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2201
timestamp 0
transform -1 0 2458 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2202
timestamp 0
transform -1 0 2459 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2203
timestamp 0
transform -1 0 2460 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2204
timestamp 0
transform -1 0 2461 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2205
timestamp 0
transform -1 0 2462 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2206
timestamp 0
transform -1 0 2463 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2207
timestamp 0
transform -1 0 2464 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2208
timestamp 0
transform -1 0 2465 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2209
timestamp 0
transform -1 0 2466 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2210
timestamp 0
transform -1 0 2467 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2211
timestamp 0
transform -1 0 2468 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2212
timestamp 0
transform -1 0 2469 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2213
timestamp 0
transform -1 0 2470 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2214
timestamp 0
transform -1 0 2471 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2215
timestamp 0
transform -1 0 2472 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2216
timestamp 0
transform -1 0 2473 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2217
timestamp 0
transform -1 0 2474 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2218
timestamp 0
transform -1 0 2475 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2219
timestamp 0
transform -1 0 2476 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2220
timestamp 0
transform -1 0 2477 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2221
timestamp 0
transform -1 0 2478 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2222
timestamp 0
transform -1 0 2479 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2223
timestamp 0
transform -1 0 2480 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2224
timestamp 0
transform -1 0 2481 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2225
timestamp 0
transform -1 0 2482 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2226
timestamp 0
transform -1 0 2483 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2227
timestamp 0
transform -1 0 2484 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2228
timestamp 0
transform -1 0 2485 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2229
timestamp 0
transform -1 0 2486 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2230
timestamp 0
transform -1 0 2487 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2231
timestamp 0
transform -1 0 2488 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2232
timestamp 0
transform -1 0 2489 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2233
timestamp 0
transform -1 0 2490 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2234
timestamp 0
transform -1 0 2491 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2235
timestamp 0
transform -1 0 2492 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2236
timestamp 0
transform -1 0 2493 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2237
timestamp 0
transform -1 0 2494 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2238
timestamp 0
transform -1 0 2495 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2239
timestamp 0
transform -1 0 2496 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2240
timestamp 0
transform -1 0 2497 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2241
timestamp 0
transform -1 0 2498 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2242
timestamp 0
transform -1 0 2499 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2243
timestamp 0
transform -1 0 2500 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2244
timestamp 0
transform -1 0 2501 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2245
timestamp 0
transform -1 0 2502 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2246
timestamp 0
transform -1 0 2503 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2247
timestamp 0
transform -1 0 2504 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2248
timestamp 0
transform -1 0 2505 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2249
timestamp 0
transform -1 0 2506 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2250
timestamp 0
transform -1 0 2507 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2251
timestamp 0
transform -1 0 2508 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2252
timestamp 0
transform -1 0 2509 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2253
timestamp 0
transform -1 0 2510 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2254
timestamp 0
transform -1 0 2511 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2255
timestamp 0
transform -1 0 2512 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2256
timestamp 0
transform -1 0 2513 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2257
timestamp 0
transform -1 0 2514 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2258
timestamp 0
transform -1 0 2515 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2259
timestamp 0
transform -1 0 2516 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2260
timestamp 0
transform -1 0 2517 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2261
timestamp 0
transform -1 0 2518 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2262
timestamp 0
transform -1 0 2519 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2263
timestamp 0
transform -1 0 2520 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2264
timestamp 0
transform -1 0 2521 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2265
timestamp 0
transform -1 0 2522 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2266
timestamp 0
transform -1 0 2523 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2267
timestamp 0
transform -1 0 2524 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2268
timestamp 0
transform -1 0 2525 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2269
timestamp 0
transform -1 0 2526 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2270
timestamp 0
transform -1 0 2527 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2271
timestamp 0
transform -1 0 2528 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2272
timestamp 0
transform -1 0 2529 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2273
timestamp 0
transform -1 0 2530 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2274
timestamp 0
transform -1 0 2531 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2275
timestamp 0
transform -1 0 2532 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2276
timestamp 0
transform -1 0 2533 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2277
timestamp 0
transform -1 0 2534 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2278
timestamp 0
transform -1 0 2535 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2279
timestamp 0
transform -1 0 2536 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2280
timestamp 0
transform -1 0 2537 0 -1 198
box 0 0 1 1
use s8iom0s8_com_bus_slice_1um  FILLER_2281
timestamp 0
transform -1 0 2538 0 -1 198
box 0 0 1 1
<< end >>
