VERSION 5.3 ;
   NAMESCASESENSITIVE ON ;
   NOWIREEXTENSIONATPIN ON ;
   DIVIDERCHAR "/" ;
   BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO lvlshiftdown
   CLASS BLOCK ;
   FOREIGN lvlshiftdown ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 9.6000 BY 4.0700 ;
   PIN vnb
      PORT
         LAYER li1 ;
	    RECT 0.0000 -0.0850 9.6000 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.1150 9.6000 0.1150 ;
      END
   END vnb
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.6150 3.6250 9.5050 3.7950 ;
	    RECT 0.6150 2.4450 1.8650 3.6250 ;
	    RECT 2.7650 2.3850 3.4350 3.6250 ;
	    RECT 4.1050 2.3850 4.9950 3.6250 ;
	    RECT 5.6650 2.3850 6.5550 3.6250 ;
	    RECT 7.2250 2.3850 8.1150 3.6250 ;
	    RECT 8.9050 3.4750 9.5050 3.6250 ;
	    RECT 9.1350 2.3850 9.5050 3.4750 ;
         LAYER met1 ;
	    RECT 0.0000 3.4450 9.6000 3.8150 ;
      END
   END vpwr
   PIN vpb
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.9850 9.6000 4.1550 ;
         LAYER met1 ;
	    RECT 0.0000 3.9550 9.6000 4.1850 ;
      END
   END vpb
   PIN vpb
   END vpb
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.6750 0.5500 1.9250 1.3850 ;
	    RECT 2.7650 0.7600 3.4950 1.4450 ;
	    RECT 2.6050 0.5500 3.4950 0.7600 ;
	    RECT 4.0450 0.5500 5.0550 1.4450 ;
	    RECT 5.6050 0.5500 6.6150 1.4450 ;
	    RECT 7.1650 0.5500 8.1750 1.4450 ;
	    RECT 9.1350 0.6000 9.5050 1.4450 ;
	    RECT 8.9750 0.5500 9.5050 0.6000 ;
	    RECT 0.6750 0.3800 9.5050 0.5500 ;
         LAYER met1 ;
	    RECT 0.0000 0.2550 9.6000 0.6250 ;
      END
   END vgnd
   PIN vnb
   END vnb
   PIN X
      PORT
         LAYER li1 ;
	    RECT 3.6050 2.2050 3.9350 3.4450 ;
	    RECT 5.1650 2.2050 5.4950 3.4450 ;
	    RECT 6.7250 2.2050 7.0550 3.4450 ;
	    RECT 8.2850 3.2300 8.7350 3.4450 ;
	    RECT 8.2850 2.2050 8.9650 3.2300 ;
	    RECT 3.6050 2.0350 8.9650 2.2050 ;
	    RECT 3.6650 1.6250 8.5550 1.7950 ;
	    RECT 3.6650 0.8050 3.8750 1.6250 ;
	    RECT 5.2250 0.8050 5.4350 1.6250 ;
	    RECT 6.7850 0.8050 6.9950 1.6250 ;
	    RECT 8.3450 0.9750 8.5550 1.6250 ;
	    RECT 8.7350 0.9750 8.9650 2.0350 ;
	    RECT 8.3450 0.8050 8.9650 0.9750 ;
      END
   END X
   PIN X
   END X
   PIN X
   END X
   PIN X
   END X
   PIN X
   END X
   PIN X
   END X
   PIN X
   END X
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.6350 1.5800 2.2450 1.8150 ;
      END
   END A
   PIN A
   END A
   PIN A
   END A
   PIN A
   END A
   OBS
         LAYER li1 ;
	    RECT 0.2450 2.2650 0.4350 3.5450 ;
	    RECT 2.0450 2.2650 2.5950 3.4450 ;
	    RECT 0.2450 2.0950 2.5950 2.2650 ;
	    RECT 0.2450 1.4750 0.4350 2.0950 ;
	    RECT 2.4250 1.9550 2.5950 2.0950 ;
	    RECT 2.4250 1.6250 3.3800 1.9550 ;
	    RECT 0.2450 0.8050 0.4550 1.4750 ;
	    RECT 2.4250 1.4000 2.5950 1.6250 ;
	    RECT 2.1050 1.2300 2.5950 1.4000 ;
	    RECT 2.1050 0.7300 2.3150 1.2300 ;
   END
END lvlshiftdown
