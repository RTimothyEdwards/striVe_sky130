magic
tech sky130A
magscale 1 2
timestamp 1586549559
<< checkpaint >>
rect -860 -908 28524 28364
<< locali >>
rect 24349 21191 24383 21497
rect 1901 16295 1935 16465
rect 3557 12045 3683 12079
rect 17725 9767 17759 9869
rect 18645 9767 18679 9937
rect 14413 7727 14447 7829
rect 10365 6129 10399 6265
rect 6593 5619 6627 5721
rect 11745 4327 11779 4429
<< viali >>
rect 6225 26733 6259 26767
rect 6777 26733 6811 26767
rect 6685 26665 6719 26699
rect 7513 26597 7547 26631
rect 23889 26597 23923 26631
rect 6685 26393 6719 26427
rect 23337 26393 23371 26427
rect 2545 26325 2579 26359
rect 18369 26325 18403 26359
rect 3005 26257 3039 26291
rect 3649 26257 3683 26291
rect 7145 26257 7179 26291
rect 8433 26257 8467 26291
rect 14505 26257 14539 26291
rect 14873 26257 14907 26291
rect 22233 26257 22267 26291
rect 24073 26257 24107 26291
rect 25821 26257 25855 26291
rect 2177 26189 2211 26223
rect 3097 26189 3131 26223
rect 3833 26189 3867 26223
rect 7237 26189 7271 26223
rect 7513 26189 7547 26223
rect 8341 26189 8375 26223
rect 11745 26189 11779 26223
rect 12389 26189 12423 26223
rect 14321 26189 14355 26223
rect 14597 26189 14631 26223
rect 15977 26189 16011 26223
rect 17725 26189 17759 26223
rect 19933 26189 19967 26223
rect 21589 26189 21623 26223
rect 23797 26189 23831 26223
rect 3557 26121 3591 26155
rect 7605 26121 7639 26155
rect 11561 26121 11595 26155
rect 12205 26121 12239 26155
rect 12297 26121 12331 26155
rect 12573 26121 12607 26155
rect 16069 26121 16103 26155
rect 16161 26121 16195 26155
rect 18001 26121 18035 26155
rect 20025 26121 20059 26155
rect 20117 26121 20151 26155
rect 21865 26121 21899 26155
rect 22325 26121 22359 26155
rect 1993 26053 2027 26087
rect 2269 26053 2303 26087
rect 4017 26053 4051 26087
rect 6225 26053 6259 26087
rect 6501 26053 6535 26087
rect 16437 26053 16471 26087
rect 18461 26053 18495 26087
rect 20393 26053 20427 26087
rect 23521 26053 23555 26087
rect 23705 26053 23739 26087
rect 7421 25849 7455 25883
rect 2085 25781 2119 25815
rect 9353 25781 9387 25815
rect 11745 25781 11779 25815
rect 14873 25781 14907 25815
rect 1165 25713 1199 25747
rect 1901 25713 1935 25747
rect 3373 25713 3407 25747
rect 4293 25713 4327 25747
rect 6685 25713 6719 25747
rect 6777 25713 6811 25747
rect 7881 25713 7915 25747
rect 10089 25713 10123 25747
rect 10181 25713 10215 25747
rect 12481 25713 12515 25747
rect 17449 25713 17483 25747
rect 18829 25713 18863 25747
rect 5857 25645 5891 25679
rect 5949 25645 5983 25679
rect 9261 25645 9295 25679
rect 11653 25645 11687 25679
rect 12573 25645 12607 25679
rect 14597 25645 14631 25679
rect 16621 25645 16655 25679
rect 18001 25645 18035 25679
rect 18553 25645 18587 25679
rect 19013 25645 19047 25679
rect 20853 25645 20887 25679
rect 21129 25645 21163 25679
rect 22877 25645 22911 25679
rect 4661 25577 4695 25611
rect 20669 25577 20703 25611
rect 7697 25509 7731 25543
rect 8249 25509 8283 25543
rect 17909 25509 17943 25543
rect 20485 25509 20519 25543
rect 23981 25509 24015 25543
rect 2637 25305 2671 25339
rect 3005 25305 3039 25339
rect 3373 25305 3407 25339
rect 3833 25305 3867 25339
rect 5673 25305 5707 25339
rect 7789 25305 7823 25339
rect 8985 25305 9019 25339
rect 11377 25305 11411 25339
rect 14689 25305 14723 25339
rect 15885 25305 15919 25339
rect 16805 25305 16839 25339
rect 19473 25305 19507 25339
rect 21957 25305 21991 25339
rect 22233 25305 22267 25339
rect 10549 25237 10583 25271
rect 14321 25237 14355 25271
rect 15701 25237 15735 25271
rect 20209 25237 20243 25271
rect 20393 25237 20427 25271
rect 21129 25237 21163 25271
rect 1073 25169 1107 25203
rect 1717 25169 1751 25203
rect 9077 25169 9111 25203
rect 14873 25169 14907 25203
rect 15333 25169 15367 25203
rect 16989 25169 17023 25203
rect 17173 25169 17207 25203
rect 17633 25169 17667 25203
rect 19933 25169 19967 25203
rect 21773 25169 21807 25203
rect 25913 25169 25947 25203
rect 1165 25101 1199 25135
rect 1809 25101 1843 25135
rect 1993 25101 2027 25135
rect 5305 25101 5339 25135
rect 6225 25101 6259 25135
rect 6869 25101 6903 25135
rect 7237 25101 7271 25135
rect 9261 25101 9295 25135
rect 10181 25101 10215 25135
rect 10917 25101 10951 25135
rect 11745 25101 11779 25135
rect 12389 25101 12423 25135
rect 15057 25101 15091 25135
rect 17357 25101 17391 25135
rect 20485 25101 20519 25135
rect 20853 25101 20887 25135
rect 21497 25101 21531 25135
rect 23889 25101 23923 25135
rect 889 25033 923 25067
rect 1625 25033 1659 25067
rect 2545 25033 2579 25067
rect 2821 25033 2855 25067
rect 3649 25033 3683 25067
rect 7145 25033 7179 25067
rect 8065 25033 8099 25067
rect 8249 25033 8283 25067
rect 8525 25033 8559 25067
rect 8801 25033 8835 25067
rect 12665 25033 12699 25067
rect 14505 25033 14539 25067
rect 19381 25033 19415 25067
rect 24165 25033 24199 25067
rect 5397 24965 5431 24999
rect 5765 24965 5799 24999
rect 7605 24965 7639 24999
rect 8341 24965 8375 24999
rect 11101 24965 11135 24999
rect 11561 24965 11595 24999
rect 19657 24965 19691 24999
rect 23521 24965 23555 24999
rect 23797 24965 23831 24999
rect 889 24761 923 24795
rect 1349 24761 1383 24795
rect 6685 24761 6719 24795
rect 6961 24761 6995 24795
rect 7421 24761 7455 24795
rect 11745 24761 11779 24795
rect 11837 24761 11871 24795
rect 12113 24761 12147 24795
rect 12389 24761 12423 24795
rect 21681 24761 21715 24795
rect 23981 24761 24015 24795
rect 24165 24761 24199 24795
rect 1533 24693 1567 24727
rect 10457 24693 10491 24727
rect 11377 24693 11411 24727
rect 4201 24625 4235 24659
rect 6409 24625 6443 24659
rect 12573 24625 12607 24659
rect 14873 24625 14907 24659
rect 18461 24625 18495 24659
rect 18829 24625 18863 24659
rect 19013 24625 19047 24659
rect 21037 24625 21071 24659
rect 22601 24625 22635 24659
rect 24441 24625 24475 24659
rect 5581 24557 5615 24591
rect 5673 24557 5707 24591
rect 6501 24557 6535 24591
rect 9261 24557 9295 24591
rect 9445 24557 9479 24591
rect 9997 24557 10031 24591
rect 10549 24557 10583 24591
rect 15149 24557 15183 24591
rect 18369 24557 18403 24591
rect 20945 24557 20979 24591
rect 24717 24557 24751 24591
rect 20485 24489 20519 24523
rect 1073 24421 1107 24455
rect 4293 24421 4327 24455
rect 7513 24421 7547 24455
rect 7789 24421 7823 24455
rect 9629 24421 9663 24455
rect 11469 24421 11503 24455
rect 14689 24421 14723 24455
rect 17357 24421 17391 24455
rect 17909 24421 17943 24455
rect 20669 24421 20703 24455
rect 21221 24421 21255 24455
rect 22417 24421 22451 24455
rect 3005 24217 3039 24251
rect 3465 24217 3499 24251
rect 4293 24217 4327 24251
rect 6133 24217 6167 24251
rect 6869 24217 6903 24251
rect 7053 24217 7087 24251
rect 9997 24217 10031 24251
rect 10273 24217 10307 24251
rect 11745 24217 11779 24251
rect 12481 24217 12515 24251
rect 12573 24217 12607 24251
rect 18461 24217 18495 24251
rect 18553 24217 18587 24251
rect 22601 24217 22635 24251
rect 23613 24217 23647 24251
rect 4201 24149 4235 24183
rect 5857 24149 5891 24183
rect 7237 24149 7271 24183
rect 10457 24149 10491 24183
rect 11377 24149 11411 24183
rect 18277 24149 18311 24183
rect 20393 24149 20427 24183
rect 20669 24149 20703 24183
rect 22417 24149 22451 24183
rect 1073 24081 1107 24115
rect 1901 24081 1935 24115
rect 5765 24081 5799 24115
rect 14137 24081 14171 24115
rect 16437 24081 16471 24115
rect 17909 24081 17943 24115
rect 20301 24081 20335 24115
rect 981 24013 1015 24047
rect 1809 24013 1843 24047
rect 5489 24013 5523 24047
rect 7421 24013 7455 24047
rect 7513 24013 7547 24047
rect 8433 24013 8467 24047
rect 13953 24013 13987 24047
rect 14413 24013 14447 24047
rect 20117 24013 20151 24047
rect 20577 24013 20611 24047
rect 21129 24013 21163 24047
rect 21589 24013 21623 24047
rect 24257 24013 24291 24047
rect 24809 24013 24843 24047
rect 705 23945 739 23979
rect 2913 23945 2947 23979
rect 3189 23945 3223 23979
rect 9077 23945 9111 23979
rect 14689 23945 14723 23979
rect 23889 23945 23923 23979
rect 14321 23877 14355 23911
rect 18001 23877 18035 23911
rect 21773 23877 21807 23911
rect 24073 23877 24107 23911
rect 14965 23673 14999 23707
rect 15149 23673 15183 23707
rect 18369 23673 18403 23707
rect 21497 23673 21531 23707
rect 24533 23673 24567 23707
rect 8065 23605 8099 23639
rect 1257 23537 1291 23571
rect 1717 23537 1751 23571
rect 4201 23537 4235 23571
rect 5121 23537 5155 23571
rect 13309 23537 13343 23571
rect 13401 23537 13435 23571
rect 16069 23537 16103 23571
rect 18093 23537 18127 23571
rect 18645 23537 18679 23571
rect 20577 23537 20611 23571
rect 20669 23537 20703 23571
rect 1809 23469 1843 23503
rect 5765 23469 5799 23503
rect 7513 23469 7547 23503
rect 12481 23469 12515 23503
rect 12573 23469 12607 23503
rect 21221 23469 21255 23503
rect 7973 23401 8007 23435
rect 981 23333 1015 23367
rect 1993 23333 2027 23367
rect 16345 23333 16379 23367
rect 20853 23333 20887 23367
rect 24165 23333 24199 23367
rect 889 23129 923 23163
rect 1073 23129 1107 23163
rect 4201 23129 4235 23163
rect 5397 23129 5431 23163
rect 7697 23129 7731 23163
rect 13309 23129 13343 23163
rect 16713 23129 16747 23163
rect 18369 23129 18403 23163
rect 18829 23129 18863 23163
rect 19381 23129 19415 23163
rect 20577 23129 20611 23163
rect 20945 23129 20979 23163
rect 2913 23061 2947 23095
rect 3189 23061 3223 23095
rect 3925 23061 3959 23095
rect 9537 23061 9571 23095
rect 9813 23061 9847 23095
rect 4661 22993 4695 23027
rect 7513 22993 7547 23027
rect 12389 22993 12423 23027
rect 13401 22993 13435 23027
rect 24165 22993 24199 23027
rect 26189 22993 26223 23027
rect 1165 22925 1199 22959
rect 2085 22925 2119 22959
rect 3097 22925 3131 22959
rect 3373 22925 3407 22959
rect 4109 22925 4143 22959
rect 4569 22925 4603 22959
rect 5121 22925 5155 22959
rect 7973 22925 8007 22959
rect 10457 22925 10491 22959
rect 10733 22925 10767 22959
rect 12573 22925 12607 22959
rect 13033 22925 13067 22959
rect 13585 22925 13619 22959
rect 16069 22925 16103 22959
rect 16897 22925 16931 22959
rect 17909 22925 17943 22959
rect 18553 22925 18587 22959
rect 18645 22925 18679 22959
rect 1901 22857 1935 22891
rect 5213 22857 5247 22891
rect 5489 22857 5523 22891
rect 9353 22857 9387 22891
rect 9629 22857 9663 22891
rect 10641 22857 10675 22891
rect 10917 22857 10951 22891
rect 11929 22857 11963 22891
rect 13125 22857 13159 22891
rect 16437 22857 16471 22891
rect 16529 22857 16563 22891
rect 18185 22857 18219 22891
rect 19289 22857 19323 22891
rect 24073 22857 24107 22891
rect 24441 22857 24475 22891
rect 2177 22789 2211 22823
rect 2361 22789 2395 22823
rect 12021 22789 12055 22823
rect 12297 22789 12331 22823
rect 15977 22789 16011 22823
rect 20853 22789 20887 22823
rect 23889 22789 23923 22823
rect 1349 22585 1383 22619
rect 2177 22585 2211 22619
rect 18553 22585 18587 22619
rect 24257 22585 24291 22619
rect 1073 22517 1107 22551
rect 1901 22517 1935 22551
rect 5213 22517 5247 22551
rect 24717 22517 24751 22551
rect 4201 22449 4235 22483
rect 4385 22449 4419 22483
rect 5029 22449 5063 22483
rect 11009 22449 11043 22483
rect 11837 22449 11871 22483
rect 12757 22449 12791 22483
rect 16345 22449 16379 22483
rect 16897 22449 16931 22483
rect 20209 22449 20243 22483
rect 21773 22449 21807 22483
rect 22785 22449 22819 22483
rect 24441 22449 24475 22483
rect 1441 22381 1475 22415
rect 1993 22381 2027 22415
rect 13401 22381 13435 22415
rect 16437 22381 16471 22415
rect 16805 22381 16839 22415
rect 20485 22381 20519 22415
rect 22693 22381 22727 22415
rect 16529 22313 16563 22347
rect 23429 22313 23463 22347
rect 4017 22245 4051 22279
rect 7789 22245 7823 22279
rect 10825 22245 10859 22279
rect 15425 22245 15459 22279
rect 19105 22245 19139 22279
rect 21773 22245 21807 22279
rect 22969 22245 23003 22279
rect 23521 22245 23555 22279
rect 23797 22245 23831 22279
rect 4017 22041 4051 22075
rect 5489 22041 5523 22075
rect 7513 22041 7547 22075
rect 11377 22041 11411 22075
rect 13585 22041 13619 22075
rect 13953 22041 13987 22075
rect 15241 22041 15275 22075
rect 16529 22041 16563 22075
rect 21589 22041 21623 22075
rect 22785 22041 22819 22075
rect 2269 21973 2303 22007
rect 3833 21973 3867 22007
rect 7329 21973 7363 22007
rect 13217 21973 13251 22007
rect 13309 21973 13343 22007
rect 15425 21973 15459 22007
rect 16713 21973 16747 22007
rect 22417 21973 22451 22007
rect 7881 21905 7915 21939
rect 8709 21905 8743 21939
rect 10181 21905 10215 21939
rect 10825 21905 10859 21939
rect 11101 21905 11135 21939
rect 13033 21905 13067 21939
rect 14873 21905 14907 21939
rect 16161 21905 16195 21939
rect 17357 21905 17391 21939
rect 18001 21905 18035 21939
rect 18829 21905 18863 21939
rect 23245 21905 23279 21939
rect 25269 21905 25303 21939
rect 981 21837 1015 21871
rect 2085 21837 2119 21871
rect 4201 21837 4235 21871
rect 4293 21837 4327 21871
rect 5213 21837 5247 21871
rect 6225 21837 6259 21871
rect 6501 21837 6535 21871
rect 7789 21837 7823 21871
rect 8586 21837 8620 21871
rect 10273 21837 10307 21871
rect 11009 21837 11043 21871
rect 11561 21837 11595 21871
rect 11745 21837 11779 21871
rect 12665 21837 12699 21871
rect 15057 21837 15091 21871
rect 15333 21837 15367 21871
rect 15885 21837 15919 21871
rect 17449 21837 17483 21871
rect 18185 21837 18219 21871
rect 19105 21837 19139 21871
rect 4937 21769 4971 21803
rect 5305 21769 5339 21803
rect 9997 21769 10031 21803
rect 10733 21769 10767 21803
rect 12389 21769 12423 21803
rect 13493 21769 13527 21803
rect 13769 21769 13803 21803
rect 17081 21769 17115 21803
rect 17909 21769 17943 21803
rect 19013 21769 19047 21803
rect 19381 21769 19415 21803
rect 21129 21769 21163 21803
rect 23153 21769 23187 21803
rect 23521 21769 23555 21803
rect 889 21701 923 21735
rect 6317 21701 6351 21735
rect 6685 21701 6719 21735
rect 12757 21701 12791 21735
rect 21773 21701 21807 21735
rect 22601 21701 22635 21735
rect 1717 21497 1751 21531
rect 1993 21497 2027 21531
rect 4293 21497 4327 21531
rect 7697 21497 7731 21531
rect 10917 21497 10951 21531
rect 15425 21497 15459 21531
rect 16161 21497 16195 21531
rect 20485 21497 20519 21531
rect 24349 21497 24383 21531
rect 24717 21497 24751 21531
rect 1073 21429 1107 21463
rect 5029 21429 5063 21463
rect 12021 21429 12055 21463
rect 15977 21429 16011 21463
rect 20301 21429 20335 21463
rect 22693 21429 22727 21463
rect 1901 21361 1935 21395
rect 5121 21361 5155 21395
rect 9261 21361 9295 21395
rect 9445 21361 9479 21395
rect 12757 21361 12791 21395
rect 16437 21361 16471 21395
rect 16713 21361 16747 21395
rect 17173 21361 17207 21395
rect 17265 21361 17299 21395
rect 21313 21361 21347 21395
rect 21681 21361 21715 21395
rect 23337 21361 23371 21395
rect 23705 21361 23739 21395
rect 4569 21293 4603 21327
rect 11924 21293 11958 21327
rect 12849 21293 12883 21327
rect 21221 21293 21255 21327
rect 21773 21293 21807 21327
rect 23245 21293 23279 21327
rect 23797 21293 23831 21327
rect 16897 21225 16931 21259
rect 1441 21157 1475 21191
rect 9537 21157 9571 21191
rect 13585 21157 13619 21191
rect 19197 21157 19231 21191
rect 20761 21157 20795 21191
rect 24349 21157 24383 21191
rect 24533 21157 24567 21191
rect 1901 20953 1935 20987
rect 2085 20953 2119 20987
rect 4753 20953 4787 20987
rect 4937 20953 4971 20987
rect 9445 20953 9479 20987
rect 9629 20953 9663 20987
rect 12205 20953 12239 20987
rect 13309 20953 13343 20987
rect 16345 20953 16379 20987
rect 16713 20953 16747 20987
rect 19933 20953 19967 20987
rect 20301 20953 20335 20987
rect 21129 20953 21163 20987
rect 22785 20953 22819 20987
rect 23521 20953 23555 20987
rect 12113 20885 12147 20919
rect 16989 20885 17023 20919
rect 4661 20817 4695 20851
rect 13217 20817 13251 20851
rect 16529 20817 16563 20851
rect 24901 20817 24935 20851
rect 25361 20817 25395 20851
rect 7605 20749 7639 20783
rect 13585 20749 13619 20783
rect 14413 20749 14447 20783
rect 14505 20749 14539 20783
rect 20117 20749 20151 20783
rect 20577 20749 20611 20783
rect 21405 20749 21439 20783
rect 24625 20749 24659 20783
rect 7421 20681 7455 20715
rect 8249 20681 8283 20715
rect 9353 20681 9387 20715
rect 12389 20681 12423 20715
rect 13033 20681 13067 20715
rect 13677 20681 13711 20715
rect 20945 20681 20979 20715
rect 23061 20681 23095 20715
rect 7329 20613 7363 20647
rect 7697 20613 7731 20647
rect 8157 20613 8191 20647
rect 11837 20613 11871 20647
rect 16805 20613 16839 20647
rect 20669 20613 20703 20647
rect 21313 20613 21347 20647
rect 23153 20613 23187 20647
rect 23337 20613 23371 20647
rect 25177 20613 25211 20647
rect 6133 20409 6167 20443
rect 8157 20409 8191 20443
rect 23797 20409 23831 20443
rect 9997 20341 10031 20375
rect 21773 20341 21807 20375
rect 889 20273 923 20307
rect 1625 20273 1659 20307
rect 4109 20273 4143 20307
rect 4293 20273 4327 20307
rect 5489 20273 5523 20307
rect 7053 20273 7087 20307
rect 9445 20273 9479 20307
rect 9629 20273 9663 20307
rect 13493 20273 13527 20307
rect 16069 20273 16103 20307
rect 16805 20273 16839 20307
rect 20209 20273 20243 20307
rect 21865 20273 21899 20307
rect 797 20205 831 20239
rect 1717 20205 1751 20239
rect 5636 20205 5670 20239
rect 5857 20205 5891 20239
rect 7421 20205 7455 20239
rect 7697 20205 7731 20239
rect 7329 20137 7363 20171
rect 13677 20137 13711 20171
rect 4385 20069 4419 20103
rect 5765 20069 5799 20103
rect 7191 20069 7225 20103
rect 7881 20069 7915 20103
rect 20485 20069 20519 20103
rect 21589 20069 21623 20103
rect 22049 20069 22083 20103
rect 889 19865 923 19899
rect 1257 19865 1291 19899
rect 1717 19865 1751 19899
rect 2085 19865 2119 19899
rect 5489 19865 5523 19899
rect 6225 19865 6259 19899
rect 6409 19865 6443 19899
rect 6777 19865 6811 19899
rect 7329 19865 7363 19899
rect 7697 19865 7731 19899
rect 8525 19865 8559 19899
rect 8709 19865 8743 19899
rect 9261 19865 9295 19899
rect 9997 19865 10031 19899
rect 10273 19865 10307 19899
rect 13493 19865 13527 19899
rect 15609 19865 15643 19899
rect 15885 19865 15919 19899
rect 19933 19865 19967 19899
rect 20485 19865 20519 19899
rect 21037 19865 21071 19899
rect 21773 19865 21807 19899
rect 22141 19865 22175 19899
rect 1073 19797 1107 19831
rect 6501 19797 6535 19831
rect 7559 19797 7593 19831
rect 8341 19797 8375 19831
rect 15517 19797 15551 19831
rect 20025 19797 20059 19831
rect 21681 19797 21715 19831
rect 7789 19729 7823 19763
rect 8157 19729 8191 19763
rect 18369 19729 18403 19763
rect 20209 19729 20243 19763
rect 23797 19729 23831 19763
rect 6869 19661 6903 19695
rect 7421 19661 7455 19695
rect 9169 19661 9203 19695
rect 9629 19661 9663 19695
rect 18461 19661 18495 19695
rect 19197 19661 19231 19695
rect 20301 19661 20335 19695
rect 20945 19661 20979 19695
rect 1625 19593 1659 19627
rect 4569 19593 4603 19627
rect 5765 19593 5799 19627
rect 8893 19593 8927 19627
rect 8985 19593 9019 19627
rect 9813 19593 9847 19627
rect 18921 19593 18955 19627
rect 19105 19593 19139 19627
rect 22049 19593 22083 19627
rect 23521 19593 23555 19627
rect 24073 19593 24107 19627
rect 25821 19593 25855 19627
rect 705 19525 739 19559
rect 1993 19525 2027 19559
rect 4201 19525 4235 19559
rect 4293 19525 4327 19559
rect 5949 19525 5983 19559
rect 7145 19525 7179 19559
rect 13677 19525 13711 19559
rect 18185 19525 18219 19559
rect 23245 19525 23279 19559
rect 23705 19525 23739 19559
rect 1349 19321 1383 19355
rect 7145 19321 7179 19355
rect 19657 19321 19691 19355
rect 20209 19321 20243 19355
rect 23061 19321 23095 19355
rect 4661 19253 4695 19287
rect 8065 19253 8099 19287
rect 17449 19253 17483 19287
rect 23429 19253 23463 19287
rect 4845 19185 4879 19219
rect 7605 19185 7639 19219
rect 10457 19185 10491 19219
rect 11101 19185 11135 19219
rect 12665 19185 12699 19219
rect 13493 19185 13527 19219
rect 18369 19185 18403 19219
rect 18737 19185 18771 19219
rect 18921 19185 18955 19219
rect 22233 19185 22267 19219
rect 23521 19185 23555 19219
rect 26097 19185 26131 19219
rect 7513 19117 7547 19151
rect 10733 19117 10767 19151
rect 11009 19117 11043 19151
rect 12757 19117 12791 19151
rect 13585 19117 13619 19151
rect 18185 19117 18219 19151
rect 21405 19117 21439 19151
rect 21957 19117 21991 19151
rect 22417 19117 22451 19151
rect 10457 19049 10491 19083
rect 17633 19049 17667 19083
rect 4937 18981 4971 19015
rect 13861 18981 13895 19015
rect 18001 18981 18035 19015
rect 23245 18981 23279 19015
rect 23705 18981 23739 19015
rect 26097 18981 26131 19015
rect 3005 18777 3039 18811
rect 3465 18777 3499 18811
rect 4385 18777 4419 18811
rect 4569 18777 4603 18811
rect 6961 18777 6995 18811
rect 7145 18777 7179 18811
rect 7697 18777 7731 18811
rect 8801 18777 8835 18811
rect 9261 18777 9295 18811
rect 10365 18777 10399 18811
rect 12849 18777 12883 18811
rect 19381 18777 19415 18811
rect 21957 18777 21991 18811
rect 22601 18777 22635 18811
rect 24993 18777 25027 18811
rect 25913 18777 25947 18811
rect 5489 18709 5523 18743
rect 7329 18709 7363 18743
rect 8065 18709 8099 18743
rect 8341 18709 8375 18743
rect 17173 18709 17207 18743
rect 17725 18709 17759 18743
rect 19013 18709 19047 18743
rect 19289 18709 19323 18743
rect 19657 18709 19691 18743
rect 21497 18709 21531 18743
rect 22785 18709 22819 18743
rect 2269 18641 2303 18675
rect 7789 18641 7823 18675
rect 10825 18641 10859 18675
rect 11285 18641 11319 18675
rect 14229 18641 14263 18675
rect 16989 18641 17023 18675
rect 18645 18641 18679 18675
rect 21865 18641 21899 18675
rect 22233 18641 22267 18675
rect 22969 18641 23003 18675
rect 23521 18641 23555 18675
rect 25361 18641 25395 18675
rect 1349 18573 1383 18607
rect 2177 18573 2211 18607
rect 3373 18573 3407 18607
rect 3833 18573 3867 18607
rect 4661 18573 4695 18607
rect 4845 18573 4879 18607
rect 7568 18573 7602 18607
rect 8985 18573 9019 18607
rect 9169 18573 9203 18607
rect 9629 18573 9663 18607
rect 10733 18573 10767 18607
rect 11101 18573 11135 18607
rect 12481 18573 12515 18607
rect 13217 18573 13251 18607
rect 13861 18573 13895 18607
rect 15609 18573 15643 18607
rect 16161 18573 16195 18607
rect 17909 18573 17943 18607
rect 18001 18573 18035 18607
rect 18369 18573 18403 18607
rect 19749 18573 19783 18607
rect 20117 18573 20151 18607
rect 20393 18573 20427 18607
rect 23613 18573 23647 18607
rect 23981 18573 24015 18607
rect 24165 18573 24199 18607
rect 25177 18573 25211 18607
rect 1073 18505 1107 18539
rect 1441 18505 1475 18539
rect 3189 18505 3223 18539
rect 6777 18505 6811 18539
rect 7421 18505 7455 18539
rect 10181 18505 10215 18539
rect 14137 18505 14171 18539
rect 15885 18505 15919 18539
rect 16345 18505 16379 18539
rect 16805 18505 16839 18539
rect 21681 18505 21715 18539
rect 889 18437 923 18471
rect 4109 18437 4143 18471
rect 4937 18437 4971 18471
rect 5397 18437 5431 18471
rect 8709 18437 8743 18471
rect 9997 18437 10031 18471
rect 10917 18437 10951 18471
rect 12573 18437 12607 18471
rect 12941 18437 12975 18471
rect 18829 18437 18863 18471
rect 22417 18437 22451 18471
rect 24257 18437 24291 18471
rect 26005 18437 26039 18471
rect 26189 18437 26223 18471
rect 4937 18233 4971 18267
rect 6593 18233 6627 18267
rect 7881 18233 7915 18267
rect 10181 18233 10215 18267
rect 18185 18233 18219 18267
rect 19657 18233 19691 18267
rect 22969 18233 23003 18267
rect 23337 18233 23371 18267
rect 13585 18165 13619 18199
rect 15793 18165 15827 18199
rect 18001 18165 18035 18199
rect 18737 18165 18771 18199
rect 20209 18165 20243 18199
rect 23797 18165 23831 18199
rect 4109 18097 4143 18131
rect 6317 18097 6351 18131
rect 6501 18097 6535 18131
rect 9261 18097 9295 18131
rect 9445 18097 9479 18131
rect 11009 18097 11043 18131
rect 13125 18097 13159 18131
rect 17541 18097 17575 18131
rect 18645 18097 18679 18131
rect 20393 18097 20427 18131
rect 23429 18097 23463 18131
rect 4477 18029 4511 18063
rect 7513 18029 7547 18063
rect 13677 18029 13711 18063
rect 15517 18029 15551 18063
rect 17817 18029 17851 18063
rect 20761 18029 20795 18063
rect 705 17893 739 17927
rect 889 17893 923 17927
rect 1257 17893 1291 17927
rect 4247 17893 4281 17927
rect 4385 17893 4419 17927
rect 4569 17893 4603 17927
rect 5121 17893 5155 17927
rect 7605 17893 7639 17927
rect 9537 17893 9571 17927
rect 10825 17893 10859 17927
rect 13861 17893 13895 17927
rect 23981 17893 24015 17927
rect 4201 17689 4235 17723
rect 5581 17689 5615 17723
rect 5765 17689 5799 17723
rect 6869 17689 6903 17723
rect 7789 17689 7823 17723
rect 8433 17689 8467 17723
rect 9813 17689 9847 17723
rect 13125 17689 13159 17723
rect 13585 17689 13619 17723
rect 15793 17689 15827 17723
rect 18461 17689 18495 17723
rect 20301 17689 20335 17723
rect 23797 17689 23831 17723
rect 24257 17689 24291 17723
rect 24625 17689 24659 17723
rect 24901 17689 24935 17723
rect 5397 17621 5431 17655
rect 13401 17621 13435 17655
rect 13953 17621 13987 17655
rect 14229 17621 14263 17655
rect 16161 17621 16195 17655
rect 18645 17621 18679 17655
rect 797 17553 831 17587
rect 889 17553 923 17587
rect 4293 17553 4327 17587
rect 5949 17553 5983 17587
rect 10181 17553 10215 17587
rect 15609 17553 15643 17587
rect 20393 17553 20427 17587
rect 1625 17485 1659 17519
rect 1717 17485 1751 17519
rect 3465 17485 3499 17519
rect 4845 17485 4879 17519
rect 6317 17485 6351 17519
rect 6685 17485 6719 17519
rect 8341 17485 8375 17519
rect 9721 17485 9755 17519
rect 10917 17485 10951 17519
rect 14137 17485 14171 17519
rect 14413 17485 14447 17519
rect 20117 17485 20151 17519
rect 20761 17485 20795 17519
rect 21129 17485 21163 17519
rect 22785 17485 22819 17519
rect 23245 17485 23279 17519
rect 24441 17485 24475 17519
rect 3189 17417 3223 17451
rect 3281 17417 3315 17451
rect 4661 17417 4695 17451
rect 6133 17417 6167 17451
rect 6961 17417 6995 17451
rect 8157 17417 8191 17451
rect 9169 17417 9203 17451
rect 9537 17417 9571 17451
rect 10365 17417 10399 17451
rect 21037 17417 21071 17451
rect 21313 17417 21347 17451
rect 23337 17417 23371 17451
rect 23613 17417 23647 17451
rect 3005 17349 3039 17383
rect 3557 17349 3591 17383
rect 4017 17349 4051 17383
rect 4569 17349 4603 17383
rect 4937 17349 4971 17383
rect 7237 17349 7271 17383
rect 7973 17349 8007 17383
rect 8893 17349 8927 17383
rect 9353 17349 9387 17383
rect 10825 17349 10859 17383
rect 15977 17349 16011 17383
rect 23521 17349 23555 17383
rect 981 17145 1015 17179
rect 2637 17145 2671 17179
rect 4293 17145 4327 17179
rect 4569 17145 4603 17179
rect 9353 17145 9387 17179
rect 14597 17145 14631 17179
rect 1717 17077 1751 17111
rect 5489 17077 5523 17111
rect 5673 17009 5707 17043
rect 6869 17009 6903 17043
rect 7053 17009 7087 17043
rect 11561 17009 11595 17043
rect 12305 17009 12339 17043
rect 15793 17009 15827 17043
rect 16345 17009 16379 17043
rect 20853 17009 20887 17043
rect 20945 17009 20979 17043
rect 21221 17009 21255 17043
rect 25821 17009 25855 17043
rect 2085 16941 2119 16975
rect 4109 16941 4143 16975
rect 9537 16941 9571 16975
rect 11469 16941 11503 16975
rect 12389 16941 12423 16975
rect 16529 16941 16563 16975
rect 21313 16941 21347 16975
rect 2177 16873 2211 16907
rect 6409 16873 6443 16907
rect 23061 16873 23095 16907
rect 705 16805 739 16839
rect 1855 16805 1889 16839
rect 1993 16805 2027 16839
rect 5765 16805 5799 16839
rect 7145 16805 7179 16839
rect 8433 16805 8467 16839
rect 14689 16805 14723 16839
rect 15425 16805 15459 16839
rect 17817 16805 17851 16839
rect 20301 16805 20335 16839
rect 23153 16805 23187 16839
rect 24993 16805 25027 16839
rect 26005 16805 26039 16839
rect 1165 16601 1199 16635
rect 1809 16601 1843 16635
rect 2269 16601 2303 16635
rect 2637 16601 2671 16635
rect 3557 16601 3591 16635
rect 4477 16601 4511 16635
rect 5581 16601 5615 16635
rect 5857 16601 5891 16635
rect 7053 16601 7087 16635
rect 9169 16601 9203 16635
rect 11101 16601 11135 16635
rect 14597 16601 14631 16635
rect 14781 16601 14815 16635
rect 15149 16601 15183 16635
rect 20485 16601 20519 16635
rect 20669 16601 20703 16635
rect 20853 16601 20887 16635
rect 22785 16601 22819 16635
rect 24809 16601 24843 16635
rect 26465 16601 26499 16635
rect 3925 16533 3959 16567
rect 4293 16533 4327 16567
rect 4937 16533 4971 16567
rect 15057 16533 15091 16567
rect 19013 16533 19047 16567
rect 20301 16533 20335 16567
rect 21037 16533 21071 16567
rect 21589 16533 21623 16567
rect 23245 16533 23279 16567
rect 26373 16533 26407 16567
rect 1901 16465 1935 16499
rect 2508 16465 2542 16499
rect 2729 16465 2763 16499
rect 3189 16465 3223 16499
rect 3741 16465 3775 16499
rect 4385 16465 4419 16499
rect 9077 16465 9111 16499
rect 12757 16465 12791 16499
rect 15425 16465 15459 16499
rect 16345 16465 16379 16499
rect 22417 16465 22451 16499
rect 24993 16465 25027 16499
rect 25729 16465 25763 16499
rect 25913 16465 25947 16499
rect 1441 16397 1475 16431
rect 2361 16397 2395 16431
rect 4017 16397 4051 16431
rect 4164 16397 4198 16431
rect 7973 16397 8007 16431
rect 8525 16397 8559 16431
rect 11837 16397 11871 16431
rect 12665 16397 12699 16431
rect 16253 16397 16287 16431
rect 16529 16397 16563 16431
rect 17633 16397 17667 16431
rect 18737 16397 18771 16431
rect 19105 16397 19139 16431
rect 21221 16397 21255 16431
rect 23429 16397 23463 16431
rect 23613 16397 23647 16431
rect 23981 16397 24015 16431
rect 24073 16397 24107 16431
rect 25637 16397 25671 16431
rect 26005 16397 26039 16431
rect 6869 16329 6903 16363
rect 8341 16329 8375 16363
rect 8709 16329 8743 16363
rect 11929 16329 11963 16363
rect 15517 16329 15551 16363
rect 17449 16329 17483 16363
rect 22601 16329 22635 16363
rect 24533 16329 24567 16363
rect 1533 16261 1567 16295
rect 1901 16261 1935 16295
rect 1993 16261 2027 16295
rect 3005 16261 3039 16295
rect 5765 16261 5799 16295
rect 7237 16261 7271 16295
rect 8249 16261 8283 16295
rect 8617 16261 8651 16295
rect 10641 16261 10675 16295
rect 10917 16261 10951 16295
rect 11193 16261 11227 16295
rect 11469 16261 11503 16295
rect 16713 16261 16747 16295
rect 20025 16261 20059 16295
rect 21497 16261 21531 16295
rect 24717 16261 24751 16295
rect 1717 16057 1751 16091
rect 4109 16057 4143 16091
rect 8433 16057 8467 16091
rect 9445 16057 9479 16091
rect 12113 16057 12147 16091
rect 15885 16057 15919 16091
rect 25085 16057 25119 16091
rect 6041 15989 6075 16023
rect 6225 15989 6259 16023
rect 6593 15989 6627 16023
rect 9537 15989 9571 16023
rect 11837 15989 11871 16023
rect 1901 15921 1935 15955
rect 2085 15921 2119 15955
rect 6133 15921 6167 15955
rect 9353 15921 9387 15955
rect 11377 15921 11411 15955
rect 16621 15921 16655 15955
rect 16989 15921 17023 15955
rect 17173 15921 17207 15955
rect 21037 15921 21071 15955
rect 21221 15921 21255 15955
rect 23889 15921 23923 15955
rect 24533 15921 24567 15955
rect 25821 15921 25855 15955
rect 5857 15853 5891 15887
rect 9169 15853 9203 15887
rect 9905 15853 9939 15887
rect 13125 15853 13159 15887
rect 13677 15853 13711 15887
rect 16529 15853 16563 15887
rect 20209 15853 20243 15887
rect 20761 15853 20795 15887
rect 24165 15853 24199 15887
rect 24809 15853 24843 15887
rect 2545 15785 2579 15819
rect 11929 15785 11963 15819
rect 13585 15785 13619 15819
rect 24073 15785 24107 15819
rect 2177 15717 2211 15751
rect 6685 15717 6719 15751
rect 7789 15717 7823 15751
rect 11561 15717 11595 15751
rect 15333 15717 15367 15751
rect 16069 15717 16103 15751
rect 23061 15717 23095 15751
rect 26097 15717 26131 15751
rect 1809 15513 1843 15547
rect 1901 15513 1935 15547
rect 2361 15513 2395 15547
rect 3005 15513 3039 15547
rect 4385 15513 4419 15547
rect 4937 15513 4971 15547
rect 7237 15513 7271 15547
rect 8157 15513 8191 15547
rect 9813 15513 9847 15547
rect 11377 15513 11411 15547
rect 11561 15513 11595 15547
rect 15241 15513 15275 15547
rect 16161 15513 16195 15547
rect 16897 15513 16931 15547
rect 20301 15513 20335 15547
rect 20669 15513 20703 15547
rect 24073 15513 24107 15547
rect 26281 15513 26315 15547
rect 2545 15445 2579 15479
rect 3097 15445 3131 15479
rect 7835 15445 7869 15479
rect 7973 15445 8007 15479
rect 9261 15445 9295 15479
rect 9537 15445 9571 15479
rect 14413 15445 14447 15479
rect 15609 15445 15643 15479
rect 15793 15445 15827 15479
rect 20761 15445 20795 15479
rect 2232 15377 2266 15411
rect 2453 15377 2487 15411
rect 4569 15377 4603 15411
rect 5765 15377 5799 15411
rect 5949 15377 5983 15411
rect 6133 15377 6167 15411
rect 6869 15377 6903 15411
rect 7513 15377 7547 15411
rect 8065 15377 8099 15411
rect 8525 15377 8559 15411
rect 12481 15377 12515 15411
rect 15425 15377 15459 15411
rect 20485 15377 20519 15411
rect 23613 15377 23647 15411
rect 24441 15377 24475 15411
rect 26189 15377 26223 15411
rect 26465 15377 26499 15411
rect 889 15309 923 15343
rect 1349 15309 1383 15343
rect 2085 15309 2119 15343
rect 4661 15309 4695 15343
rect 4753 15309 4787 15343
rect 5397 15309 5431 15343
rect 6409 15309 6443 15343
rect 7053 15309 7087 15343
rect 13125 15309 13159 15343
rect 14045 15309 14079 15343
rect 16069 15309 16103 15343
rect 16529 15309 16563 15343
rect 16713 15309 16747 15343
rect 22601 15309 22635 15343
rect 23245 15309 23279 15343
rect 24165 15309 24199 15343
rect 1257 15241 1291 15275
rect 1625 15241 1659 15275
rect 6493 15241 6527 15275
rect 7697 15241 7731 15275
rect 15885 15241 15919 15275
rect 5489 15173 5523 15207
rect 6317 15173 6351 15207
rect 7329 15173 7363 15207
rect 9353 15173 9387 15207
rect 9905 15173 9939 15207
rect 12665 15173 12699 15207
rect 12849 15173 12883 15207
rect 13033 15173 13067 15207
rect 22693 15173 22727 15207
rect 23245 15173 23279 15207
rect 23797 15173 23831 15207
rect 1993 14969 2027 15003
rect 4293 14969 4327 15003
rect 5949 14969 5983 15003
rect 6685 14969 6719 15003
rect 12021 14969 12055 15003
rect 12205 14969 12239 15003
rect 13217 14969 13251 15003
rect 15885 14969 15919 15003
rect 23705 14969 23739 15003
rect 24257 14969 24291 15003
rect 2453 14901 2487 14935
rect 4109 14901 4143 14935
rect 5489 14901 5523 14935
rect 6593 14901 6627 14935
rect 13309 14901 13343 14935
rect 23797 14901 23831 14935
rect 24349 14901 24383 14935
rect 24625 14901 24659 14935
rect 2177 14833 2211 14867
rect 3465 14833 3499 14867
rect 5305 14833 5339 14867
rect 5397 14833 5431 14867
rect 6409 14833 6443 14867
rect 7329 14833 7363 14867
rect 8985 14833 9019 14867
rect 9169 14833 9203 14867
rect 11377 14833 11411 14867
rect 16989 14833 17023 14867
rect 17173 14833 17207 14867
rect 18001 14833 18035 14867
rect 22785 14833 22819 14867
rect 22969 14833 23003 14867
rect 23337 14833 23371 14867
rect 3373 14765 3407 14799
rect 5121 14765 5155 14799
rect 5857 14765 5891 14799
rect 7697 14765 7731 14799
rect 11745 14765 11779 14799
rect 16161 14765 16195 14799
rect 16713 14765 16747 14799
rect 22325 14765 22359 14799
rect 23245 14765 23279 14799
rect 7605 14697 7639 14731
rect 11542 14697 11576 14731
rect 12389 14697 12423 14731
rect 2361 14629 2395 14663
rect 3649 14629 3683 14663
rect 6133 14629 6167 14663
rect 7467 14629 7501 14663
rect 7973 14629 8007 14663
rect 9261 14629 9295 14663
rect 9905 14629 9939 14663
rect 10181 14629 10215 14663
rect 11653 14629 11687 14663
rect 17817 14629 17851 14663
rect 18277 14629 18311 14663
rect 19841 14629 19875 14663
rect 1533 14425 1567 14459
rect 2269 14425 2303 14459
rect 3097 14425 3131 14459
rect 3557 14425 3591 14459
rect 3833 14425 3867 14459
rect 4090 14425 4124 14459
rect 4569 14425 4603 14459
rect 6501 14425 6535 14459
rect 6777 14425 6811 14459
rect 6961 14425 6995 14459
rect 8433 14425 8467 14459
rect 8617 14425 8651 14459
rect 9169 14425 9203 14459
rect 9353 14425 9387 14459
rect 9537 14425 9571 14459
rect 10733 14425 10767 14459
rect 12205 14425 12239 14459
rect 12941 14425 12975 14459
rect 13861 14425 13895 14459
rect 16713 14425 16747 14459
rect 17081 14425 17115 14459
rect 17449 14425 17483 14459
rect 22601 14425 22635 14459
rect 1349 14357 1383 14391
rect 1901 14357 1935 14391
rect 4201 14357 4235 14391
rect 7513 14357 7547 14391
rect 8249 14357 8283 14391
rect 9077 14357 9111 14391
rect 11883 14357 11917 14391
rect 12021 14357 12055 14391
rect 16437 14357 16471 14391
rect 16621 14357 16655 14391
rect 20577 14357 20611 14391
rect 22233 14357 22267 14391
rect 22785 14357 22819 14391
rect 2140 14289 2174 14323
rect 2361 14289 2395 14323
rect 4293 14289 4327 14323
rect 5121 14289 5155 14323
rect 7384 14289 7418 14323
rect 7605 14289 7639 14323
rect 10641 14289 10675 14323
rect 12113 14289 12147 14323
rect 12573 14289 12607 14323
rect 18461 14289 18495 14323
rect 19657 14289 19691 14323
rect 19933 14289 19967 14323
rect 22969 14289 23003 14323
rect 23521 14289 23555 14323
rect 25637 14289 25671 14323
rect 26189 14289 26223 14323
rect 5765 14221 5799 14255
rect 7145 14221 7179 14255
rect 7237 14221 7271 14255
rect 9905 14221 9939 14255
rect 10181 14221 10215 14255
rect 13585 14221 13619 14255
rect 18369 14221 18403 14255
rect 18737 14221 18771 14255
rect 18921 14221 18955 14255
rect 19473 14221 19507 14255
rect 20117 14221 20151 14255
rect 20577 14221 20611 14255
rect 22417 14221 22451 14255
rect 23797 14221 23831 14255
rect 23981 14221 24015 14255
rect 24073 14221 24107 14255
rect 25453 14221 25487 14255
rect 26005 14221 26039 14255
rect 1993 14153 2027 14187
rect 2729 14153 2763 14187
rect 3925 14153 3959 14187
rect 4753 14153 4787 14187
rect 7973 14153 8007 14187
rect 8801 14153 8835 14187
rect 10273 14153 10307 14187
rect 11101 14153 11135 14187
rect 11285 14153 11319 14187
rect 11745 14153 11779 14187
rect 12849 14153 12883 14187
rect 16253 14153 16287 14187
rect 17725 14153 17759 14187
rect 1625 14085 1659 14119
rect 2821 14085 2855 14119
rect 3281 14085 3315 14119
rect 3373 14085 3407 14119
rect 5397 14085 5431 14119
rect 5581 14085 5615 14119
rect 5949 14085 5983 14119
rect 6317 14085 6351 14119
rect 8065 14085 8099 14119
rect 9721 14085 9755 14119
rect 10089 14085 10123 14119
rect 11469 14085 11503 14119
rect 13677 14085 13711 14119
rect 14045 14085 14079 14119
rect 16989 14085 17023 14119
rect 17633 14085 17667 14119
rect 22049 14085 22083 14119
rect 4293 13881 4327 13915
rect 4753 13881 4787 13915
rect 12113 13881 12147 13915
rect 18001 13881 18035 13915
rect 19841 13881 19875 13915
rect 22325 13881 22359 13915
rect 23061 13881 23095 13915
rect 23429 13881 23463 13915
rect 23705 13881 23739 13915
rect 4017 13813 4051 13847
rect 7605 13813 7639 13847
rect 7697 13813 7731 13847
rect 9997 13813 10031 13847
rect 10181 13813 10215 13847
rect 10549 13813 10583 13847
rect 20209 13813 20243 13847
rect 1809 13745 1843 13779
rect 1993 13745 2027 13779
rect 4201 13745 4235 13779
rect 7513 13745 7547 13779
rect 10089 13745 10123 13779
rect 11377 13745 11411 13779
rect 11561 13745 11595 13779
rect 15793 13745 15827 13779
rect 18553 13745 18587 13779
rect 18700 13745 18734 13779
rect 20393 13745 20427 13779
rect 21681 13745 21715 13779
rect 23245 13745 23279 13779
rect 7329 13677 7363 13711
rect 8065 13677 8099 13711
rect 9813 13677 9847 13711
rect 12205 13677 12239 13711
rect 18921 13677 18955 13711
rect 21589 13677 21623 13711
rect 15885 13609 15919 13643
rect 18829 13609 18863 13643
rect 2085 13541 2119 13575
rect 6133 13541 6167 13575
rect 8157 13541 8191 13575
rect 9261 13541 9295 13575
rect 11653 13541 11687 13575
rect 13309 13541 13343 13575
rect 17817 13541 17851 13575
rect 19197 13541 19231 13575
rect 20485 13541 20519 13575
rect 20945 13541 20979 13575
rect 21865 13541 21899 13575
rect 1717 13337 1751 13371
rect 1901 13337 1935 13371
rect 2269 13337 2303 13371
rect 2821 13337 2855 13371
rect 3281 13337 3315 13371
rect 3557 13337 3591 13371
rect 5121 13337 5155 13371
rect 5581 13337 5615 13371
rect 7421 13337 7455 13371
rect 7973 13337 8007 13371
rect 8157 13337 8191 13371
rect 10089 13337 10123 13371
rect 10549 13337 10583 13371
rect 11377 13337 11411 13371
rect 15793 13337 15827 13371
rect 15977 13337 16011 13371
rect 17817 13337 17851 13371
rect 18553 13337 18587 13371
rect 18737 13337 18771 13371
rect 18921 13337 18955 13371
rect 19197 13337 19231 13371
rect 20025 13337 20059 13371
rect 21957 13337 21991 13371
rect 22141 13337 22175 13371
rect 23153 13337 23187 13371
rect 24073 13337 24107 13371
rect 24441 13337 24475 13371
rect 3649 13269 3683 13303
rect 6961 13269 6995 13303
rect 7145 13269 7179 13303
rect 9353 13269 9387 13303
rect 11193 13269 11227 13303
rect 12941 13269 12975 13303
rect 19749 13269 19783 13303
rect 20393 13269 20427 13303
rect 4109 13201 4143 13235
rect 4201 13201 4235 13235
rect 4937 13201 4971 13235
rect 7605 13201 7639 13235
rect 8065 13201 8099 13235
rect 8525 13201 8559 13235
rect 11009 13201 11043 13235
rect 13401 13201 13435 13235
rect 14229 13201 14263 13235
rect 21221 13201 21255 13235
rect 22325 13201 22359 13235
rect 23061 13201 23095 13235
rect 23613 13201 23647 13235
rect 1993 13133 2027 13167
rect 2177 13133 2211 13167
rect 4477 13133 4511 13167
rect 5673 13133 5707 13167
rect 5949 13133 5983 13167
rect 7697 13133 7731 13167
rect 7844 13133 7878 13167
rect 9261 13133 9295 13167
rect 9537 13133 9571 13167
rect 10641 13133 10675 13167
rect 11929 13133 11963 13167
rect 12389 13133 12423 13167
rect 13309 13133 13343 13167
rect 14137 13133 14171 13167
rect 17633 13133 17667 13167
rect 19289 13133 19323 13167
rect 20209 13133 20243 13167
rect 21313 13133 21347 13167
rect 21681 13133 21715 13167
rect 21865 13133 21899 13167
rect 23981 13133 24015 13167
rect 25453 13133 25487 13167
rect 2637 13065 2671 13099
rect 4385 13065 4419 13099
rect 4569 13065 4603 13099
rect 6133 13065 6167 13099
rect 6501 13065 6535 13099
rect 6869 13065 6903 13099
rect 9169 13065 9203 13099
rect 11745 13065 11779 13099
rect 12297 13065 12331 13099
rect 13125 13065 13159 13099
rect 17725 13065 17759 13099
rect 18001 13065 18035 13099
rect 20669 13065 20703 13099
rect 23797 13065 23831 13099
rect 24717 13065 24751 13099
rect 25545 13065 25579 13099
rect 25637 13065 25671 13099
rect 1349 12997 1383 13031
rect 1533 12997 1567 13031
rect 3925 12997 3959 13031
rect 6317 12997 6351 13031
rect 6409 12997 6443 13031
rect 8893 12997 8927 13031
rect 9721 12997 9755 13031
rect 10365 12997 10399 13031
rect 12573 12997 12607 13031
rect 20577 12997 20611 13031
rect 25821 12997 25855 13031
rect 1901 12793 1935 12827
rect 8065 12793 8099 12827
rect 9261 12793 9295 12827
rect 12205 12793 12239 12827
rect 13309 12793 13343 12827
rect 20485 12793 20519 12827
rect 20853 12793 20887 12827
rect 4201 12725 4235 12759
rect 5857 12725 5891 12759
rect 7605 12725 7639 12759
rect 17449 12725 17483 12759
rect 1625 12657 1659 12691
rect 1809 12657 1843 12691
rect 4385 12657 4419 12691
rect 5949 12657 5983 12691
rect 7789 12657 7823 12691
rect 11009 12657 11043 12691
rect 11469 12657 11503 12691
rect 11837 12657 11871 12691
rect 15241 12657 15275 12691
rect 17633 12657 17667 12691
rect 20485 12657 20519 12691
rect 21681 12657 21715 12691
rect 21865 12657 21899 12691
rect 23429 12657 23463 12691
rect 23705 12657 23739 12691
rect 24073 12657 24107 12691
rect 4753 12589 4787 12623
rect 6317 12589 6351 12623
rect 7881 12589 7915 12623
rect 8249 12589 8283 12623
rect 9813 12589 9847 12623
rect 11929 12589 11963 12623
rect 15425 12589 15459 12623
rect 20761 12589 20795 12623
rect 21957 12589 21991 12623
rect 23981 12589 24015 12623
rect 3741 12521 3775 12555
rect 6225 12521 6259 12555
rect 6777 12521 6811 12555
rect 23521 12521 23555 12555
rect 2269 12453 2303 12487
rect 4109 12453 4143 12487
rect 6114 12453 6148 12487
rect 6593 12453 6627 12487
rect 7421 12453 7455 12487
rect 14321 12453 14355 12487
rect 17725 12453 17759 12487
rect 1257 12249 1291 12283
rect 1901 12249 1935 12283
rect 5857 12249 5891 12283
rect 6409 12249 6443 12283
rect 6593 12249 6627 12283
rect 7145 12249 7179 12283
rect 7513 12249 7547 12283
rect 11469 12249 11503 12283
rect 17633 12249 17667 12283
rect 17817 12249 17851 12283
rect 20301 12249 20335 12283
rect 21865 12249 21899 12283
rect 22785 12249 22819 12283
rect 23337 12249 23371 12283
rect 23521 12249 23555 12283
rect 1533 12181 1567 12215
rect 2361 12181 2395 12215
rect 4569 12181 4603 12215
rect 5121 12181 5155 12215
rect 5581 12181 5615 12215
rect 6271 12181 6305 12215
rect 7053 12181 7087 12215
rect 11745 12181 11779 12215
rect 17541 12181 17575 12215
rect 20485 12181 20519 12215
rect 22601 12181 22635 12215
rect 2232 12113 2266 12147
rect 2453 12113 2487 12147
rect 3465 12113 3499 12147
rect 4385 12113 4419 12147
rect 5765 12113 5799 12147
rect 6501 12113 6535 12147
rect 14321 12113 14355 12147
rect 21681 12113 21715 12147
rect 23153 12113 23187 12147
rect 23981 12113 24015 12147
rect 2085 12045 2119 12079
rect 2913 12045 2947 12079
rect 7329 12045 7363 12079
rect 7973 12045 8007 12079
rect 23705 12045 23739 12079
rect 3373 11977 3407 12011
rect 4017 11977 4051 12011
rect 5397 11977 5431 12011
rect 6133 11977 6167 12011
rect 8065 11977 8099 12011
rect 8249 11977 8283 12011
rect 8433 11977 8467 12011
rect 8801 11977 8835 12011
rect 14229 11977 14263 12011
rect 14597 11977 14631 12011
rect 16345 11977 16379 12011
rect 21497 11977 21531 12011
rect 25729 11977 25763 12011
rect 1625 11909 1659 11943
rect 2729 11909 2763 11943
rect 3833 11909 3867 11943
rect 3925 11909 3959 11943
rect 4661 11909 4695 11943
rect 4937 11909 4971 11943
rect 7697 11909 7731 11943
rect 8341 11909 8375 11943
rect 8893 11909 8927 11943
rect 11009 11909 11043 11943
rect 11285 11909 11319 11943
rect 14045 11909 14079 11943
rect 2269 11705 2303 11739
rect 3925 11705 3959 11739
rect 4477 11705 4511 11739
rect 9445 11705 9479 11739
rect 10825 11705 10859 11739
rect 15425 11705 15459 11739
rect 23153 11705 23187 11739
rect 24165 11705 24199 11739
rect 1533 11637 1567 11671
rect 3649 11637 3683 11671
rect 4385 11637 4419 11671
rect 5949 11637 5983 11671
rect 7329 11637 7363 11671
rect 9537 11637 9571 11671
rect 14413 11637 14447 11671
rect 23797 11637 23831 11671
rect 24717 11637 24751 11671
rect 1717 11569 1751 11603
rect 4553 11569 4587 11603
rect 6777 11569 6811 11603
rect 9353 11569 9387 11603
rect 10733 11569 10767 11603
rect 12849 11569 12883 11603
rect 15333 11569 15367 11603
rect 23889 11569 23923 11603
rect 24441 11569 24475 11603
rect 4201 11501 4235 11535
rect 4937 11501 4971 11535
rect 6501 11501 6535 11535
rect 6961 11501 6995 11535
rect 9169 11501 9203 11535
rect 9905 11501 9939 11535
rect 14597 11433 14631 11467
rect 1809 11365 1843 11399
rect 2361 11365 2395 11399
rect 8065 11365 8099 11399
rect 13033 11365 13067 11399
rect 13217 11365 13251 11399
rect 13401 11365 13435 11399
rect 1625 11161 1659 11195
rect 1809 11161 1843 11195
rect 2361 11161 2395 11195
rect 3373 11161 3407 11195
rect 3833 11161 3867 11195
rect 4385 11161 4419 11195
rect 4753 11161 4787 11195
rect 6501 11161 6535 11195
rect 6685 11161 6719 11195
rect 9997 11161 10031 11195
rect 10825 11161 10859 11195
rect 13953 11161 13987 11195
rect 14670 11161 14704 11195
rect 15333 11161 15367 11195
rect 24441 11161 24475 11195
rect 24717 11161 24751 11195
rect 4201 11093 4235 11127
rect 6133 11093 6167 11127
rect 6409 11093 6443 11127
rect 7605 11093 7639 11127
rect 13861 11093 13895 11127
rect 14781 11093 14815 11127
rect 18185 11093 18219 11127
rect 18553 11093 18587 11127
rect 2821 11025 2855 11059
rect 3649 11025 3683 11059
rect 4293 11025 4327 11059
rect 9721 11025 9755 11059
rect 10917 11025 10951 11059
rect 12297 11025 12331 11059
rect 12665 11025 12699 11059
rect 12849 11025 12883 11059
rect 13677 11025 13711 11059
rect 14413 11025 14447 11059
rect 14873 11025 14907 11059
rect 21681 11025 21715 11059
rect 2269 10957 2303 10991
rect 3281 10957 3315 10991
rect 4072 10957 4106 10991
rect 4937 10957 4971 10991
rect 7053 10957 7087 10991
rect 7789 10957 7823 10991
rect 7973 10957 8007 10991
rect 8157 10957 8191 10991
rect 9169 10957 9203 10991
rect 9629 10957 9663 10991
rect 11929 10957 11963 10991
rect 12389 10957 12423 10991
rect 13125 10957 13159 10991
rect 13309 10957 13343 10991
rect 18369 10957 18403 10991
rect 18737 10957 18771 10991
rect 19197 10957 19231 10991
rect 19289 10957 19323 10991
rect 21129 10957 21163 10991
rect 1901 10889 1935 10923
rect 2085 10889 2119 10923
rect 3925 10889 3959 10923
rect 9353 10889 9387 10923
rect 11561 10889 11595 10923
rect 11745 10889 11779 10923
rect 14229 10889 14263 10923
rect 14505 10889 14539 10923
rect 21405 10889 21439 10923
rect 21865 10889 21899 10923
rect 3005 10821 3039 10855
rect 5213 10821 5247 10855
rect 7237 10821 7271 10855
rect 12941 10821 12975 10855
rect 15149 10821 15183 10855
rect 1809 10617 1843 10651
rect 2177 10617 2211 10651
rect 4569 10617 4603 10651
rect 7421 10617 7455 10651
rect 19289 10617 19323 10651
rect 23153 10617 23187 10651
rect 23797 10617 23831 10651
rect 4385 10549 4419 10583
rect 5673 10549 5707 10583
rect 8985 10549 9019 10583
rect 9169 10549 9203 10583
rect 9353 10549 9387 10583
rect 9721 10549 9755 10583
rect 3741 10481 3775 10515
rect 3925 10481 3959 10515
rect 4293 10481 4327 10515
rect 5121 10481 5155 10515
rect 5305 10481 5339 10515
rect 9261 10481 9295 10515
rect 12297 10481 12331 10515
rect 12757 10481 12791 10515
rect 13125 10481 13159 10515
rect 15241 10481 15275 10515
rect 15609 10481 15643 10515
rect 15701 10481 15735 10515
rect 17817 10481 17851 10515
rect 18001 10481 18035 10515
rect 18369 10481 18403 10515
rect 18553 10481 18587 10515
rect 20209 10481 20243 10515
rect 23337 10481 23371 10515
rect 24441 10481 24475 10515
rect 8617 10413 8651 10447
rect 15333 10413 15367 10447
rect 20485 10413 20519 10447
rect 22233 10413 22267 10447
rect 24717 10413 24751 10447
rect 13125 10345 13159 10379
rect 19473 10345 19507 10379
rect 14413 10277 14447 10311
rect 14689 10277 14723 10311
rect 17633 10277 17667 10311
rect 19105 10277 19139 10311
rect 24073 10277 24107 10311
rect 1441 10073 1475 10107
rect 1855 10073 1889 10107
rect 2637 10073 2671 10107
rect 3005 10073 3039 10107
rect 3189 10073 3223 10107
rect 4201 10073 4235 10107
rect 4569 10073 4603 10107
rect 5213 10073 5247 10107
rect 5581 10073 5615 10107
rect 6777 10073 6811 10107
rect 7237 10073 7271 10107
rect 8157 10073 8191 10107
rect 9813 10073 9847 10107
rect 11469 10073 11503 10107
rect 11837 10073 11871 10107
rect 12665 10073 12699 10107
rect 13125 10073 13159 10107
rect 13861 10073 13895 10107
rect 14413 10073 14447 10107
rect 16989 10073 17023 10107
rect 19013 10073 19047 10107
rect 20669 10073 20703 10107
rect 20945 10073 20979 10107
rect 23245 10073 23279 10107
rect 23521 10073 23555 10107
rect 1625 10005 1659 10039
rect 1993 10005 2027 10039
rect 7881 10005 7915 10039
rect 9629 10005 9663 10039
rect 14045 10005 14079 10039
rect 17173 10005 17207 10039
rect 17909 10005 17943 10039
rect 18461 10005 18495 10039
rect 2085 9937 2119 9971
rect 4293 9937 4327 9971
rect 7605 9937 7639 9971
rect 12297 9937 12331 9971
rect 14505 9937 14539 9971
rect 16069 9937 16103 9971
rect 16253 9937 16287 9971
rect 18645 9937 18679 9971
rect 19105 9937 19139 9971
rect 20393 9937 20427 9971
rect 25821 9937 25855 9971
rect 3465 9869 3499 9903
rect 3649 9869 3683 9903
rect 6961 9869 6995 9903
rect 7053 9869 7087 9903
rect 8801 9869 8835 9903
rect 9997 9869 10031 9903
rect 10181 9869 10215 9903
rect 12021 9869 12055 9903
rect 12481 9869 12515 9903
rect 14965 9869 14999 9903
rect 15149 9869 15183 9903
rect 15333 9869 15367 9903
rect 15609 9869 15643 9903
rect 15977 9869 16011 9903
rect 17725 9869 17759 9903
rect 17817 9869 17851 9903
rect 1717 9801 1751 9835
rect 4017 9801 4051 9835
rect 5305 9801 5339 9835
rect 8617 9801 8651 9835
rect 8985 9801 9019 9835
rect 9353 9801 9387 9835
rect 12941 9801 12975 9835
rect 19565 9869 19599 9903
rect 19749 9869 19783 9903
rect 20025 9869 20059 9903
rect 20577 9869 20611 9903
rect 21129 9869 21163 9903
rect 23797 9869 23831 9903
rect 24073 9801 24107 9835
rect 2361 9733 2395 9767
rect 3373 9733 3407 9767
rect 8249 9733 8283 9767
rect 8525 9733 8559 9767
rect 8893 9733 8927 9767
rect 9445 9733 9479 9767
rect 13585 9733 13619 9767
rect 14137 9733 14171 9767
rect 17357 9733 17391 9767
rect 17541 9733 17575 9767
rect 17725 9733 17759 9767
rect 18277 9733 18311 9767
rect 18645 9733 18679 9767
rect 18829 9733 18863 9767
rect 23061 9733 23095 9767
rect 23613 9733 23647 9767
rect 705 9529 739 9563
rect 981 9529 1015 9563
rect 1809 9529 1843 9563
rect 8617 9529 8651 9563
rect 12573 9529 12607 9563
rect 15425 9529 15459 9563
rect 17449 9529 17483 9563
rect 19473 9529 19507 9563
rect 20301 9529 20335 9563
rect 24533 9529 24567 9563
rect 24717 9529 24751 9563
rect 1901 9461 1935 9495
rect 6133 9461 6167 9495
rect 14413 9461 14447 9495
rect 19289 9461 19323 9495
rect 2085 9393 2119 9427
rect 3833 9393 3867 9427
rect 4293 9393 4327 9427
rect 4569 9393 4603 9427
rect 4753 9393 4787 9427
rect 6685 9393 6719 9427
rect 6961 9393 6995 9427
rect 9077 9393 9111 9427
rect 11193 9393 11227 9427
rect 12481 9393 12515 9427
rect 14689 9393 14723 9427
rect 16621 9393 16655 9427
rect 18737 9393 18771 9427
rect 18921 9393 18955 9427
rect 23429 9393 23463 9427
rect 23705 9393 23739 9427
rect 24165 9393 24199 9427
rect 2453 9325 2487 9359
rect 5121 9325 5155 9359
rect 5213 9325 5247 9359
rect 7145 9325 7179 9359
rect 8985 9325 9019 9359
rect 11101 9325 11135 9359
rect 14597 9325 14631 9359
rect 24349 9325 24383 9359
rect 16437 9257 16471 9291
rect 23429 9257 23463 9291
rect 9261 9189 9295 9223
rect 11377 9189 11411 9223
rect 14873 9189 14907 9223
rect 15241 9189 15275 9223
rect 2085 8985 2119 9019
rect 3005 8985 3039 9019
rect 3189 8985 3223 9019
rect 3557 8985 3591 9019
rect 4293 8985 4327 9019
rect 4937 8985 4971 9019
rect 5581 8985 5615 9019
rect 7605 8985 7639 9019
rect 8065 8985 8099 9019
rect 9077 8985 9111 9019
rect 9261 8985 9295 9019
rect 9353 8985 9387 9019
rect 11193 8985 11227 9019
rect 12297 8985 12331 9019
rect 12389 8985 12423 9019
rect 15333 8985 15367 9019
rect 16437 8985 16471 9019
rect 16529 8985 16563 9019
rect 19105 8985 19139 9019
rect 19289 8985 19323 9019
rect 21129 8985 21163 9019
rect 21681 8985 21715 9019
rect 22233 8985 22267 9019
rect 22601 8985 22635 9019
rect 22785 8985 22819 9019
rect 23061 8985 23095 9019
rect 23429 8985 23463 9019
rect 24165 8985 24199 9019
rect 24349 8985 24383 9019
rect 25453 8985 25487 9019
rect 1993 8917 2027 8951
rect 3281 8917 3315 8951
rect 3741 8917 3775 8951
rect 5765 8917 5799 8951
rect 11837 8917 11871 8951
rect 13401 8917 13435 8951
rect 14229 8917 14263 8951
rect 17817 8917 17851 8951
rect 18921 8917 18955 8951
rect 23318 8917 23352 8951
rect 1717 8849 1751 8883
rect 3925 8849 3959 8883
rect 6961 8849 6995 8883
rect 8617 8849 8651 8883
rect 11469 8849 11503 8883
rect 12665 8849 12699 8883
rect 14965 8849 14999 8883
rect 23521 8849 23555 8883
rect 23889 8849 23923 8883
rect 24533 8849 24567 8883
rect 25177 8849 25211 8883
rect 25269 8849 25303 8883
rect 797 8781 831 8815
rect 1625 8781 1659 8815
rect 4017 8781 4051 8815
rect 4109 8781 4143 8815
rect 5949 8781 5983 8815
rect 7789 8781 7823 8815
rect 7881 8781 7915 8815
rect 11285 8781 11319 8815
rect 13125 8781 13159 8815
rect 13401 8781 13435 8815
rect 14689 8781 14723 8815
rect 15149 8781 15183 8815
rect 17909 8781 17943 8815
rect 18093 8781 18127 8815
rect 18461 8781 18495 8815
rect 21313 8781 21347 8815
rect 22417 8781 22451 8815
rect 23153 8781 23187 8815
rect 23981 8781 24015 8815
rect 25085 8781 25119 8815
rect 889 8713 923 8747
rect 6133 8713 6167 8747
rect 6501 8713 6535 8747
rect 6869 8713 6903 8747
rect 8525 8713 8559 8747
rect 12113 8713 12147 8747
rect 13953 8713 13987 8747
rect 14413 8713 14447 8747
rect 14505 8713 14539 8747
rect 18737 8713 18771 8747
rect 2361 8645 2395 8679
rect 4753 8645 4787 8679
rect 5397 8645 5431 8679
rect 6317 8645 6351 8679
rect 6409 8645 6443 8679
rect 7145 8645 7179 8679
rect 18553 8645 18587 8679
rect 21589 8645 21623 8679
rect 705 8441 739 8475
rect 889 8441 923 8475
rect 3833 8441 3867 8475
rect 6225 8441 6259 8475
rect 9077 8441 9111 8475
rect 12849 8441 12883 8475
rect 14689 8441 14723 8475
rect 23153 8441 23187 8475
rect 4109 8373 4143 8407
rect 6409 8373 6443 8407
rect 6685 8373 6719 8407
rect 11285 8373 11319 8407
rect 11837 8373 11871 8407
rect 1441 8305 1475 8339
rect 1625 8305 1659 8339
rect 4293 8305 4327 8339
rect 4661 8305 4695 8339
rect 5765 8305 5799 8339
rect 8985 8305 9019 8339
rect 11469 8305 11503 8339
rect 15241 8305 15275 8339
rect 15425 8305 15459 8339
rect 15609 8305 15643 8339
rect 17725 8305 17759 8339
rect 18277 8305 18311 8339
rect 23613 8305 23647 8339
rect 24257 8305 24291 8339
rect 26097 8305 26131 8339
rect 14781 8237 14815 8271
rect 23521 8237 23555 8271
rect 23981 8237 24015 8271
rect 24533 8237 24567 8271
rect 12665 8169 12699 8203
rect 1717 8101 1751 8135
rect 6041 8101 6075 8135
rect 12481 8101 12515 8135
rect 17817 8101 17851 8135
rect 18553 8101 18587 8135
rect 18829 8101 18863 8135
rect 26097 8101 26131 8135
rect 1625 7897 1659 7931
rect 1809 7897 1843 7931
rect 4201 7897 4235 7931
rect 4385 7897 4419 7931
rect 4569 7897 4603 7931
rect 5765 7897 5799 7931
rect 6133 7897 6167 7931
rect 9077 7897 9111 7931
rect 11377 7897 11411 7931
rect 11837 7897 11871 7931
rect 12205 7897 12239 7931
rect 15241 7897 15275 7931
rect 16989 7897 17023 7931
rect 20577 7897 20611 7931
rect 20945 7897 20979 7931
rect 21497 7897 21531 7931
rect 23153 7897 23187 7931
rect 23705 7897 23739 7931
rect 23981 7897 24015 7931
rect 26281 7897 26315 7931
rect 9169 7829 9203 7863
rect 12113 7829 12147 7863
rect 14413 7829 14447 7863
rect 15057 7829 15091 7863
rect 23337 7829 23371 7863
rect 1533 7761 1567 7795
rect 12941 7761 12975 7795
rect 19105 7761 19139 7795
rect 20669 7761 20703 7795
rect 21313 7761 21347 7795
rect 24441 7761 24475 7795
rect 13033 7693 13067 7727
rect 13401 7693 13435 7727
rect 13585 7693 13619 7727
rect 14413 7693 14447 7727
rect 15701 7693 15735 7727
rect 15885 7693 15919 7727
rect 17173 7693 17207 7727
rect 18461 7693 18495 7727
rect 18645 7693 18679 7727
rect 18921 7693 18955 7727
rect 19473 7693 19507 7727
rect 20761 7693 20795 7727
rect 24165 7693 24199 7727
rect 12389 7625 12423 7659
rect 14597 7625 14631 7659
rect 15793 7625 15827 7659
rect 16069 7625 16103 7659
rect 17909 7625 17943 7659
rect 18001 7625 18035 7659
rect 26189 7625 26223 7659
rect 26465 7625 26499 7659
rect 11469 7557 11503 7591
rect 14873 7557 14907 7591
rect 17541 7557 17575 7591
rect 17725 7557 17759 7591
rect 23521 7557 23555 7591
rect 23889 7557 23923 7591
rect 12481 7353 12515 7387
rect 17725 7353 17759 7387
rect 18093 7353 18127 7387
rect 20945 7353 20979 7387
rect 24349 7353 24383 7387
rect 24625 7353 24659 7387
rect 12573 7285 12607 7319
rect 24257 7285 24291 7319
rect 1625 7217 1659 7251
rect 6317 7217 6351 7251
rect 6501 7217 6535 7251
rect 6685 7217 6719 7251
rect 9445 7217 9479 7251
rect 9629 7217 9663 7251
rect 9905 7217 9939 7251
rect 11285 7217 11319 7251
rect 12849 7217 12883 7251
rect 15609 7217 15643 7251
rect 15977 7217 16011 7251
rect 16161 7217 16195 7251
rect 18829 7217 18863 7251
rect 19105 7217 19139 7251
rect 20301 7217 20335 7251
rect 21589 7217 21623 7251
rect 2177 7149 2211 7183
rect 8985 7149 9019 7183
rect 10089 7149 10123 7183
rect 10365 7149 10399 7183
rect 12757 7149 12791 7183
rect 15701 7149 15735 7183
rect 18277 7149 18311 7183
rect 19289 7149 19323 7183
rect 20209 7149 20243 7183
rect 1533 7081 1567 7115
rect 2085 7081 2119 7115
rect 6133 7081 6167 7115
rect 11377 7013 11411 7047
rect 13033 7013 13067 7047
rect 15057 7013 15091 7047
rect 20485 7013 20519 7047
rect 21129 7013 21163 7047
rect 21681 7013 21715 7047
rect 981 6809 1015 6843
rect 1349 6809 1383 6843
rect 2453 6809 2487 6843
rect 6133 6809 6167 6843
rect 6593 6809 6627 6843
rect 8617 6809 8651 6843
rect 8893 6809 8927 6843
rect 9261 6809 9295 6843
rect 9537 6809 9571 6843
rect 10457 6809 10491 6843
rect 13125 6809 13159 6843
rect 14597 6809 14631 6843
rect 19105 6809 19139 6843
rect 19933 6809 19967 6843
rect 22049 6809 22083 6843
rect 5949 6741 5983 6775
rect 9445 6741 9479 6775
rect 11469 6741 11503 6775
rect 14781 6741 14815 6775
rect 20485 6741 20519 6775
rect 20945 6741 20979 6775
rect 9077 6673 9111 6707
rect 14413 6673 14447 6707
rect 15517 6673 15551 6707
rect 16161 6673 16195 6707
rect 21497 6673 21531 6707
rect 25361 6673 25395 6707
rect 25913 6673 25947 6707
rect 1441 6605 1475 6639
rect 2085 6605 2119 6639
rect 3189 6605 3223 6639
rect 3465 6605 3499 6639
rect 7053 6605 7087 6639
rect 7329 6605 7363 6639
rect 9905 6605 9939 6639
rect 10733 6605 10767 6639
rect 13033 6605 13067 6639
rect 15057 6605 15091 6639
rect 15149 6605 15183 6639
rect 15333 6605 15367 6639
rect 17725 6605 17759 6639
rect 18001 6605 18035 6639
rect 18093 6605 18127 6639
rect 18277 6605 18311 6639
rect 18829 6605 18863 6639
rect 20945 6605 20979 6639
rect 21221 6605 21255 6639
rect 21681 6605 21715 6639
rect 22233 6605 22267 6639
rect 24257 6605 24291 6639
rect 25177 6605 25211 6639
rect 25729 6605 25763 6639
rect 1165 6537 1199 6571
rect 2361 6537 2395 6571
rect 3373 6537 3407 6571
rect 3649 6537 3683 6571
rect 6409 6537 6443 6571
rect 9721 6537 9755 6571
rect 10273 6537 10307 6571
rect 10549 6537 10583 6571
rect 14873 6537 14907 6571
rect 17173 6537 17207 6571
rect 17909 6537 17943 6571
rect 20117 6537 20151 6571
rect 20301 6537 20335 6571
rect 24349 6537 24383 6571
rect 24441 6537 24475 6571
rect 6869 6469 6903 6503
rect 7145 6469 7179 6503
rect 11377 6469 11411 6503
rect 12757 6469 12791 6503
rect 14229 6469 14263 6503
rect 15885 6469 15919 6503
rect 17449 6469 17483 6503
rect 18461 6469 18495 6503
rect 19657 6469 19691 6503
rect 24625 6469 24659 6503
rect 1993 6265 2027 6299
rect 3373 6265 3407 6299
rect 10365 6265 10399 6299
rect 11929 6265 11963 6299
rect 15425 6265 15459 6299
rect 18553 6265 18587 6299
rect 20945 6265 20979 6299
rect 797 6129 831 6163
rect 1625 6129 1659 6163
rect 1717 6129 1751 6163
rect 3557 6129 3591 6163
rect 5305 6129 5339 6163
rect 6409 6129 6443 6163
rect 7145 6129 7179 6163
rect 7329 6129 7363 6163
rect 9537 6129 9571 6163
rect 10281 6129 10315 6163
rect 14597 6197 14631 6231
rect 15241 6197 15275 6231
rect 18645 6197 18679 6231
rect 20209 6197 20243 6231
rect 14781 6129 14815 6163
rect 16069 6129 16103 6163
rect 17633 6129 17667 6163
rect 20393 6129 20427 6163
rect 22141 6129 22175 6163
rect 24257 6129 24291 6163
rect 24441 6129 24475 6163
rect 889 6061 923 6095
rect 4845 6061 4879 6095
rect 5397 6061 5431 6095
rect 9445 6061 9479 6095
rect 15149 6061 15183 6095
rect 15977 6061 16011 6095
rect 17780 6061 17814 6095
rect 18001 6061 18035 6095
rect 24165 6061 24199 6095
rect 11837 5993 11871 6027
rect 18093 5993 18127 6027
rect 23981 5993 24015 6027
rect 4201 5925 4235 5959
rect 8709 5925 8743 5959
rect 16253 5925 16287 5959
rect 17909 5925 17943 5959
rect 20485 5925 20519 5959
rect 22141 5925 22175 5959
rect 24533 5925 24567 5959
rect 889 5721 923 5755
rect 1165 5721 1199 5755
rect 3465 5721 3499 5755
rect 5305 5721 5339 5755
rect 5489 5721 5523 5755
rect 5673 5721 5707 5755
rect 5949 5721 5983 5755
rect 6409 5721 6443 5755
rect 6593 5721 6627 5755
rect 7421 5721 7455 5755
rect 15977 5721 16011 5755
rect 16161 5721 16195 5755
rect 16345 5721 16379 5755
rect 17633 5721 17667 5755
rect 17909 5721 17943 5755
rect 20301 5721 20335 5755
rect 20485 5721 20519 5755
rect 22325 5721 22359 5755
rect 23429 5721 23463 5755
rect 23613 5721 23647 5755
rect 797 5653 831 5687
rect 3925 5653 3959 5687
rect 6317 5653 6351 5687
rect 7145 5653 7179 5687
rect 14229 5653 14263 5687
rect 23797 5653 23831 5687
rect 2361 5585 2395 5619
rect 3005 5585 3039 5619
rect 3833 5585 3867 5619
rect 6593 5585 6627 5619
rect 6685 5585 6719 5619
rect 7237 5585 7271 5619
rect 7513 5585 7547 5619
rect 8617 5585 8651 5619
rect 10733 5585 10767 5619
rect 11193 5585 11227 5619
rect 13861 5585 13895 5619
rect 18277 5585 18311 5619
rect 20025 5585 20059 5619
rect 20577 5585 20611 5619
rect 23889 5585 23923 5619
rect 24165 5585 24199 5619
rect 25913 5585 25947 5619
rect 2453 5517 2487 5551
rect 2913 5517 2947 5551
rect 4201 5517 4235 5551
rect 5029 5517 5063 5551
rect 5121 5517 5155 5551
rect 8709 5517 8743 5551
rect 11377 5517 11411 5551
rect 12205 5517 12239 5551
rect 12389 5517 12423 5551
rect 12757 5517 12791 5551
rect 12849 5517 12883 5551
rect 14045 5517 14079 5551
rect 14965 5517 14999 5551
rect 15149 5517 15183 5551
rect 15517 5517 15551 5551
rect 15609 5517 15643 5551
rect 17449 5517 17483 5551
rect 18001 5517 18035 5551
rect 21589 5517 21623 5551
rect 3097 5449 3131 5483
rect 3373 5449 3407 5483
rect 4293 5449 4327 5483
rect 8433 5449 8467 5483
rect 8985 5449 9019 5483
rect 11561 5449 11595 5483
rect 11745 5449 11779 5483
rect 14413 5449 14447 5483
rect 14505 5449 14539 5483
rect 15793 5449 15827 5483
rect 17081 5449 17115 5483
rect 21865 5449 21899 5483
rect 22233 5449 22267 5483
rect 1257 5381 1291 5415
rect 13677 5381 13711 5415
rect 21405 5381 21439 5415
rect 22509 5381 22543 5415
rect 3373 5177 3407 5211
rect 4201 5177 4235 5211
rect 6501 5177 6535 5211
rect 6777 5177 6811 5211
rect 8709 5177 8743 5211
rect 9629 5177 9663 5211
rect 9997 5177 10031 5211
rect 10273 5177 10307 5211
rect 15057 5177 15091 5211
rect 15241 5177 15275 5211
rect 17909 5177 17943 5211
rect 18369 5177 18403 5211
rect 23889 5177 23923 5211
rect 24257 5177 24291 5211
rect 6869 5109 6903 5143
rect 9353 5109 9387 5143
rect 9905 5109 9939 5143
rect 11193 5109 11227 5143
rect 12941 5109 12975 5143
rect 14965 5109 14999 5143
rect 17725 5109 17759 5143
rect 19105 5109 19139 5143
rect 21313 5109 21347 5143
rect 24717 5109 24751 5143
rect 4385 5041 4419 5075
rect 5857 5041 5891 5075
rect 9077 5041 9111 5075
rect 14873 5041 14907 5075
rect 15885 5041 15919 5075
rect 18737 5041 18771 5075
rect 24441 5041 24475 5075
rect 10917 4973 10951 5007
rect 15793 4973 15827 5007
rect 18277 4973 18311 5007
rect 21037 4973 21071 5007
rect 23061 4973 23095 5007
rect 5673 4905 5707 4939
rect 18093 4905 18127 4939
rect 2453 4837 2487 4871
rect 16069 4837 16103 4871
rect 2177 4633 2211 4667
rect 4477 4633 4511 4667
rect 4845 4633 4879 4667
rect 6777 4633 6811 4667
rect 6961 4633 6995 4667
rect 9353 4633 9387 4667
rect 11009 4633 11043 4667
rect 13217 4633 13251 4667
rect 13769 4633 13803 4667
rect 14873 4633 14907 4667
rect 15977 4633 16011 4667
rect 16161 4633 16195 4667
rect 18737 4633 18771 4667
rect 19933 4633 19967 4667
rect 21313 4633 21347 4667
rect 21681 4633 21715 4667
rect 24441 4633 24475 4667
rect 24625 4633 24659 4667
rect 11561 4565 11595 4599
rect 14689 4565 14723 4599
rect 18921 4565 18955 4599
rect 19841 4565 19875 4599
rect 21497 4565 21531 4599
rect 4569 4497 4603 4531
rect 11193 4497 11227 4531
rect 12021 4497 12055 4531
rect 12573 4497 12607 4531
rect 15885 4497 15919 4531
rect 19381 4497 19415 4531
rect 21129 4497 21163 4531
rect 2453 4429 2487 4463
rect 3925 4429 3959 4463
rect 11745 4429 11779 4463
rect 11837 4429 11871 4463
rect 13125 4429 13159 4463
rect 13585 4429 13619 4463
rect 19197 4429 19231 4463
rect 2361 4361 2395 4395
rect 4017 4361 4051 4395
rect 11377 4361 11411 4395
rect 9077 4293 9111 4327
rect 11745 4293 11779 4327
rect 12389 4293 12423 4327
rect 23705 4089 23739 4123
rect 2269 4021 2303 4055
rect 3373 4021 3407 4055
rect 15517 4021 15551 4055
rect 22601 4021 22635 4055
rect 705 3953 739 3987
rect 1625 3953 1659 3987
rect 3557 3953 3591 3987
rect 9169 3953 9203 3987
rect 22785 3953 22819 3987
rect 15241 3885 15275 3919
rect 17265 3885 17299 3919
rect 3741 3817 3775 3851
rect 9169 3749 9203 3783
rect 22877 3749 22911 3783
rect 23889 3749 23923 3783
rect 24073 3749 24107 3783
rect 797 3545 831 3579
rect 3557 3545 3591 3579
rect 3833 3545 3867 3579
rect 4569 3545 4603 3579
rect 8433 3545 8467 3579
rect 8617 3545 8651 3579
rect 15241 3545 15275 3579
rect 15885 3545 15919 3579
rect 21037 3545 21071 3579
rect 22509 3545 22543 3579
rect 22969 3545 23003 3579
rect 25315 3545 25349 3579
rect 1349 3477 1383 3511
rect 4937 3477 4971 3511
rect 15517 3477 15551 3511
rect 889 3409 923 3443
rect 1533 3409 1567 3443
rect 5673 3409 5707 3443
rect 17541 3409 17575 3443
rect 18093 3409 18127 3443
rect 4201 3341 4235 3375
rect 4569 3341 4603 3375
rect 6133 3341 6167 3375
rect 6593 3341 6627 3375
rect 8249 3341 8283 3375
rect 9445 3341 9479 3375
rect 9721 3341 9755 3375
rect 17357 3341 17391 3375
rect 17909 3341 17943 3375
rect 23613 3341 23647 3375
rect 1441 3273 1475 3307
rect 1717 3273 1751 3307
rect 4661 3273 4695 3307
rect 6961 3273 6995 3307
rect 11929 3273 11963 3307
rect 12205 3273 12239 3307
rect 15701 3273 15735 3307
rect 23889 3273 23923 3307
rect 3373 3205 3407 3239
rect 5121 3205 5155 3239
rect 5949 3205 5983 3239
rect 6225 3205 6259 3239
rect 11745 3205 11779 3239
rect 12021 3205 12055 3239
rect 22693 3205 22727 3239
rect 23337 3205 23371 3239
rect 23521 3205 23555 3239
rect 25637 3205 25671 3239
rect 797 3001 831 3035
rect 981 3001 1015 3035
rect 9077 3001 9111 3035
rect 24257 3001 24291 3035
rect 1625 2933 1659 2967
rect 1717 2933 1751 2967
rect 18093 2933 18127 2967
rect 1441 2865 1475 2899
rect 4477 2865 4511 2899
rect 6961 2865 6995 2899
rect 11745 2865 11779 2899
rect 13217 2865 13251 2899
rect 15517 2865 15551 2899
rect 18829 2865 18863 2899
rect 21405 2865 21439 2899
rect 21497 2865 21531 2899
rect 22141 2865 22175 2899
rect 22417 2865 22451 2899
rect 23521 2865 23555 2899
rect 23705 2865 23739 2899
rect 1165 2797 1199 2831
rect 7513 2797 7547 2831
rect 13309 2797 13343 2831
rect 14965 2797 14999 2831
rect 18001 2797 18035 2831
rect 18921 2797 18955 2831
rect 20485 2797 20519 2831
rect 21129 2797 21163 2831
rect 7421 2729 7455 2763
rect 15425 2729 15459 2763
rect 20669 2729 20703 2763
rect 20761 2729 20795 2763
rect 6777 2661 6811 2695
rect 9997 2661 10031 2695
rect 15701 2661 15735 2695
rect 23797 2661 23831 2695
rect 24441 2661 24475 2695
rect 2361 2457 2395 2491
rect 5121 2457 5155 2491
rect 6501 2457 6535 2491
rect 6685 2457 6719 2491
rect 11837 2457 11871 2491
rect 12573 2457 12607 2491
rect 14413 2457 14447 2491
rect 14597 2457 14631 2491
rect 14781 2457 14815 2491
rect 17449 2457 17483 2491
rect 17633 2457 17667 2491
rect 17909 2457 17943 2491
rect 22141 2457 22175 2491
rect 22325 2457 22359 2491
rect 23797 2457 23831 2491
rect 23981 2457 24015 2491
rect 25867 2457 25901 2491
rect 8065 2389 8099 2423
rect 20301 2389 20335 2423
rect 22601 2389 22635 2423
rect 23061 2389 23095 2423
rect 889 2321 923 2355
rect 1073 2321 1107 2355
rect 9629 2321 9663 2355
rect 11929 2321 11963 2355
rect 12481 2321 12515 2355
rect 12757 2321 12791 2355
rect 17173 2321 17207 2355
rect 20945 2321 20979 2355
rect 24165 2321 24199 2355
rect 24441 2321 24475 2355
rect 26189 2321 26223 2355
rect 1349 2253 1383 2287
rect 2269 2253 2303 2287
rect 3281 2253 3315 2287
rect 3557 2253 3591 2287
rect 6777 2253 6811 2287
rect 7789 2253 7823 2287
rect 9905 2253 9939 2287
rect 10641 2253 10675 2287
rect 12389 2253 12423 2287
rect 13861 2253 13895 2287
rect 14137 2253 14171 2287
rect 14873 2253 14907 2287
rect 15793 2253 15827 2287
rect 16529 2253 16563 2287
rect 18001 2253 18035 2287
rect 19703 2253 19737 2287
rect 20485 2253 20519 2287
rect 21497 2253 21531 2287
rect 21773 2253 21807 2287
rect 21957 2253 21991 2287
rect 22969 2253 23003 2287
rect 1993 2185 2027 2219
rect 4477 2185 4511 2219
rect 4661 2185 4695 2219
rect 4937 2185 4971 2219
rect 10825 2185 10859 2219
rect 11377 2185 11411 2219
rect 11561 2185 11595 2219
rect 16437 2185 16471 2219
rect 18277 2185 18311 2219
rect 20669 2185 20703 2219
rect 22693 2185 22727 2219
rect 1257 2117 1291 2151
rect 3097 2117 3131 2151
rect 3373 2117 3407 2151
rect 4753 2117 4787 2151
rect 6225 2117 6259 2151
rect 9813 2117 9847 2151
rect 13677 2117 13711 2151
rect 13953 2117 13987 2151
rect 20025 2117 20059 2151
rect 20853 2117 20887 2151
rect 23521 2117 23555 2151
rect 7053 1913 7087 1947
rect 11837 1913 11871 1947
rect 18369 1913 18403 1947
rect 18645 1913 18679 1947
rect 20669 1913 20703 1947
rect 23521 1913 23555 1947
rect 23889 1913 23923 1947
rect 24257 1913 24291 1947
rect 24441 1913 24475 1947
rect 25913 1913 25947 1947
rect 6777 1845 6811 1879
rect 7145 1845 7179 1879
rect 9169 1845 9203 1879
rect 11377 1845 11411 1879
rect 15517 1845 15551 1879
rect 15701 1845 15735 1879
rect 18093 1845 18127 1879
rect 19289 1845 19323 1879
rect 23245 1845 23279 1879
rect 24165 1845 24199 1879
rect 1533 1777 1567 1811
rect 2269 1777 2303 1811
rect 3741 1777 3775 1811
rect 4569 1777 4603 1811
rect 5857 1777 5891 1811
rect 6593 1777 6627 1811
rect 7789 1777 7823 1811
rect 9077 1777 9111 1811
rect 9905 1777 9939 1811
rect 12573 1777 12607 1811
rect 13401 1777 13435 1811
rect 14597 1777 14631 1811
rect 15241 1777 15275 1811
rect 16529 1777 16563 1811
rect 18737 1777 18771 1811
rect 18921 1777 18955 1811
rect 20853 1777 20887 1811
rect 23429 1777 23463 1811
rect 26097 1777 26131 1811
rect 1441 1709 1475 1743
rect 2361 1709 2395 1743
rect 3833 1709 3867 1743
rect 4661 1709 4695 1743
rect 9997 1709 10031 1743
rect 10917 1709 10951 1743
rect 11469 1709 11503 1743
rect 12665 1709 12699 1743
rect 13493 1709 13527 1743
rect 18185 1709 18219 1743
rect 21773 1709 21807 1743
rect 7605 1573 7639 1607
rect 16345 1573 16379 1607
rect 17909 1573 17943 1607
rect 1257 1369 1291 1403
rect 2085 1369 2119 1403
rect 2269 1369 2303 1403
rect 3097 1369 3131 1403
rect 3465 1369 3499 1403
rect 7053 1369 7087 1403
rect 7789 1369 7823 1403
rect 8341 1369 8375 1403
rect 8893 1369 8927 1403
rect 9721 1369 9755 1403
rect 10089 1369 10123 1403
rect 10917 1369 10951 1403
rect 11193 1369 11227 1403
rect 11745 1369 11779 1403
rect 12021 1369 12055 1403
rect 12205 1369 12239 1403
rect 12757 1369 12791 1403
rect 16345 1369 16379 1403
rect 16713 1369 16747 1403
rect 19013 1369 19047 1403
rect 19289 1369 19323 1403
rect 19749 1369 19783 1403
rect 20577 1369 20611 1403
rect 20945 1369 20979 1403
rect 21497 1369 21531 1403
rect 23061 1369 23095 1403
rect 23245 1369 23279 1403
rect 23429 1369 23463 1403
rect 23797 1369 23831 1403
rect 26373 1369 26407 1403
rect 4201 1301 4235 1335
rect 9629 1301 9663 1335
rect 9997 1301 10031 1335
rect 12849 1301 12883 1335
rect 13033 1301 13067 1335
rect 15977 1301 16011 1335
rect 16529 1301 16563 1335
rect 19473 1301 19507 1335
rect 21221 1301 21255 1335
rect 4017 1233 4051 1267
rect 6685 1233 6719 1267
rect 7605 1233 7639 1267
rect 8157 1233 8191 1267
rect 9077 1233 9111 1267
rect 11377 1233 11411 1267
rect 14413 1233 14447 1267
rect 15057 1233 15091 1267
rect 15241 1233 15275 1267
rect 15333 1233 15367 1267
rect 21313 1233 21347 1267
rect 24349 1233 24383 1267
rect 26097 1233 26131 1267
rect 1073 1165 1107 1199
rect 1349 1165 1383 1199
rect 3373 1165 3407 1199
rect 5857 1165 5891 1199
rect 6133 1165 6167 1199
rect 6777 1165 6811 1199
rect 9261 1165 9295 1199
rect 11929 1165 11963 1199
rect 14505 1165 14539 1199
rect 15885 1165 15919 1199
rect 16161 1165 16195 1199
rect 17909 1165 17943 1199
rect 18369 1165 18403 1199
rect 19289 1165 19323 1199
rect 19841 1165 19875 1199
rect 20669 1165 20703 1199
rect 24073 1165 24107 1199
rect 25775 1165 25809 1199
rect 889 1097 923 1131
rect 1809 1097 1843 1131
rect 1901 1097 1935 1131
rect 3189 1097 3223 1131
rect 5581 1097 5615 1131
rect 5765 1097 5799 1131
rect 6593 1097 6627 1131
rect 7513 1097 7547 1131
rect 7973 1097 8007 1131
rect 9445 1097 9479 1131
rect 14045 1097 14079 1131
rect 14229 1097 14263 1131
rect 14965 1097 14999 1131
rect 18829 1097 18863 1131
rect 3925 1029 3959 1063
rect 4385 1029 4419 1063
rect 12481 1029 12515 1063
rect 18185 1029 18219 1063
rect 18645 1029 18679 1063
rect 23981 1029 24015 1063
rect 26281 1029 26315 1063
rect 1349 825 1383 859
rect 1625 825 1659 859
rect 3649 825 3683 859
rect 3833 825 3867 859
rect 5949 825 5983 859
rect 14873 825 14907 859
rect 24165 825 24199 859
rect 24349 757 24383 791
<< metal1 >>
rect 25438 27268 25444 27320
rect 25496 27308 25502 27320
rect 26358 27308 26364 27320
rect 25496 27280 26364 27308
rect 25496 27268 25502 27280
rect 26358 27268 26364 27280
rect 26416 27268 26422 27320
rect 400 27082 27264 27104
rect 400 27030 18870 27082
rect 18922 27030 18934 27082
rect 18986 27030 18998 27082
rect 19050 27030 19062 27082
rect 19114 27030 19126 27082
rect 19178 27030 27264 27082
rect 400 27008 27264 27030
rect 6210 26764 6216 26776
rect 6171 26736 6216 26764
rect 6210 26724 6216 26736
rect 6268 26724 6274 26776
rect 6486 26724 6492 26776
rect 6544 26764 6550 26776
rect 6765 26767 6823 26773
rect 6765 26764 6777 26767
rect 6544 26736 6777 26764
rect 6544 26724 6550 26736
rect 6765 26733 6777 26736
rect 6811 26733 6823 26767
rect 6765 26727 6823 26733
rect 6670 26696 6676 26708
rect 6631 26668 6676 26696
rect 6670 26656 6676 26668
rect 6728 26656 6734 26708
rect 7501 26631 7559 26637
rect 7501 26597 7513 26631
rect 7547 26628 7559 26631
rect 7682 26628 7688 26640
rect 7547 26600 7688 26628
rect 7547 26597 7559 26600
rect 7501 26591 7559 26597
rect 7682 26588 7688 26600
rect 7740 26588 7746 26640
rect 23877 26631 23935 26637
rect 23877 26597 23889 26631
rect 23923 26628 23935 26631
rect 24058 26628 24064 26640
rect 23923 26600 24064 26628
rect 23923 26597 23935 26600
rect 23877 26591 23935 26597
rect 24058 26588 24064 26600
rect 24116 26588 24122 26640
rect 400 26538 27264 26560
rect 400 26486 3510 26538
rect 3562 26486 3574 26538
rect 3626 26486 3638 26538
rect 3690 26486 3702 26538
rect 3754 26486 3766 26538
rect 3818 26486 27264 26538
rect 400 26464 27264 26486
rect 6670 26424 6676 26436
rect 6631 26396 6676 26424
rect 6670 26384 6676 26396
rect 6728 26384 6734 26436
rect 23325 26427 23383 26433
rect 23325 26393 23337 26427
rect 23371 26424 23383 26427
rect 23598 26424 23604 26436
rect 23371 26396 23604 26424
rect 23371 26393 23383 26396
rect 23325 26387 23383 26393
rect 23598 26384 23604 26396
rect 23656 26424 23662 26436
rect 23656 26396 25852 26424
rect 23656 26384 23662 26396
rect 2533 26359 2591 26365
rect 2533 26325 2545 26359
rect 2579 26356 2591 26359
rect 3910 26356 3916 26368
rect 2579 26328 3916 26356
rect 2579 26325 2591 26328
rect 2533 26319 2591 26325
rect 2162 26220 2168 26232
rect 2075 26192 2168 26220
rect 2162 26180 2168 26192
rect 2220 26220 2226 26232
rect 2548 26220 2576 26319
rect 3910 26316 3916 26328
rect 3968 26316 3974 26368
rect 4278 26316 4284 26368
rect 4336 26356 4342 26368
rect 4336 26328 14352 26356
rect 4336 26316 4342 26328
rect 2990 26288 2996 26300
rect 2903 26260 2996 26288
rect 2990 26248 2996 26260
rect 3048 26288 3054 26300
rect 3637 26291 3695 26297
rect 3637 26288 3649 26291
rect 3048 26260 3649 26288
rect 3048 26248 3054 26260
rect 3637 26257 3649 26260
rect 3683 26257 3695 26291
rect 3637 26251 3695 26257
rect 7133 26291 7191 26297
rect 7133 26257 7145 26291
rect 7179 26288 7191 26291
rect 8421 26291 8479 26297
rect 8421 26288 8433 26291
rect 7179 26260 8433 26288
rect 7179 26257 7191 26260
rect 7133 26251 7191 26257
rect 8421 26257 8433 26260
rect 8467 26288 8479 26291
rect 12190 26288 12196 26300
rect 8467 26260 12196 26288
rect 8467 26257 8479 26260
rect 8421 26251 8479 26257
rect 12190 26248 12196 26260
rect 12248 26248 12254 26300
rect 2220 26192 2576 26220
rect 3085 26223 3143 26229
rect 2220 26180 2226 26192
rect 3085 26189 3097 26223
rect 3131 26220 3143 26223
rect 3358 26220 3364 26232
rect 3131 26192 3364 26220
rect 3131 26189 3143 26192
rect 3085 26183 3143 26189
rect 3358 26180 3364 26192
rect 3416 26220 3422 26232
rect 3821 26223 3879 26229
rect 3821 26220 3833 26223
rect 3416 26192 3833 26220
rect 3416 26180 3422 26192
rect 3821 26189 3833 26192
rect 3867 26220 3879 26223
rect 3867 26192 4554 26220
rect 3867 26189 3879 26192
rect 3821 26183 3879 26189
rect 3545 26155 3603 26161
rect 3545 26121 3557 26155
rect 3591 26121 3603 26155
rect 4526 26152 4554 26192
rect 6394 26180 6400 26232
rect 6452 26220 6458 26232
rect 7225 26223 7283 26229
rect 7225 26220 7237 26223
rect 6452 26192 7237 26220
rect 6452 26180 6458 26192
rect 7225 26189 7237 26192
rect 7271 26220 7283 26223
rect 7314 26220 7320 26232
rect 7271 26192 7320 26220
rect 7271 26189 7283 26192
rect 7225 26183 7283 26189
rect 7314 26180 7320 26192
rect 7372 26180 7378 26232
rect 7501 26223 7559 26229
rect 7501 26189 7513 26223
rect 7547 26220 7559 26223
rect 7682 26220 7688 26232
rect 7547 26192 7688 26220
rect 7547 26189 7559 26192
rect 7501 26183 7559 26189
rect 7682 26180 7688 26192
rect 7740 26180 7746 26232
rect 8329 26223 8387 26229
rect 8329 26189 8341 26223
rect 8375 26189 8387 26223
rect 11730 26220 11736 26232
rect 11643 26192 11736 26220
rect 8329 26183 8387 26189
rect 7406 26152 7412 26164
rect 4526 26124 7412 26152
rect 3545 26115 3603 26121
rect 1702 26044 1708 26096
rect 1760 26084 1766 26096
rect 1981 26087 2039 26093
rect 1981 26084 1993 26087
rect 1760 26056 1993 26084
rect 1760 26044 1766 26056
rect 1981 26053 1993 26056
rect 2027 26084 2039 26087
rect 2257 26087 2315 26093
rect 2257 26084 2269 26087
rect 2027 26056 2269 26084
rect 2027 26053 2039 26056
rect 1981 26047 2039 26053
rect 2257 26053 2269 26056
rect 2303 26053 2315 26087
rect 3560 26084 3588 26115
rect 7406 26112 7412 26124
rect 7464 26152 7470 26164
rect 7593 26155 7651 26161
rect 7593 26152 7605 26155
rect 7464 26124 7605 26152
rect 7464 26112 7470 26124
rect 7593 26121 7605 26124
rect 7639 26121 7651 26155
rect 7593 26115 7651 26121
rect 4005 26087 4063 26093
rect 4005 26084 4017 26087
rect 3560 26056 4017 26084
rect 2257 26047 2315 26053
rect 4005 26053 4017 26056
rect 4051 26084 4063 26087
rect 4186 26084 4192 26096
rect 4051 26056 4192 26084
rect 4051 26053 4063 26056
rect 4005 26047 4063 26053
rect 4186 26044 4192 26056
rect 4244 26044 4250 26096
rect 6210 26084 6216 26096
rect 6171 26056 6216 26084
rect 6210 26044 6216 26056
rect 6268 26044 6274 26096
rect 6486 26084 6492 26096
rect 6447 26056 6492 26084
rect 6486 26044 6492 26056
rect 6544 26044 6550 26096
rect 7314 26044 7320 26096
rect 7372 26084 7378 26096
rect 8344 26084 8372 26183
rect 11730 26180 11736 26192
rect 11788 26220 11794 26232
rect 14324 26229 14352 26328
rect 17710 26316 17716 26368
rect 17768 26356 17774 26368
rect 18357 26359 18415 26365
rect 18357 26356 18369 26359
rect 17768 26328 18369 26356
rect 17768 26316 17774 26328
rect 18357 26325 18369 26328
rect 18403 26356 18415 26359
rect 18403 26328 21620 26356
rect 18403 26325 18415 26328
rect 18357 26319 18415 26325
rect 14493 26291 14551 26297
rect 14493 26257 14505 26291
rect 14539 26288 14551 26291
rect 14861 26291 14919 26297
rect 14861 26288 14873 26291
rect 14539 26260 14873 26288
rect 14539 26257 14551 26260
rect 14493 26251 14551 26257
rect 14861 26257 14873 26260
rect 14907 26288 14919 26291
rect 19274 26288 19280 26300
rect 14907 26260 19280 26288
rect 14907 26257 14919 26260
rect 14861 26251 14919 26257
rect 19274 26248 19280 26260
rect 19332 26248 19338 26300
rect 21592 26288 21620 26328
rect 22221 26291 22279 26297
rect 22221 26288 22233 26291
rect 21592 26260 22233 26288
rect 12377 26223 12435 26229
rect 12377 26220 12389 26223
rect 11788 26192 12389 26220
rect 11788 26180 11794 26192
rect 12377 26189 12389 26192
rect 12423 26189 12435 26223
rect 12377 26183 12435 26189
rect 14309 26223 14367 26229
rect 14309 26189 14321 26223
rect 14355 26220 14367 26223
rect 14585 26223 14643 26229
rect 14585 26220 14597 26223
rect 14355 26192 14597 26220
rect 14355 26189 14367 26192
rect 14309 26183 14367 26189
rect 14585 26189 14597 26192
rect 14631 26189 14643 26223
rect 14585 26183 14643 26189
rect 15965 26223 16023 26229
rect 15965 26189 15977 26223
rect 16011 26220 16023 26223
rect 16011 26192 16468 26220
rect 16011 26189 16023 26192
rect 15965 26183 16023 26189
rect 11549 26155 11607 26161
rect 11549 26121 11561 26155
rect 11595 26152 11607 26155
rect 12190 26152 12196 26164
rect 11595 26124 12196 26152
rect 11595 26121 11607 26124
rect 11549 26115 11607 26121
rect 12190 26112 12196 26124
rect 12248 26112 12254 26164
rect 12285 26155 12343 26161
rect 12285 26121 12297 26155
rect 12331 26152 12343 26155
rect 12466 26152 12472 26164
rect 12331 26124 12472 26152
rect 12331 26121 12343 26124
rect 12285 26115 12343 26121
rect 12466 26112 12472 26124
rect 12524 26152 12530 26164
rect 12561 26155 12619 26161
rect 12561 26152 12573 26155
rect 12524 26124 12573 26152
rect 12524 26112 12530 26124
rect 12561 26121 12573 26124
rect 12607 26121 12619 26155
rect 12561 26115 12619 26121
rect 14858 26112 14864 26164
rect 14916 26152 14922 26164
rect 16057 26155 16115 26161
rect 16057 26152 16069 26155
rect 14916 26124 16069 26152
rect 14916 26112 14922 26124
rect 16057 26121 16069 26124
rect 16103 26152 16115 26155
rect 16149 26155 16207 26161
rect 16149 26152 16161 26155
rect 16103 26124 16161 26152
rect 16103 26121 16115 26124
rect 16057 26115 16115 26121
rect 16149 26121 16161 26124
rect 16195 26121 16207 26155
rect 16149 26115 16207 26121
rect 9062 26084 9068 26096
rect 7372 26056 9068 26084
rect 7372 26044 7378 26056
rect 9062 26044 9068 26056
rect 9120 26044 9126 26096
rect 16440 26093 16468 26192
rect 16514 26180 16520 26232
rect 16572 26220 16578 26232
rect 17710 26220 17716 26232
rect 16572 26192 17716 26220
rect 16572 26180 16578 26192
rect 17710 26180 17716 26192
rect 17768 26180 17774 26232
rect 21592 26229 21620 26260
rect 22221 26257 22233 26260
rect 22267 26288 22279 26291
rect 23690 26288 23696 26300
rect 22267 26260 23696 26288
rect 22267 26257 22279 26260
rect 22221 26251 22279 26257
rect 23690 26248 23696 26260
rect 23748 26248 23754 26300
rect 24058 26288 24064 26300
rect 24019 26260 24064 26288
rect 24058 26248 24064 26260
rect 24116 26248 24122 26300
rect 25824 26297 25852 26396
rect 25809 26291 25867 26297
rect 25809 26257 25821 26291
rect 25855 26257 25867 26291
rect 25809 26251 25867 26257
rect 19921 26223 19979 26229
rect 19921 26189 19933 26223
rect 19967 26189 19979 26223
rect 19921 26183 19979 26189
rect 21577 26223 21635 26229
rect 21577 26189 21589 26223
rect 21623 26189 21635 26223
rect 23785 26223 23843 26229
rect 23785 26220 23797 26223
rect 21577 26183 21635 26189
rect 23524 26192 23797 26220
rect 17989 26155 18047 26161
rect 17989 26121 18001 26155
rect 18035 26152 18047 26155
rect 18035 26124 18400 26152
rect 18035 26121 18047 26124
rect 17989 26115 18047 26121
rect 18372 26096 18400 26124
rect 16425 26087 16483 26093
rect 16425 26053 16437 26087
rect 16471 26084 16483 26087
rect 17894 26084 17900 26096
rect 16471 26056 17900 26084
rect 16471 26053 16483 26056
rect 16425 26047 16483 26053
rect 17894 26044 17900 26056
rect 17952 26044 17958 26096
rect 18354 26044 18360 26096
rect 18412 26084 18418 26096
rect 18449 26087 18507 26093
rect 18449 26084 18461 26087
rect 18412 26056 18461 26084
rect 18412 26044 18418 26056
rect 18449 26053 18461 26056
rect 18495 26053 18507 26087
rect 19936 26084 19964 26183
rect 20013 26155 20071 26161
rect 20013 26121 20025 26155
rect 20059 26152 20071 26155
rect 20105 26155 20163 26161
rect 20105 26152 20117 26155
rect 20059 26124 20117 26152
rect 20059 26121 20071 26124
rect 20013 26115 20071 26121
rect 20105 26121 20117 26124
rect 20151 26152 20163 26155
rect 20470 26152 20476 26164
rect 20151 26124 20476 26152
rect 20151 26121 20163 26124
rect 20105 26115 20163 26121
rect 20470 26112 20476 26124
rect 20528 26112 20534 26164
rect 21850 26152 21856 26164
rect 21763 26124 21856 26152
rect 21850 26112 21856 26124
rect 21908 26152 21914 26164
rect 22313 26155 22371 26161
rect 22313 26152 22325 26155
rect 21908 26124 22325 26152
rect 21908 26112 21914 26124
rect 22313 26121 22325 26124
rect 22359 26121 22371 26155
rect 22313 26115 22371 26121
rect 23524 26096 23552 26192
rect 23785 26189 23797 26192
rect 23831 26189 23843 26223
rect 23785 26183 23843 26189
rect 20381 26087 20439 26093
rect 20381 26084 20393 26087
rect 19936 26056 20393 26084
rect 18449 26047 18507 26053
rect 20381 26053 20393 26056
rect 20427 26084 20439 26087
rect 20562 26084 20568 26096
rect 20427 26056 20568 26084
rect 20427 26053 20439 26056
rect 20381 26047 20439 26053
rect 20562 26044 20568 26056
rect 20620 26044 20626 26096
rect 23506 26084 23512 26096
rect 23467 26056 23512 26084
rect 23506 26044 23512 26056
rect 23564 26044 23570 26096
rect 23690 26084 23696 26096
rect 23603 26056 23696 26084
rect 23690 26044 23696 26056
rect 23748 26084 23754 26096
rect 24426 26084 24432 26096
rect 23748 26056 24432 26084
rect 23748 26044 23754 26056
rect 24426 26044 24432 26056
rect 24484 26084 24490 26096
rect 24536 26084 24564 26152
rect 24484 26056 24564 26084
rect 24484 26044 24490 26056
rect 400 25994 27264 26016
rect 400 25942 18870 25994
rect 18922 25942 18934 25994
rect 18986 25942 18998 25994
rect 19050 25942 19062 25994
rect 19114 25942 19126 25994
rect 19178 25942 27264 25994
rect 400 25920 27264 25942
rect 7406 25880 7412 25892
rect 7367 25852 7412 25880
rect 7406 25840 7412 25852
rect 7464 25840 7470 25892
rect 2073 25815 2131 25821
rect 2073 25781 2085 25815
rect 2119 25812 2131 25815
rect 2162 25812 2168 25824
rect 2119 25784 2168 25812
rect 2119 25781 2131 25784
rect 2073 25775 2131 25781
rect 2162 25772 2168 25784
rect 2220 25772 2226 25824
rect 8326 25812 8332 25824
rect 6780 25784 8332 25812
rect 6780 25756 6808 25784
rect 8326 25772 8332 25784
rect 8384 25772 8390 25824
rect 9246 25772 9252 25824
rect 9304 25812 9310 25824
rect 9341 25815 9399 25821
rect 9341 25812 9353 25815
rect 9304 25784 9353 25812
rect 9304 25772 9310 25784
rect 9341 25781 9353 25784
rect 9387 25781 9399 25815
rect 11730 25812 11736 25824
rect 11691 25784 11736 25812
rect 9341 25775 9399 25781
rect 11730 25772 11736 25784
rect 11788 25772 11794 25824
rect 14858 25812 14864 25824
rect 14819 25784 14864 25812
rect 14858 25772 14864 25784
rect 14916 25772 14922 25824
rect 15870 25772 15876 25824
rect 15928 25772 15934 25824
rect 21850 25772 21856 25824
rect 21908 25772 21914 25824
rect 966 25704 972 25756
rect 1024 25744 1030 25756
rect 1153 25747 1211 25753
rect 1153 25744 1165 25747
rect 1024 25716 1165 25744
rect 1024 25704 1030 25716
rect 1153 25713 1165 25716
rect 1199 25713 1211 25747
rect 1886 25744 1892 25756
rect 1847 25716 1892 25744
rect 1153 25707 1211 25713
rect 1886 25704 1892 25716
rect 1944 25704 1950 25756
rect 3358 25744 3364 25756
rect 3319 25716 3364 25744
rect 3358 25704 3364 25716
rect 3416 25704 3422 25756
rect 4278 25744 4284 25756
rect 4239 25716 4284 25744
rect 4278 25704 4284 25716
rect 4336 25704 4342 25756
rect 6394 25704 6400 25756
rect 6452 25744 6458 25756
rect 6673 25747 6731 25753
rect 6673 25744 6685 25747
rect 6452 25716 6685 25744
rect 6452 25704 6458 25716
rect 6673 25713 6685 25716
rect 6719 25713 6731 25747
rect 6673 25707 6731 25713
rect 6762 25704 6768 25756
rect 6820 25744 6826 25756
rect 7869 25747 7927 25753
rect 6820 25716 6913 25744
rect 6820 25704 6826 25716
rect 7869 25713 7881 25747
rect 7915 25744 7927 25747
rect 10074 25744 10080 25756
rect 7915 25716 8280 25744
rect 10035 25716 10080 25744
rect 7915 25713 7927 25716
rect 7869 25707 7927 25713
rect 5382 25636 5388 25688
rect 5440 25676 5446 25688
rect 5845 25679 5903 25685
rect 5845 25676 5857 25679
rect 5440 25648 5857 25676
rect 5440 25636 5446 25648
rect 5845 25645 5857 25648
rect 5891 25645 5903 25679
rect 5845 25639 5903 25645
rect 5937 25679 5995 25685
rect 5937 25645 5949 25679
rect 5983 25676 5995 25679
rect 6210 25676 6216 25688
rect 5983 25648 6216 25676
rect 5983 25645 5995 25648
rect 5937 25639 5995 25645
rect 6210 25636 6216 25648
rect 6268 25636 6274 25688
rect 4186 25568 4192 25620
rect 4244 25608 4250 25620
rect 4649 25611 4707 25617
rect 4649 25608 4661 25611
rect 4244 25580 4661 25608
rect 4244 25568 4250 25580
rect 4649 25577 4661 25580
rect 4695 25577 4707 25611
rect 4649 25571 4707 25577
rect 6486 25500 6492 25552
rect 6544 25540 6550 25552
rect 7685 25543 7743 25549
rect 7685 25540 7697 25543
rect 6544 25512 7697 25540
rect 6544 25500 6550 25512
rect 7685 25509 7697 25512
rect 7731 25540 7743 25543
rect 7774 25540 7780 25552
rect 7731 25512 7780 25540
rect 7731 25509 7743 25512
rect 7685 25503 7743 25509
rect 7774 25500 7780 25512
rect 7832 25500 7838 25552
rect 8252 25549 8280 25716
rect 10074 25704 10080 25716
rect 10132 25704 10138 25756
rect 10169 25747 10227 25753
rect 10169 25713 10181 25747
rect 10215 25744 10227 25747
rect 10258 25744 10264 25756
rect 10215 25716 10264 25744
rect 10215 25713 10227 25716
rect 10169 25707 10227 25713
rect 10258 25704 10264 25716
rect 10316 25744 10322 25756
rect 12374 25744 12380 25756
rect 10316 25716 12380 25744
rect 10316 25704 10322 25716
rect 12374 25704 12380 25716
rect 12432 25744 12438 25756
rect 12469 25747 12527 25753
rect 12469 25744 12481 25747
rect 12432 25716 12481 25744
rect 12432 25704 12438 25716
rect 12469 25713 12481 25716
rect 12515 25713 12527 25747
rect 12469 25707 12527 25713
rect 17437 25747 17495 25753
rect 17437 25713 17449 25747
rect 17483 25744 17495 25747
rect 18354 25744 18360 25756
rect 17483 25716 18360 25744
rect 17483 25713 17495 25716
rect 17437 25707 17495 25713
rect 18354 25704 18360 25716
rect 18412 25704 18418 25756
rect 18817 25747 18875 25753
rect 18817 25713 18829 25747
rect 18863 25744 18875 25747
rect 19642 25744 19648 25756
rect 18863 25716 19648 25744
rect 18863 25713 18875 25716
rect 18817 25707 18875 25713
rect 19642 25704 19648 25716
rect 19700 25704 19706 25756
rect 9154 25636 9160 25688
rect 9212 25676 9218 25688
rect 9249 25679 9307 25685
rect 9249 25676 9261 25679
rect 9212 25648 9261 25676
rect 9212 25636 9218 25648
rect 9249 25645 9261 25648
rect 9295 25645 9307 25679
rect 9249 25639 9307 25645
rect 11086 25636 11092 25688
rect 11144 25676 11150 25688
rect 11641 25679 11699 25685
rect 11641 25676 11653 25679
rect 11144 25648 11653 25676
rect 11144 25636 11150 25648
rect 11641 25645 11653 25648
rect 11687 25645 11699 25679
rect 12558 25676 12564 25688
rect 12519 25648 12564 25676
rect 11641 25639 11699 25645
rect 12558 25636 12564 25648
rect 12616 25676 12622 25688
rect 14214 25676 14220 25688
rect 12616 25648 14220 25676
rect 12616 25636 12622 25648
rect 14214 25636 14220 25648
rect 14272 25636 14278 25688
rect 14398 25636 14404 25688
rect 14456 25676 14462 25688
rect 14585 25679 14643 25685
rect 14585 25676 14597 25679
rect 14456 25648 14597 25676
rect 14456 25636 14462 25648
rect 14585 25645 14597 25648
rect 14631 25645 14643 25679
rect 14585 25639 14643 25645
rect 15226 25636 15232 25688
rect 15284 25676 15290 25688
rect 16146 25676 16152 25688
rect 15284 25648 16152 25676
rect 15284 25636 15290 25648
rect 16146 25636 16152 25648
rect 16204 25676 16210 25688
rect 16609 25679 16667 25685
rect 16609 25676 16621 25679
rect 16204 25648 16621 25676
rect 16204 25636 16210 25648
rect 16609 25645 16621 25648
rect 16655 25645 16667 25679
rect 16609 25639 16667 25645
rect 17618 25636 17624 25688
rect 17676 25676 17682 25688
rect 17989 25679 18047 25685
rect 17989 25676 18001 25679
rect 17676 25648 18001 25676
rect 17676 25636 17682 25648
rect 17989 25645 18001 25648
rect 18035 25645 18047 25679
rect 17989 25639 18047 25645
rect 18541 25679 18599 25685
rect 18541 25645 18553 25679
rect 18587 25645 18599 25679
rect 18998 25676 19004 25688
rect 18959 25648 19004 25676
rect 18541 25639 18599 25645
rect 17710 25568 17716 25620
rect 17768 25608 17774 25620
rect 18556 25608 18584 25639
rect 18998 25636 19004 25648
rect 19056 25636 19062 25688
rect 20838 25676 20844 25688
rect 20799 25648 20844 25676
rect 20838 25636 20844 25648
rect 20896 25636 20902 25688
rect 21114 25676 21120 25688
rect 21075 25648 21120 25676
rect 21114 25636 21120 25648
rect 21172 25636 21178 25688
rect 22862 25676 22868 25688
rect 22823 25648 22868 25676
rect 22862 25636 22868 25648
rect 22920 25636 22926 25688
rect 19458 25608 19464 25620
rect 17768 25580 19464 25608
rect 17768 25568 17774 25580
rect 19458 25568 19464 25580
rect 19516 25608 19522 25620
rect 20654 25608 20660 25620
rect 19516 25580 20660 25608
rect 19516 25568 19522 25580
rect 20654 25568 20660 25580
rect 20712 25568 20718 25620
rect 8237 25543 8295 25549
rect 8237 25509 8249 25543
rect 8283 25540 8295 25543
rect 8418 25540 8424 25552
rect 8283 25512 8424 25540
rect 8283 25509 8295 25512
rect 8237 25503 8295 25509
rect 8418 25500 8424 25512
rect 8476 25500 8482 25552
rect 16790 25500 16796 25552
rect 16848 25540 16854 25552
rect 17897 25543 17955 25549
rect 17897 25540 17909 25543
rect 16848 25512 17909 25540
rect 16848 25500 16854 25512
rect 17897 25509 17909 25512
rect 17943 25540 17955 25543
rect 18998 25540 19004 25552
rect 17943 25512 19004 25540
rect 17943 25509 17955 25512
rect 17897 25503 17955 25509
rect 18998 25500 19004 25512
rect 19056 25500 19062 25552
rect 20470 25540 20476 25552
rect 20431 25512 20476 25540
rect 20470 25500 20476 25512
rect 20528 25500 20534 25552
rect 23969 25543 24027 25549
rect 23969 25509 23981 25543
rect 24015 25540 24027 25543
rect 24242 25540 24248 25552
rect 24015 25512 24248 25540
rect 24015 25509 24027 25512
rect 23969 25503 24027 25509
rect 24242 25500 24248 25512
rect 24300 25500 24306 25552
rect 400 25450 27264 25472
rect 400 25398 3510 25450
rect 3562 25398 3574 25450
rect 3626 25398 3638 25450
rect 3690 25398 3702 25450
rect 3754 25398 3766 25450
rect 3818 25398 27264 25450
rect 400 25376 27264 25398
rect 2625 25339 2683 25345
rect 2625 25305 2637 25339
rect 2671 25336 2683 25339
rect 2990 25336 2996 25348
rect 2671 25308 2996 25336
rect 2671 25305 2683 25308
rect 2625 25299 2683 25305
rect 2990 25296 2996 25308
rect 3048 25296 3054 25348
rect 3358 25336 3364 25348
rect 3319 25308 3364 25336
rect 3358 25296 3364 25308
rect 3416 25296 3422 25348
rect 3821 25339 3879 25345
rect 3821 25305 3833 25339
rect 3867 25336 3879 25339
rect 3910 25336 3916 25348
rect 3867 25308 3916 25336
rect 3867 25305 3879 25308
rect 3821 25299 3879 25305
rect 3910 25296 3916 25308
rect 3968 25336 3974 25348
rect 4278 25336 4284 25348
rect 3968 25308 4284 25336
rect 3968 25296 3974 25308
rect 4278 25296 4284 25308
rect 4336 25296 4342 25348
rect 5661 25339 5719 25345
rect 5661 25305 5673 25339
rect 5707 25336 5719 25339
rect 6762 25336 6768 25348
rect 5707 25308 6768 25336
rect 5707 25305 5719 25308
rect 5661 25299 5719 25305
rect 6762 25296 6768 25308
rect 6820 25296 6826 25348
rect 7774 25336 7780 25348
rect 7735 25308 7780 25336
rect 7774 25296 7780 25308
rect 7832 25296 7838 25348
rect 8973 25339 9031 25345
rect 8973 25305 8985 25339
rect 9019 25336 9031 25339
rect 10074 25336 10080 25348
rect 9019 25308 10080 25336
rect 9019 25305 9031 25308
rect 8973 25299 9031 25305
rect 10074 25296 10080 25308
rect 10132 25296 10138 25348
rect 11365 25339 11423 25345
rect 11365 25305 11377 25339
rect 11411 25336 11423 25339
rect 12558 25336 12564 25348
rect 11411 25308 12564 25336
rect 11411 25305 11423 25308
rect 11365 25299 11423 25305
rect 12558 25296 12564 25308
rect 12616 25296 12622 25348
rect 14677 25339 14735 25345
rect 14677 25305 14689 25339
rect 14723 25336 14735 25339
rect 14858 25336 14864 25348
rect 14723 25308 14864 25336
rect 14723 25305 14735 25308
rect 14677 25299 14735 25305
rect 14858 25296 14864 25308
rect 14916 25296 14922 25348
rect 15870 25336 15876 25348
rect 15336 25308 15876 25336
rect 10442 25268 10448 25280
rect 8528 25240 10448 25268
rect 1061 25203 1119 25209
rect 1061 25169 1073 25203
rect 1107 25200 1119 25203
rect 1702 25200 1708 25212
rect 1107 25172 1708 25200
rect 1107 25169 1119 25172
rect 1061 25163 1119 25169
rect 1702 25160 1708 25172
rect 1760 25160 1766 25212
rect 966 25092 972 25144
rect 1024 25132 1030 25144
rect 1153 25135 1211 25141
rect 1153 25132 1165 25135
rect 1024 25104 1165 25132
rect 1024 25092 1030 25104
rect 1153 25101 1165 25104
rect 1199 25132 1211 25135
rect 1797 25135 1855 25141
rect 1797 25132 1809 25135
rect 1199 25104 1809 25132
rect 1199 25101 1211 25104
rect 1153 25095 1211 25101
rect 1797 25101 1809 25104
rect 1843 25132 1855 25135
rect 1981 25135 2039 25141
rect 1981 25132 1993 25135
rect 1843 25104 1993 25132
rect 1843 25101 1855 25104
rect 1797 25095 1855 25101
rect 1981 25101 1993 25104
rect 2027 25101 2039 25135
rect 1981 25095 2039 25101
rect 5293 25135 5351 25141
rect 5293 25101 5305 25135
rect 5339 25132 5351 25135
rect 6210 25132 6216 25144
rect 5339 25104 6216 25132
rect 5339 25101 5351 25104
rect 5293 25095 5351 25101
rect 6210 25092 6216 25104
rect 6268 25092 6274 25144
rect 6670 25092 6676 25144
rect 6728 25132 6734 25144
rect 6857 25135 6915 25141
rect 6857 25132 6869 25135
rect 6728 25104 6869 25132
rect 6728 25092 6734 25104
rect 6857 25101 6869 25104
rect 6903 25132 6915 25135
rect 7225 25135 7283 25141
rect 7225 25132 7237 25135
rect 6903 25104 7237 25132
rect 6903 25101 6915 25104
rect 6857 25095 6915 25101
rect 7225 25101 7237 25104
rect 7271 25132 7283 25135
rect 7406 25132 7412 25144
rect 7271 25104 7412 25132
rect 7271 25101 7283 25104
rect 7225 25095 7283 25101
rect 7406 25092 7412 25104
rect 7464 25092 7470 25144
rect 877 25067 935 25073
rect 877 25033 889 25067
rect 923 25064 935 25067
rect 1613 25067 1671 25073
rect 1613 25064 1625 25067
rect 923 25036 1625 25064
rect 923 25033 935 25036
rect 877 25027 935 25033
rect 1613 25033 1625 25036
rect 1659 25064 1671 25067
rect 1886 25064 1892 25076
rect 1659 25036 1892 25064
rect 1659 25033 1671 25036
rect 1613 25027 1671 25033
rect 1886 25024 1892 25036
rect 1944 25064 1950 25076
rect 2533 25067 2591 25073
rect 2533 25064 2545 25067
rect 1944 25036 2545 25064
rect 1944 25024 1950 25036
rect 2533 25033 2545 25036
rect 2579 25064 2591 25067
rect 2809 25067 2867 25073
rect 2809 25064 2821 25067
rect 2579 25036 2821 25064
rect 2579 25033 2591 25036
rect 2533 25027 2591 25033
rect 2809 25033 2821 25036
rect 2855 25033 2867 25067
rect 2809 25027 2867 25033
rect 3637 25067 3695 25073
rect 3637 25033 3649 25067
rect 3683 25064 3695 25067
rect 4186 25064 4192 25076
rect 3683 25036 4192 25064
rect 3683 25033 3695 25036
rect 3637 25027 3695 25033
rect 4186 25024 4192 25036
rect 4244 25024 4250 25076
rect 8528 25073 8556 25240
rect 10442 25228 10448 25240
rect 10500 25268 10506 25280
rect 10537 25271 10595 25277
rect 10537 25268 10549 25271
rect 10500 25240 10549 25268
rect 10500 25228 10506 25240
rect 10537 25237 10549 25240
rect 10583 25237 10595 25271
rect 10537 25231 10595 25237
rect 14309 25271 14367 25277
rect 14309 25237 14321 25271
rect 14355 25268 14367 25271
rect 15226 25268 15232 25280
rect 14355 25240 15232 25268
rect 14355 25237 14367 25240
rect 14309 25231 14367 25237
rect 15226 25228 15232 25240
rect 15284 25228 15290 25280
rect 9062 25200 9068 25212
rect 9023 25172 9068 25200
rect 9062 25160 9068 25172
rect 9120 25200 9126 25212
rect 10258 25200 10264 25212
rect 9120 25172 10264 25200
rect 9120 25160 9126 25172
rect 10258 25160 10264 25172
rect 10316 25160 10322 25212
rect 15336 25209 15364 25308
rect 15870 25296 15876 25308
rect 15928 25296 15934 25348
rect 16790 25336 16796 25348
rect 16751 25308 16796 25336
rect 16790 25296 16796 25308
rect 16848 25296 16854 25348
rect 19458 25336 19464 25348
rect 19419 25308 19464 25336
rect 19458 25296 19464 25308
rect 19516 25296 19522 25348
rect 21942 25336 21948 25348
rect 21903 25308 21948 25336
rect 21942 25296 21948 25308
rect 22000 25296 22006 25348
rect 22221 25339 22279 25345
rect 22221 25305 22233 25339
rect 22267 25336 22279 25339
rect 22862 25336 22868 25348
rect 22267 25308 22868 25336
rect 22267 25305 22279 25308
rect 22221 25299 22279 25305
rect 22862 25296 22868 25308
rect 22920 25296 22926 25348
rect 15689 25271 15747 25277
rect 15689 25237 15701 25271
rect 15735 25268 15747 25271
rect 16514 25268 16520 25280
rect 15735 25240 16520 25268
rect 15735 25237 15747 25240
rect 15689 25231 15747 25237
rect 14861 25203 14919 25209
rect 14861 25169 14873 25203
rect 14907 25200 14919 25203
rect 15321 25203 15379 25209
rect 15321 25200 15333 25203
rect 14907 25172 15333 25200
rect 14907 25169 14919 25172
rect 14861 25163 14919 25169
rect 15321 25169 15333 25172
rect 15367 25169 15379 25203
rect 15321 25163 15379 25169
rect 9246 25132 9252 25144
rect 9207 25104 9252 25132
rect 9246 25092 9252 25104
rect 9304 25092 9310 25144
rect 9798 25092 9804 25144
rect 9856 25132 9862 25144
rect 10169 25135 10227 25141
rect 10169 25132 10181 25135
rect 9856 25104 10181 25132
rect 9856 25092 9862 25104
rect 10169 25101 10181 25104
rect 10215 25132 10227 25135
rect 10905 25135 10963 25141
rect 10905 25132 10917 25135
rect 10215 25104 10917 25132
rect 10215 25101 10227 25104
rect 10169 25095 10227 25101
rect 10905 25101 10917 25104
rect 10951 25101 10963 25135
rect 11730 25132 11736 25144
rect 11691 25104 11736 25132
rect 10905 25095 10963 25101
rect 7133 25067 7191 25073
rect 7133 25033 7145 25067
rect 7179 25033 7191 25067
rect 7133 25027 7191 25033
rect 8053 25067 8111 25073
rect 8053 25033 8065 25067
rect 8099 25064 8111 25067
rect 8237 25067 8295 25073
rect 8237 25064 8249 25067
rect 8099 25036 8249 25064
rect 8099 25033 8111 25036
rect 8053 25027 8111 25033
rect 8237 25033 8249 25036
rect 8283 25064 8295 25067
rect 8513 25067 8571 25073
rect 8513 25064 8525 25067
rect 8283 25036 8525 25064
rect 8283 25033 8295 25036
rect 8237 25027 8295 25033
rect 8513 25033 8525 25036
rect 8559 25033 8571 25067
rect 8513 25027 8571 25033
rect 8789 25067 8847 25073
rect 8789 25033 8801 25067
rect 8835 25064 8847 25067
rect 9154 25064 9160 25076
rect 8835 25036 9160 25064
rect 8835 25033 8847 25036
rect 8789 25027 8847 25033
rect 5382 24996 5388 25008
rect 5343 24968 5388 24996
rect 5382 24956 5388 24968
rect 5440 24956 5446 25008
rect 5474 24956 5480 25008
rect 5532 24996 5538 25008
rect 5753 24999 5811 25005
rect 5753 24996 5765 24999
rect 5532 24968 5765 24996
rect 5532 24956 5538 24968
rect 5753 24965 5765 24968
rect 5799 24965 5811 24999
rect 5753 24959 5811 24965
rect 6946 24956 6952 25008
rect 7004 24996 7010 25008
rect 7148 24996 7176 25027
rect 9154 25024 9160 25036
rect 9212 25024 9218 25076
rect 10920 25064 10948 25095
rect 11730 25092 11736 25104
rect 11788 25092 11794 25144
rect 12190 25092 12196 25144
rect 12248 25132 12254 25144
rect 12377 25135 12435 25141
rect 12377 25132 12389 25135
rect 12248 25104 12389 25132
rect 12248 25092 12254 25104
rect 12377 25101 12389 25104
rect 12423 25101 12435 25135
rect 12377 25095 12435 25101
rect 14950 25092 14956 25144
rect 15008 25132 15014 25144
rect 15045 25135 15103 25141
rect 15045 25132 15057 25135
rect 15008 25104 15057 25132
rect 15008 25092 15014 25104
rect 15045 25101 15057 25104
rect 15091 25132 15103 25135
rect 15704 25132 15732 25231
rect 16514 25228 16520 25240
rect 16572 25228 16578 25280
rect 20197 25271 20255 25277
rect 20197 25237 20209 25271
rect 20243 25268 20255 25271
rect 20381 25271 20439 25277
rect 20381 25268 20393 25271
rect 20243 25240 20393 25268
rect 20243 25237 20255 25240
rect 20197 25231 20255 25237
rect 20381 25237 20393 25240
rect 20427 25268 20439 25271
rect 21114 25268 21120 25280
rect 20427 25240 21120 25268
rect 20427 25237 20439 25240
rect 20381 25231 20439 25237
rect 21114 25228 21120 25240
rect 21172 25228 21178 25280
rect 16977 25203 17035 25209
rect 16977 25169 16989 25203
rect 17023 25200 17035 25203
rect 17161 25203 17219 25209
rect 17161 25200 17173 25203
rect 17023 25172 17173 25200
rect 17023 25169 17035 25172
rect 16977 25163 17035 25169
rect 17161 25169 17173 25172
rect 17207 25200 17219 25203
rect 17618 25200 17624 25212
rect 17207 25172 17624 25200
rect 17207 25169 17219 25172
rect 17161 25163 17219 25169
rect 17618 25160 17624 25172
rect 17676 25160 17682 25212
rect 17986 25160 17992 25212
rect 18044 25200 18050 25212
rect 19921 25203 19979 25209
rect 19921 25200 19933 25203
rect 18044 25172 19933 25200
rect 18044 25160 18050 25172
rect 19921 25169 19933 25172
rect 19967 25200 19979 25203
rect 21761 25203 21819 25209
rect 19967 25172 20976 25200
rect 19967 25169 19979 25172
rect 19921 25163 19979 25169
rect 17342 25132 17348 25144
rect 15091 25104 15732 25132
rect 17303 25104 17348 25132
rect 15091 25101 15103 25104
rect 15045 25095 15103 25101
rect 17342 25092 17348 25104
rect 17400 25092 17406 25144
rect 20470 25132 20476 25144
rect 20431 25104 20476 25132
rect 20470 25092 20476 25104
rect 20528 25092 20534 25144
rect 20654 25092 20660 25144
rect 20712 25132 20718 25144
rect 20841 25135 20899 25141
rect 20841 25132 20853 25135
rect 20712 25104 20853 25132
rect 20712 25092 20718 25104
rect 20841 25101 20853 25104
rect 20887 25101 20899 25135
rect 20948 25132 20976 25172
rect 21761 25169 21773 25203
rect 21807 25200 21819 25203
rect 22402 25200 22408 25212
rect 21807 25172 22408 25200
rect 21807 25169 21819 25172
rect 21761 25163 21819 25169
rect 22402 25160 22408 25172
rect 22460 25160 22466 25212
rect 24150 25160 24156 25212
rect 24208 25200 24214 25212
rect 25901 25203 25959 25209
rect 25901 25200 25913 25203
rect 24208 25172 25913 25200
rect 24208 25160 24214 25172
rect 25901 25169 25913 25172
rect 25947 25169 25959 25203
rect 25901 25163 25959 25169
rect 21485 25135 21543 25141
rect 21485 25132 21497 25135
rect 20948 25104 21497 25132
rect 20841 25095 20899 25101
rect 21485 25101 21497 25104
rect 21531 25132 21543 25135
rect 23414 25132 23420 25144
rect 21531 25104 23420 25132
rect 21531 25101 21543 25104
rect 21485 25095 21543 25101
rect 23414 25092 23420 25104
rect 23472 25092 23478 25144
rect 23877 25135 23935 25141
rect 23877 25132 23889 25135
rect 23524 25104 23889 25132
rect 12558 25064 12564 25076
rect 10920 25036 12564 25064
rect 12558 25024 12564 25036
rect 12616 25064 12622 25076
rect 12653 25067 12711 25073
rect 12653 25064 12665 25067
rect 12616 25036 12665 25064
rect 12616 25024 12622 25036
rect 12653 25033 12665 25036
rect 12699 25033 12711 25067
rect 12653 25027 12711 25033
rect 14398 25024 14404 25076
rect 14456 25064 14462 25076
rect 14493 25067 14551 25073
rect 14493 25064 14505 25067
rect 14456 25036 14505 25064
rect 14456 25024 14462 25036
rect 14493 25033 14505 25036
rect 14539 25064 14551 25067
rect 17360 25064 17388 25092
rect 14539 25036 17388 25064
rect 14539 25033 14551 25036
rect 14493 25027 14551 25033
rect 18354 25024 18360 25076
rect 18412 25024 18418 25076
rect 18998 25024 19004 25076
rect 19056 25064 19062 25076
rect 19369 25067 19427 25073
rect 19369 25064 19381 25067
rect 19056 25036 19381 25064
rect 19056 25024 19062 25036
rect 19369 25033 19381 25036
rect 19415 25064 19427 25067
rect 20562 25064 20568 25076
rect 19415 25036 20568 25064
rect 19415 25033 19427 25036
rect 19369 25027 19427 25033
rect 20562 25024 20568 25036
rect 20620 25024 20626 25076
rect 23524 25008 23552 25104
rect 23877 25101 23889 25104
rect 23923 25101 23935 25135
rect 23877 25095 23935 25101
rect 24153 25067 24211 25073
rect 24153 25033 24165 25067
rect 24199 25064 24211 25067
rect 24242 25064 24248 25076
rect 24199 25036 24248 25064
rect 24199 25033 24211 25036
rect 24153 25027 24211 25033
rect 24242 25024 24248 25036
rect 24300 25024 24306 25076
rect 24702 25024 24708 25076
rect 24760 25024 24766 25076
rect 7593 24999 7651 25005
rect 7593 24996 7605 24999
rect 7004 24968 7605 24996
rect 7004 24956 7010 24968
rect 7593 24965 7605 24968
rect 7639 24996 7651 24999
rect 8329 24999 8387 25005
rect 8329 24996 8341 24999
rect 7639 24968 8341 24996
rect 7639 24965 7651 24968
rect 7593 24959 7651 24965
rect 8329 24965 8341 24968
rect 8375 24996 8387 24999
rect 8418 24996 8424 25008
rect 8375 24968 8424 24996
rect 8375 24965 8387 24968
rect 8329 24959 8387 24965
rect 8418 24956 8424 24968
rect 8476 24956 8482 25008
rect 11086 24996 11092 25008
rect 11047 24968 11092 24996
rect 11086 24956 11092 24968
rect 11144 24956 11150 25008
rect 11549 24999 11607 25005
rect 11549 24965 11561 24999
rect 11595 24996 11607 24999
rect 12374 24996 12380 25008
rect 11595 24968 12380 24996
rect 11595 24965 11607 24968
rect 11549 24959 11607 24965
rect 12374 24956 12380 24968
rect 12432 24956 12438 25008
rect 19642 24996 19648 25008
rect 19603 24968 19648 24996
rect 19642 24956 19648 24968
rect 19700 24956 19706 25008
rect 23506 24996 23512 25008
rect 23467 24968 23512 24996
rect 23506 24956 23512 24968
rect 23564 24956 23570 25008
rect 23785 24999 23843 25005
rect 23785 24965 23797 24999
rect 23831 24996 23843 24999
rect 24720 24996 24748 25024
rect 23831 24968 24748 24996
rect 23831 24965 23843 24968
rect 23785 24959 23843 24965
rect 400 24906 27264 24928
rect 400 24854 18870 24906
rect 18922 24854 18934 24906
rect 18986 24854 18998 24906
rect 19050 24854 19062 24906
rect 19114 24854 19126 24906
rect 19178 24854 27264 24906
rect 400 24832 27264 24854
rect 874 24792 880 24804
rect 835 24764 880 24792
rect 874 24752 880 24764
rect 932 24752 938 24804
rect 1337 24795 1395 24801
rect 1337 24761 1349 24795
rect 1383 24792 1395 24795
rect 1886 24792 1892 24804
rect 1383 24764 1892 24792
rect 1383 24761 1395 24764
rect 1337 24755 1395 24761
rect 1886 24752 1892 24764
rect 1944 24752 1950 24804
rect 6210 24752 6216 24804
rect 6268 24792 6274 24804
rect 6673 24795 6731 24801
rect 6673 24792 6685 24795
rect 6268 24764 6685 24792
rect 6268 24752 6274 24764
rect 6673 24761 6685 24764
rect 6719 24761 6731 24795
rect 6946 24792 6952 24804
rect 6907 24764 6952 24792
rect 6673 24755 6731 24761
rect 6946 24752 6952 24764
rect 7004 24752 7010 24804
rect 7406 24792 7412 24804
rect 7367 24764 7412 24792
rect 7406 24752 7412 24764
rect 7464 24752 7470 24804
rect 11730 24792 11736 24804
rect 11691 24764 11736 24792
rect 11730 24752 11736 24764
rect 11788 24792 11794 24804
rect 11825 24795 11883 24801
rect 11825 24792 11837 24795
rect 11788 24764 11837 24792
rect 11788 24752 11794 24764
rect 11825 24761 11837 24764
rect 11871 24761 11883 24795
rect 11825 24755 11883 24761
rect 12101 24795 12159 24801
rect 12101 24761 12113 24795
rect 12147 24792 12159 24795
rect 12190 24792 12196 24804
rect 12147 24764 12196 24792
rect 12147 24761 12159 24764
rect 12101 24755 12159 24761
rect 1521 24727 1579 24733
rect 1521 24693 1533 24727
rect 1567 24724 1579 24727
rect 2162 24724 2168 24736
rect 1567 24696 2168 24724
rect 1567 24693 1579 24696
rect 1521 24687 1579 24693
rect 2162 24684 2168 24696
rect 2220 24684 2226 24736
rect 10442 24724 10448 24736
rect 10403 24696 10448 24724
rect 10442 24684 10448 24696
rect 10500 24684 10506 24736
rect 11362 24724 11368 24736
rect 11275 24696 11368 24724
rect 11362 24684 11368 24696
rect 11420 24724 11426 24736
rect 12116 24724 12144 24755
rect 12190 24752 12196 24764
rect 12248 24752 12254 24804
rect 12377 24795 12435 24801
rect 12377 24761 12389 24795
rect 12423 24792 12435 24795
rect 12466 24792 12472 24804
rect 12423 24764 12472 24792
rect 12423 24761 12435 24764
rect 12377 24755 12435 24761
rect 12466 24752 12472 24764
rect 12524 24752 12530 24804
rect 20838 24752 20844 24804
rect 20896 24792 20902 24804
rect 21669 24795 21727 24801
rect 21669 24792 21681 24795
rect 20896 24764 21681 24792
rect 20896 24752 20902 24764
rect 21669 24761 21681 24764
rect 21715 24792 21727 24795
rect 23230 24792 23236 24804
rect 21715 24764 23236 24792
rect 21715 24761 21727 24764
rect 21669 24755 21727 24761
rect 23230 24752 23236 24764
rect 23288 24792 23294 24804
rect 23506 24792 23512 24804
rect 23288 24764 23512 24792
rect 23288 24752 23294 24764
rect 23506 24752 23512 24764
rect 23564 24752 23570 24804
rect 23969 24795 24027 24801
rect 23969 24761 23981 24795
rect 24015 24792 24027 24795
rect 24058 24792 24064 24804
rect 24015 24764 24064 24792
rect 24015 24761 24027 24764
rect 23969 24755 24027 24761
rect 24058 24752 24064 24764
rect 24116 24792 24122 24804
rect 24153 24795 24211 24801
rect 24153 24792 24165 24795
rect 24116 24764 24165 24792
rect 24116 24752 24122 24764
rect 24153 24761 24165 24764
rect 24199 24761 24211 24795
rect 24153 24755 24211 24761
rect 11420 24696 12144 24724
rect 11420 24684 11426 24696
rect 4186 24656 4192 24668
rect 4147 24628 4192 24656
rect 4186 24616 4192 24628
rect 4244 24616 4250 24668
rect 5474 24616 5480 24668
rect 5532 24656 5538 24668
rect 6394 24656 6400 24668
rect 5532 24628 6400 24656
rect 5532 24616 5538 24628
rect 6394 24616 6400 24628
rect 6452 24616 6458 24668
rect 12558 24656 12564 24668
rect 12519 24628 12564 24656
rect 12558 24616 12564 24628
rect 12616 24616 12622 24668
rect 14861 24659 14919 24665
rect 14861 24625 14873 24659
rect 14907 24656 14919 24659
rect 14950 24656 14956 24668
rect 14907 24628 14956 24656
rect 14907 24625 14919 24628
rect 14861 24619 14919 24625
rect 14950 24616 14956 24628
rect 15008 24616 15014 24668
rect 18446 24656 18452 24668
rect 18407 24628 18452 24656
rect 18446 24616 18452 24628
rect 18504 24616 18510 24668
rect 18814 24656 18820 24668
rect 18775 24628 18820 24656
rect 18814 24616 18820 24628
rect 18872 24616 18878 24668
rect 19001 24659 19059 24665
rect 19001 24625 19013 24659
rect 19047 24656 19059 24659
rect 19642 24656 19648 24668
rect 19047 24628 19648 24656
rect 19047 24625 19059 24628
rect 19001 24619 19059 24625
rect 5566 24588 5572 24600
rect 5527 24560 5572 24588
rect 5566 24548 5572 24560
rect 5624 24548 5630 24600
rect 5658 24548 5664 24600
rect 5716 24588 5722 24600
rect 6486 24588 6492 24600
rect 5716 24560 5761 24588
rect 6447 24560 6492 24588
rect 5716 24548 5722 24560
rect 6486 24548 6492 24560
rect 6544 24548 6550 24600
rect 9246 24588 9252 24600
rect 9159 24560 9252 24588
rect 9246 24548 9252 24560
rect 9304 24588 9310 24600
rect 9433 24591 9491 24597
rect 9433 24588 9445 24591
rect 9304 24560 9445 24588
rect 9304 24548 9310 24560
rect 9433 24557 9445 24560
rect 9479 24588 9491 24591
rect 9982 24588 9988 24600
rect 9479 24560 9988 24588
rect 9479 24557 9491 24560
rect 9433 24551 9491 24557
rect 9982 24548 9988 24560
rect 10040 24548 10046 24600
rect 10537 24591 10595 24597
rect 10537 24557 10549 24591
rect 10583 24557 10595 24591
rect 15134 24588 15140 24600
rect 15095 24560 15140 24588
rect 10537 24551 10595 24557
rect 1058 24452 1064 24464
rect 1019 24424 1064 24452
rect 1058 24412 1064 24424
rect 1116 24412 1122 24464
rect 4278 24452 4284 24464
rect 4239 24424 4284 24452
rect 4278 24412 4284 24424
rect 4336 24412 4342 24464
rect 7498 24452 7504 24464
rect 7459 24424 7504 24452
rect 7498 24412 7504 24424
rect 7556 24412 7562 24464
rect 7777 24455 7835 24461
rect 7777 24421 7789 24455
rect 7823 24452 7835 24455
rect 7958 24452 7964 24464
rect 7823 24424 7964 24452
rect 7823 24421 7835 24424
rect 7777 24415 7835 24421
rect 7958 24412 7964 24424
rect 8016 24412 8022 24464
rect 9617 24455 9675 24461
rect 9617 24421 9629 24455
rect 9663 24452 9675 24455
rect 9798 24452 9804 24464
rect 9663 24424 9804 24452
rect 9663 24421 9675 24424
rect 9617 24415 9675 24421
rect 9798 24412 9804 24424
rect 9856 24412 9862 24464
rect 10552 24452 10580 24551
rect 15134 24548 15140 24560
rect 15192 24548 15198 24600
rect 17986 24548 17992 24600
rect 18044 24588 18050 24600
rect 18357 24591 18415 24597
rect 18357 24588 18369 24591
rect 18044 24560 18369 24588
rect 18044 24548 18050 24560
rect 18357 24557 18369 24560
rect 18403 24557 18415 24591
rect 18357 24551 18415 24557
rect 18722 24548 18728 24600
rect 18780 24588 18786 24600
rect 19016 24588 19044 24619
rect 19642 24616 19648 24628
rect 19700 24616 19706 24668
rect 21025 24659 21083 24665
rect 21025 24625 21037 24659
rect 21071 24656 21083 24659
rect 21482 24656 21488 24668
rect 21071 24628 21488 24656
rect 21071 24625 21083 24628
rect 21025 24619 21083 24625
rect 21482 24616 21488 24628
rect 21540 24616 21546 24668
rect 22589 24659 22647 24665
rect 22589 24625 22601 24659
rect 22635 24656 22647 24659
rect 22862 24656 22868 24668
rect 22635 24628 22868 24656
rect 22635 24625 22647 24628
rect 22589 24619 22647 24625
rect 22862 24616 22868 24628
rect 22920 24616 22926 24668
rect 24426 24656 24432 24668
rect 24387 24628 24432 24656
rect 24426 24616 24432 24628
rect 24484 24616 24490 24668
rect 18780 24560 19044 24588
rect 18780 24548 18786 24560
rect 20562 24548 20568 24600
rect 20620 24588 20626 24600
rect 20933 24591 20991 24597
rect 20933 24588 20945 24591
rect 20620 24560 20945 24588
rect 20620 24548 20626 24560
rect 20933 24557 20945 24560
rect 20979 24557 20991 24591
rect 24702 24588 24708 24600
rect 24663 24560 24708 24588
rect 20933 24551 20991 24557
rect 24702 24548 24708 24560
rect 24760 24548 24766 24600
rect 20473 24523 20531 24529
rect 20473 24489 20485 24523
rect 20519 24520 20531 24523
rect 20746 24520 20752 24532
rect 20519 24492 20752 24520
rect 20519 24489 20531 24492
rect 20473 24483 20531 24489
rect 20746 24480 20752 24492
rect 20804 24480 20810 24532
rect 11454 24452 11460 24464
rect 10552 24424 11460 24452
rect 11454 24412 11460 24424
rect 11512 24412 11518 24464
rect 14677 24455 14735 24461
rect 14677 24421 14689 24455
rect 14723 24452 14735 24455
rect 16422 24452 16428 24464
rect 14723 24424 16428 24452
rect 14723 24421 14735 24424
rect 14677 24415 14735 24421
rect 16422 24412 16428 24424
rect 16480 24412 16486 24464
rect 17342 24452 17348 24464
rect 17303 24424 17348 24452
rect 17342 24412 17348 24424
rect 17400 24412 17406 24464
rect 17894 24452 17900 24464
rect 17807 24424 17900 24452
rect 17894 24412 17900 24424
rect 17952 24452 17958 24464
rect 18538 24452 18544 24464
rect 17952 24424 18544 24452
rect 17952 24412 17958 24424
rect 18538 24412 18544 24424
rect 18596 24412 18602 24464
rect 20654 24452 20660 24464
rect 20615 24424 20660 24452
rect 20654 24412 20660 24424
rect 20712 24412 20718 24464
rect 21022 24412 21028 24464
rect 21080 24452 21086 24464
rect 21209 24455 21267 24461
rect 21209 24452 21221 24455
rect 21080 24424 21221 24452
rect 21080 24412 21086 24424
rect 21209 24421 21221 24424
rect 21255 24452 21267 24455
rect 21390 24452 21396 24464
rect 21255 24424 21396 24452
rect 21255 24421 21267 24424
rect 21209 24415 21267 24421
rect 21390 24412 21396 24424
rect 21448 24412 21454 24464
rect 22402 24452 22408 24464
rect 22363 24424 22408 24452
rect 22402 24412 22408 24424
rect 22460 24412 22466 24464
rect 400 24362 27264 24384
rect 400 24310 3510 24362
rect 3562 24310 3574 24362
rect 3626 24310 3638 24362
rect 3690 24310 3702 24362
rect 3754 24310 3766 24362
rect 3818 24310 27264 24362
rect 400 24288 27264 24310
rect 2993 24251 3051 24257
rect 2993 24217 3005 24251
rect 3039 24248 3051 24251
rect 3453 24251 3511 24257
rect 3453 24248 3465 24251
rect 3039 24220 3465 24248
rect 3039 24217 3051 24220
rect 2993 24211 3051 24217
rect 3453 24217 3465 24220
rect 3499 24248 3511 24251
rect 3910 24248 3916 24260
rect 3499 24220 3916 24248
rect 3499 24217 3511 24220
rect 3453 24211 3511 24217
rect 3910 24208 3916 24220
rect 3968 24208 3974 24260
rect 4278 24248 4284 24260
rect 4239 24220 4284 24248
rect 4278 24208 4284 24220
rect 4336 24208 4342 24260
rect 5658 24208 5664 24260
rect 5716 24248 5722 24260
rect 6121 24251 6179 24257
rect 6121 24248 6133 24251
rect 5716 24220 6133 24248
rect 5716 24208 5722 24220
rect 6121 24217 6133 24220
rect 6167 24217 6179 24251
rect 6121 24211 6179 24217
rect 6857 24251 6915 24257
rect 6857 24217 6869 24251
rect 6903 24248 6915 24251
rect 6946 24248 6952 24260
rect 6903 24220 6952 24248
rect 6903 24217 6915 24220
rect 6857 24211 6915 24217
rect 6946 24208 6952 24220
rect 7004 24208 7010 24260
rect 7041 24251 7099 24257
rect 7041 24217 7053 24251
rect 7087 24248 7099 24251
rect 7498 24248 7504 24260
rect 7087 24220 7504 24248
rect 7087 24217 7099 24220
rect 7041 24211 7099 24217
rect 7498 24208 7504 24220
rect 7556 24208 7562 24260
rect 9982 24248 9988 24260
rect 9943 24220 9988 24248
rect 9982 24208 9988 24220
rect 10040 24208 10046 24260
rect 10261 24251 10319 24257
rect 10261 24217 10273 24251
rect 10307 24248 10319 24251
rect 11454 24248 11460 24260
rect 10307 24220 11460 24248
rect 10307 24217 10319 24220
rect 10261 24211 10319 24217
rect 11454 24208 11460 24220
rect 11512 24248 11518 24260
rect 11733 24251 11791 24257
rect 11733 24248 11745 24251
rect 11512 24220 11745 24248
rect 11512 24208 11518 24220
rect 11733 24217 11745 24220
rect 11779 24217 11791 24251
rect 12466 24248 12472 24260
rect 12427 24220 12472 24248
rect 11733 24211 11791 24217
rect 12466 24208 12472 24220
rect 12524 24208 12530 24260
rect 12558 24208 12564 24260
rect 12616 24248 12622 24260
rect 18446 24248 18452 24260
rect 12616 24220 12661 24248
rect 18407 24220 18452 24248
rect 12616 24208 12622 24220
rect 18446 24208 18452 24220
rect 18504 24208 18510 24260
rect 18538 24208 18544 24260
rect 18596 24248 18602 24260
rect 18596 24220 18641 24248
rect 18596 24208 18602 24220
rect 21482 24208 21488 24260
rect 21540 24248 21546 24260
rect 22589 24251 22647 24257
rect 22589 24248 22601 24251
rect 21540 24220 22601 24248
rect 21540 24208 21546 24220
rect 22589 24217 22601 24220
rect 22635 24248 22647 24251
rect 22862 24248 22868 24260
rect 22635 24220 22868 24248
rect 22635 24217 22647 24220
rect 22589 24211 22647 24217
rect 22862 24208 22868 24220
rect 22920 24208 22926 24260
rect 23598 24248 23604 24260
rect 23559 24220 23604 24248
rect 23598 24208 23604 24220
rect 23656 24248 23662 24260
rect 23656 24220 24380 24248
rect 23656 24208 23662 24220
rect 874 24140 880 24192
rect 932 24180 938 24192
rect 4186 24180 4192 24192
rect 932 24152 1932 24180
rect 4147 24152 4192 24180
rect 932 24140 938 24152
rect 1058 24112 1064 24124
rect 1019 24084 1064 24112
rect 1058 24072 1064 24084
rect 1116 24072 1122 24124
rect 1904 24121 1932 24152
rect 4186 24140 4192 24152
rect 4244 24140 4250 24192
rect 5566 24140 5572 24192
rect 5624 24180 5630 24192
rect 5845 24183 5903 24189
rect 5845 24180 5857 24183
rect 5624 24152 5857 24180
rect 5624 24140 5630 24152
rect 5845 24149 5857 24152
rect 5891 24149 5903 24183
rect 5845 24143 5903 24149
rect 7225 24183 7283 24189
rect 7225 24149 7237 24183
rect 7271 24180 7283 24183
rect 7406 24180 7412 24192
rect 7271 24152 7412 24180
rect 7271 24149 7283 24152
rect 7225 24143 7283 24149
rect 7406 24140 7412 24152
rect 7464 24140 7470 24192
rect 10442 24180 10448 24192
rect 10403 24152 10448 24180
rect 10442 24140 10448 24152
rect 10500 24140 10506 24192
rect 11362 24180 11368 24192
rect 11323 24152 11368 24180
rect 11362 24140 11368 24152
rect 11420 24140 11426 24192
rect 18265 24183 18323 24189
rect 18265 24149 18277 24183
rect 18311 24180 18323 24183
rect 18722 24180 18728 24192
rect 18311 24152 18728 24180
rect 18311 24149 18323 24152
rect 18265 24143 18323 24149
rect 18722 24140 18728 24152
rect 18780 24140 18786 24192
rect 20381 24183 20439 24189
rect 20381 24180 20393 24183
rect 18832 24152 20393 24180
rect 18832 24124 18860 24152
rect 20381 24149 20393 24152
rect 20427 24180 20439 24183
rect 20470 24180 20476 24192
rect 20427 24152 20476 24180
rect 20427 24149 20439 24152
rect 20381 24143 20439 24149
rect 20470 24140 20476 24152
rect 20528 24140 20534 24192
rect 20654 24180 20660 24192
rect 20615 24152 20660 24180
rect 20654 24140 20660 24152
rect 20712 24140 20718 24192
rect 22402 24180 22408 24192
rect 22363 24152 22408 24180
rect 22402 24140 22408 24152
rect 22460 24140 22466 24192
rect 1889 24115 1947 24121
rect 1889 24081 1901 24115
rect 1935 24081 1947 24115
rect 1889 24075 1947 24081
rect 5753 24115 5811 24121
rect 5753 24081 5765 24115
rect 5799 24112 5811 24115
rect 6486 24112 6492 24124
rect 5799 24084 6492 24112
rect 5799 24081 5811 24084
rect 5753 24075 5811 24081
rect 6486 24072 6492 24084
rect 6544 24072 6550 24124
rect 14125 24115 14183 24121
rect 14125 24081 14137 24115
rect 14171 24112 14183 24115
rect 15134 24112 15140 24124
rect 14171 24084 15140 24112
rect 14171 24081 14183 24084
rect 14125 24075 14183 24081
rect 15134 24072 15140 24084
rect 15192 24072 15198 24124
rect 16422 24112 16428 24124
rect 16383 24084 16428 24112
rect 16422 24072 16428 24084
rect 16480 24072 16486 24124
rect 17897 24115 17955 24121
rect 17897 24081 17909 24115
rect 17943 24112 17955 24115
rect 18814 24112 18820 24124
rect 17943 24084 18820 24112
rect 17943 24081 17955 24084
rect 17897 24075 17955 24081
rect 18814 24072 18820 24084
rect 18872 24072 18878 24124
rect 20289 24115 20347 24121
rect 20289 24081 20301 24115
rect 20335 24112 20347 24115
rect 20746 24112 20752 24124
rect 20335 24084 20752 24112
rect 20335 24081 20347 24084
rect 20289 24075 20347 24081
rect 20746 24072 20752 24084
rect 20804 24112 20810 24124
rect 20804 24084 21252 24112
rect 20804 24072 20810 24084
rect 782 24004 788 24056
rect 840 24044 846 24056
rect 969 24047 1027 24053
rect 969 24044 981 24047
rect 840 24016 981 24044
rect 840 24004 846 24016
rect 969 24013 981 24016
rect 1015 24013 1027 24047
rect 969 24007 1027 24013
rect 1518 24004 1524 24056
rect 1576 24044 1582 24056
rect 1797 24047 1855 24053
rect 1797 24044 1809 24047
rect 1576 24016 1809 24044
rect 1576 24004 1582 24016
rect 1797 24013 1809 24016
rect 1843 24044 1855 24047
rect 5474 24044 5480 24056
rect 1843 24016 5480 24044
rect 1843 24013 1855 24016
rect 1797 24007 1855 24013
rect 5474 24004 5480 24016
rect 5532 24004 5538 24056
rect 7406 24044 7412 24056
rect 7319 24016 7412 24044
rect 7406 24004 7412 24016
rect 7464 24044 7470 24056
rect 7501 24047 7559 24053
rect 7501 24044 7513 24047
rect 7464 24016 7513 24044
rect 7464 24004 7470 24016
rect 7501 24013 7513 24016
rect 7547 24013 7559 24047
rect 8418 24044 8424 24056
rect 8379 24016 8424 24044
rect 7501 24007 7559 24013
rect 8418 24004 8424 24016
rect 8476 24004 8482 24056
rect 13941 24047 13999 24053
rect 13941 24013 13953 24047
rect 13987 24044 13999 24047
rect 14398 24044 14404 24056
rect 13987 24016 14404 24044
rect 13987 24013 13999 24016
rect 13941 24007 13999 24013
rect 14398 24004 14404 24016
rect 14456 24004 14462 24056
rect 20105 24047 20163 24053
rect 20105 24013 20117 24047
rect 20151 24044 20163 24047
rect 20565 24047 20623 24053
rect 20565 24044 20577 24047
rect 20151 24016 20577 24044
rect 20151 24013 20163 24016
rect 20105 24007 20163 24013
rect 20565 24013 20577 24016
rect 20611 24044 20623 24047
rect 21022 24044 21028 24056
rect 20611 24016 21028 24044
rect 20611 24013 20623 24016
rect 20565 24007 20623 24013
rect 21022 24004 21028 24016
rect 21080 24004 21086 24056
rect 21117 24047 21175 24053
rect 21117 24013 21129 24047
rect 21163 24013 21175 24047
rect 21224 24044 21252 24084
rect 21577 24047 21635 24053
rect 21577 24044 21589 24047
rect 21224 24016 21589 24044
rect 21117 24007 21175 24013
rect 21577 24013 21589 24016
rect 21623 24044 21635 24047
rect 22420 24044 22448 24140
rect 21623 24016 22448 24044
rect 21623 24013 21635 24016
rect 21577 24007 21635 24013
rect 693 23979 751 23985
rect 693 23945 705 23979
rect 739 23976 751 23979
rect 1536 23976 1564 24004
rect 739 23948 1564 23976
rect 739 23945 751 23948
rect 693 23939 751 23945
rect 2162 23936 2168 23988
rect 2220 23976 2226 23988
rect 2901 23979 2959 23985
rect 2901 23976 2913 23979
rect 2220 23948 2913 23976
rect 2220 23936 2226 23948
rect 2901 23945 2913 23948
rect 2947 23976 2959 23979
rect 3177 23979 3235 23985
rect 3177 23976 3189 23979
rect 2947 23948 3189 23976
rect 2947 23945 2959 23948
rect 2901 23939 2959 23945
rect 3177 23945 3189 23948
rect 3223 23945 3235 23979
rect 9062 23976 9068 23988
rect 9023 23948 9068 23976
rect 3177 23939 3235 23945
rect 9062 23936 9068 23948
rect 9120 23936 9126 23988
rect 14677 23979 14735 23985
rect 14677 23945 14689 23979
rect 14723 23945 14735 23979
rect 14677 23939 14735 23945
rect 14309 23911 14367 23917
rect 14309 23877 14321 23911
rect 14355 23908 14367 23911
rect 14692 23908 14720 23939
rect 15134 23936 15140 23988
rect 15192 23936 15198 23988
rect 20470 23936 20476 23988
rect 20528 23976 20534 23988
rect 21132 23976 21160 24007
rect 24058 24004 24064 24056
rect 24116 24044 24122 24056
rect 24245 24047 24303 24053
rect 24245 24044 24257 24047
rect 24116 24016 24257 24044
rect 24116 24004 24122 24016
rect 24245 24013 24257 24016
rect 24291 24013 24303 24047
rect 24352 24044 24380 24220
rect 24797 24047 24855 24053
rect 24797 24044 24809 24047
rect 24352 24016 24809 24044
rect 24245 24007 24303 24013
rect 24797 24013 24809 24016
rect 24843 24013 24855 24047
rect 24797 24007 24855 24013
rect 20528 23948 21160 23976
rect 20528 23936 20534 23948
rect 23414 23936 23420 23988
rect 23472 23976 23478 23988
rect 23877 23979 23935 23985
rect 23877 23976 23889 23979
rect 23472 23948 23889 23976
rect 23472 23936 23478 23948
rect 23877 23945 23889 23948
rect 23923 23976 23935 23979
rect 23923 23948 25208 23976
rect 23923 23945 23935 23948
rect 23877 23939 23935 23945
rect 16514 23908 16520 23920
rect 14355 23880 16520 23908
rect 14355 23877 14367 23880
rect 14309 23871 14367 23877
rect 16514 23868 16520 23880
rect 16572 23868 16578 23920
rect 16882 23868 16888 23920
rect 16940 23908 16946 23920
rect 17986 23908 17992 23920
rect 16940 23880 17992 23908
rect 16940 23868 16946 23880
rect 17986 23868 17992 23880
rect 18044 23868 18050 23920
rect 21390 23868 21396 23920
rect 21448 23908 21454 23920
rect 21761 23911 21819 23917
rect 21761 23908 21773 23911
rect 21448 23880 21773 23908
rect 21448 23868 21454 23880
rect 21761 23877 21773 23880
rect 21807 23877 21819 23911
rect 21761 23871 21819 23877
rect 24061 23911 24119 23917
rect 24061 23877 24073 23911
rect 24107 23908 24119 23911
rect 24426 23908 24432 23920
rect 24107 23880 24432 23908
rect 24107 23877 24119 23880
rect 24061 23871 24119 23877
rect 24426 23868 24432 23880
rect 24484 23868 24490 23920
rect 400 23818 27264 23840
rect 400 23766 18870 23818
rect 18922 23766 18934 23818
rect 18986 23766 18998 23818
rect 19050 23766 19062 23818
rect 19114 23766 19126 23818
rect 19178 23766 27264 23818
rect 400 23744 27264 23766
rect 14950 23704 14956 23716
rect 14911 23676 14956 23704
rect 14950 23664 14956 23676
rect 15008 23664 15014 23716
rect 15134 23704 15140 23716
rect 15095 23676 15140 23704
rect 15134 23664 15140 23676
rect 15192 23664 15198 23716
rect 18354 23704 18360 23716
rect 18315 23676 18360 23704
rect 18354 23664 18360 23676
rect 18412 23664 18418 23716
rect 21482 23704 21488 23716
rect 21443 23676 21488 23704
rect 21482 23664 21488 23676
rect 21540 23664 21546 23716
rect 24521 23707 24579 23713
rect 24521 23673 24533 23707
rect 24567 23704 24579 23707
rect 24702 23704 24708 23716
rect 24567 23676 24708 23704
rect 24567 23673 24579 23676
rect 24521 23667 24579 23673
rect 24702 23664 24708 23676
rect 24760 23664 24766 23716
rect 7498 23596 7504 23648
rect 7556 23636 7562 23648
rect 8053 23639 8111 23645
rect 8053 23636 8065 23639
rect 7556 23608 8065 23636
rect 7556 23596 7562 23608
rect 8053 23605 8065 23608
rect 8099 23605 8111 23639
rect 8053 23599 8111 23605
rect 12466 23596 12472 23648
rect 12524 23636 12530 23648
rect 16238 23636 16244 23648
rect 12524 23608 13340 23636
rect 12524 23596 12530 23608
rect 1058 23528 1064 23580
rect 1116 23568 1122 23580
rect 1245 23571 1303 23577
rect 1245 23568 1257 23571
rect 1116 23540 1257 23568
rect 1116 23528 1122 23540
rect 1245 23537 1257 23540
rect 1291 23537 1303 23571
rect 1245 23531 1303 23537
rect 1705 23571 1763 23577
rect 1705 23537 1717 23571
rect 1751 23568 1763 23571
rect 1886 23568 1892 23580
rect 1751 23540 1892 23568
rect 1751 23537 1763 23540
rect 1705 23531 1763 23537
rect 1886 23528 1892 23540
rect 1944 23528 1950 23580
rect 4186 23568 4192 23580
rect 4147 23540 4192 23568
rect 4186 23528 4192 23540
rect 4244 23528 4250 23580
rect 4278 23528 4284 23580
rect 4336 23568 4342 23580
rect 13312 23577 13340 23608
rect 14186 23608 16244 23636
rect 5109 23571 5167 23577
rect 5109 23568 5121 23571
rect 4336 23540 5121 23568
rect 4336 23528 4342 23540
rect 5109 23537 5121 23540
rect 5155 23537 5167 23571
rect 5109 23531 5167 23537
rect 13297 23571 13355 23577
rect 13297 23537 13309 23571
rect 13343 23537 13355 23571
rect 13297 23531 13355 23537
rect 13386 23528 13392 23580
rect 13444 23568 13450 23580
rect 14186 23568 14214 23608
rect 16238 23596 16244 23608
rect 16296 23596 16302 23648
rect 13444 23540 14214 23568
rect 13444 23528 13450 23540
rect 15962 23528 15968 23580
rect 16020 23568 16026 23580
rect 16057 23571 16115 23577
rect 16057 23568 16069 23571
rect 16020 23540 16069 23568
rect 16020 23528 16026 23540
rect 16057 23537 16069 23540
rect 16103 23568 16115 23571
rect 16422 23568 16428 23580
rect 16103 23540 16428 23568
rect 16103 23537 16115 23540
rect 16057 23531 16115 23537
rect 16422 23528 16428 23540
rect 16480 23528 16486 23580
rect 18078 23568 18084 23580
rect 18039 23540 18084 23568
rect 18078 23528 18084 23540
rect 18136 23528 18142 23580
rect 18630 23568 18636 23580
rect 18591 23540 18636 23568
rect 18630 23528 18636 23540
rect 18688 23528 18694 23580
rect 20562 23568 20568 23580
rect 20523 23540 20568 23568
rect 20562 23528 20568 23540
rect 20620 23528 20626 23580
rect 20654 23528 20660 23580
rect 20712 23568 20718 23580
rect 20712 23540 20757 23568
rect 20712 23528 20718 23540
rect 1794 23500 1800 23512
rect 1755 23472 1800 23500
rect 1794 23460 1800 23472
rect 1852 23460 1858 23512
rect 5750 23500 5756 23512
rect 5711 23472 5756 23500
rect 5750 23460 5756 23472
rect 5808 23460 5814 23512
rect 7406 23460 7412 23512
rect 7464 23500 7470 23512
rect 7501 23503 7559 23509
rect 7501 23500 7513 23503
rect 7464 23472 7513 23500
rect 7464 23460 7470 23472
rect 7501 23469 7513 23472
rect 7547 23469 7559 23503
rect 7501 23463 7559 23469
rect 12282 23460 12288 23512
rect 12340 23500 12346 23512
rect 12469 23503 12527 23509
rect 12469 23500 12481 23503
rect 12340 23472 12481 23500
rect 12340 23460 12346 23472
rect 12469 23469 12481 23472
rect 12515 23469 12527 23503
rect 12469 23463 12527 23469
rect 12558 23460 12564 23512
rect 12616 23500 12622 23512
rect 20580 23500 20608 23528
rect 20930 23500 20936 23512
rect 12616 23472 12661 23500
rect 20580 23472 20936 23500
rect 12616 23460 12622 23472
rect 20930 23460 20936 23472
rect 20988 23500 20994 23512
rect 21209 23503 21267 23509
rect 21209 23500 21221 23503
rect 20988 23472 21221 23500
rect 20988 23460 20994 23472
rect 21209 23469 21221 23472
rect 21255 23469 21267 23503
rect 21209 23463 21267 23469
rect 7958 23432 7964 23444
rect 7919 23404 7964 23432
rect 7958 23392 7964 23404
rect 8016 23392 8022 23444
rect 782 23324 788 23376
rect 840 23364 846 23376
rect 969 23367 1027 23373
rect 969 23364 981 23367
rect 840 23336 981 23364
rect 840 23324 846 23336
rect 969 23333 981 23336
rect 1015 23364 1027 23367
rect 1150 23364 1156 23376
rect 1015 23336 1156 23364
rect 1015 23333 1027 23336
rect 969 23327 1027 23333
rect 1150 23324 1156 23336
rect 1208 23324 1214 23376
rect 1978 23364 1984 23376
rect 1939 23336 1984 23364
rect 1978 23324 1984 23336
rect 2036 23324 2042 23376
rect 16333 23367 16391 23373
rect 16333 23333 16345 23367
rect 16379 23364 16391 23367
rect 16698 23364 16704 23376
rect 16379 23336 16704 23364
rect 16379 23333 16391 23336
rect 16333 23327 16391 23333
rect 16698 23324 16704 23336
rect 16756 23324 16762 23376
rect 20838 23364 20844 23376
rect 20799 23336 20844 23364
rect 20838 23324 20844 23336
rect 20896 23324 20902 23376
rect 24150 23364 24156 23376
rect 24111 23336 24156 23364
rect 24150 23324 24156 23336
rect 24208 23324 24214 23376
rect 400 23274 27264 23296
rect 400 23222 3510 23274
rect 3562 23222 3574 23274
rect 3626 23222 3638 23274
rect 3690 23222 3702 23274
rect 3754 23222 3766 23274
rect 3818 23222 27264 23274
rect 400 23200 27264 23222
rect 877 23163 935 23169
rect 877 23129 889 23163
rect 923 23160 935 23163
rect 1058 23160 1064 23172
rect 923 23132 1064 23160
rect 923 23129 935 23132
rect 877 23123 935 23129
rect 1058 23120 1064 23132
rect 1116 23120 1122 23172
rect 4186 23160 4192 23172
rect 4147 23132 4192 23160
rect 4186 23120 4192 23132
rect 4244 23160 4250 23172
rect 5385 23163 5443 23169
rect 5385 23160 5397 23163
rect 4244 23132 5397 23160
rect 4244 23120 4250 23132
rect 1794 23052 1800 23104
rect 1852 23092 1858 23104
rect 2901 23095 2959 23101
rect 2901 23092 2913 23095
rect 1852 23064 2913 23092
rect 1852 23052 1858 23064
rect 2901 23061 2913 23064
rect 2947 23092 2959 23095
rect 3177 23095 3235 23101
rect 3177 23092 3189 23095
rect 2947 23064 3189 23092
rect 2947 23061 2959 23064
rect 2901 23055 2959 23061
rect 3177 23061 3189 23064
rect 3223 23061 3235 23095
rect 3177 23055 3235 23061
rect 3913 23095 3971 23101
rect 3913 23061 3925 23095
rect 3959 23092 3971 23095
rect 4278 23092 4284 23104
rect 3959 23064 4284 23092
rect 3959 23061 3971 23064
rect 3913 23055 3971 23061
rect 4278 23052 4284 23064
rect 4336 23052 4342 23104
rect 4664 23033 4692 23132
rect 5385 23129 5397 23132
rect 5431 23160 5443 23163
rect 5658 23160 5664 23172
rect 5431 23132 5664 23160
rect 5431 23129 5443 23132
rect 5385 23123 5443 23129
rect 5658 23120 5664 23132
rect 5716 23120 5722 23172
rect 7498 23120 7504 23172
rect 7556 23160 7562 23172
rect 7685 23163 7743 23169
rect 7685 23160 7697 23163
rect 7556 23132 7697 23160
rect 7556 23120 7562 23132
rect 7685 23129 7697 23132
rect 7731 23129 7743 23163
rect 7685 23123 7743 23129
rect 13297 23163 13355 23169
rect 13297 23129 13309 23163
rect 13343 23160 13355 23163
rect 13386 23160 13392 23172
rect 13343 23132 13392 23160
rect 13343 23129 13355 23132
rect 13297 23123 13355 23129
rect 13386 23120 13392 23132
rect 13444 23120 13450 23172
rect 16698 23160 16704 23172
rect 16659 23132 16704 23160
rect 16698 23120 16704 23132
rect 16756 23120 16762 23172
rect 18354 23160 18360 23172
rect 18315 23132 18360 23160
rect 18354 23120 18360 23132
rect 18412 23120 18418 23172
rect 18722 23120 18728 23172
rect 18780 23160 18786 23172
rect 18817 23163 18875 23169
rect 18817 23160 18829 23163
rect 18780 23132 18829 23160
rect 18780 23120 18786 23132
rect 18817 23129 18829 23132
rect 18863 23160 18875 23163
rect 19369 23163 19427 23169
rect 19369 23160 19381 23163
rect 18863 23132 19381 23160
rect 18863 23129 18875 23132
rect 18817 23123 18875 23129
rect 19369 23129 19381 23132
rect 19415 23160 19427 23163
rect 20565 23163 20623 23169
rect 20565 23160 20577 23163
rect 19415 23132 20577 23160
rect 19415 23129 19427 23132
rect 19369 23123 19427 23129
rect 20565 23129 20577 23132
rect 20611 23160 20623 23163
rect 20654 23160 20660 23172
rect 20611 23132 20660 23160
rect 20611 23129 20623 23132
rect 20565 23123 20623 23129
rect 20654 23120 20660 23132
rect 20712 23120 20718 23172
rect 20930 23160 20936 23172
rect 20891 23132 20936 23160
rect 20930 23120 20936 23132
rect 20988 23120 20994 23172
rect 9525 23095 9583 23101
rect 9525 23061 9537 23095
rect 9571 23092 9583 23095
rect 9798 23092 9804 23104
rect 9571 23064 9804 23092
rect 9571 23061 9583 23064
rect 9525 23055 9583 23061
rect 9798 23052 9804 23064
rect 9856 23052 9862 23104
rect 4649 23027 4707 23033
rect 4649 22993 4661 23027
rect 4695 22993 4707 23027
rect 4649 22987 4707 22993
rect 7406 22984 7412 23036
rect 7464 23024 7470 23036
rect 7501 23027 7559 23033
rect 7501 23024 7513 23027
rect 7464 22996 7513 23024
rect 7464 22984 7470 22996
rect 7501 22993 7513 22996
rect 7547 22993 7559 23027
rect 7501 22987 7559 22993
rect 11822 22984 11828 23036
rect 11880 23024 11886 23036
rect 12377 23027 12435 23033
rect 12377 23024 12389 23027
rect 11880 22996 12389 23024
rect 11880 22984 11886 22996
rect 12377 22993 12389 22996
rect 12423 22993 12435 23027
rect 13389 23027 13447 23033
rect 13389 23024 13401 23027
rect 12377 22987 12435 22993
rect 12576 22996 13401 23024
rect 12576 22968 12604 22996
rect 13389 22993 13401 22996
rect 13435 22993 13447 23027
rect 24150 23024 24156 23036
rect 13389 22987 13447 22993
rect 23846 22996 24156 23024
rect 1058 22916 1064 22968
rect 1116 22956 1122 22968
rect 1153 22959 1211 22965
rect 1153 22956 1165 22959
rect 1116 22928 1165 22956
rect 1116 22916 1122 22928
rect 1153 22925 1165 22928
rect 1199 22925 1211 22959
rect 1153 22919 1211 22925
rect 1978 22916 1984 22968
rect 2036 22956 2042 22968
rect 2073 22959 2131 22965
rect 2073 22956 2085 22959
rect 2036 22928 2085 22956
rect 2036 22916 2042 22928
rect 2073 22925 2085 22928
rect 2119 22956 2131 22959
rect 3085 22959 3143 22965
rect 3085 22956 3097 22959
rect 2119 22928 3097 22956
rect 2119 22925 2131 22928
rect 2073 22919 2131 22925
rect 3085 22925 3097 22928
rect 3131 22956 3143 22959
rect 3361 22959 3419 22965
rect 3361 22956 3373 22959
rect 3131 22928 3373 22956
rect 3131 22925 3143 22928
rect 3085 22919 3143 22925
rect 3361 22925 3373 22928
rect 3407 22925 3419 22959
rect 3361 22919 3419 22925
rect 4097 22959 4155 22965
rect 4097 22925 4109 22959
rect 4143 22956 4155 22959
rect 4557 22959 4615 22965
rect 4557 22956 4569 22959
rect 4143 22928 4569 22956
rect 4143 22925 4155 22928
rect 4097 22919 4155 22925
rect 4557 22925 4569 22928
rect 4603 22956 4615 22959
rect 5109 22959 5167 22965
rect 5109 22956 5121 22959
rect 4603 22928 5121 22956
rect 4603 22925 4615 22928
rect 4557 22919 4615 22925
rect 5109 22925 5121 22928
rect 5155 22956 5167 22959
rect 5750 22956 5756 22968
rect 5155 22928 5756 22956
rect 5155 22925 5167 22928
rect 5109 22919 5167 22925
rect 5750 22916 5756 22928
rect 5808 22916 5814 22968
rect 7958 22956 7964 22968
rect 7871 22928 7964 22956
rect 7958 22916 7964 22928
rect 8016 22956 8022 22968
rect 9062 22956 9068 22968
rect 8016 22928 9068 22956
rect 8016 22916 8022 22928
rect 9062 22916 9068 22928
rect 9120 22956 9126 22968
rect 10445 22959 10503 22965
rect 10445 22956 10457 22959
rect 9120 22928 10457 22956
rect 9120 22916 9126 22928
rect 10445 22925 10457 22928
rect 10491 22956 10503 22959
rect 10721 22959 10779 22965
rect 10721 22956 10733 22959
rect 10491 22928 10733 22956
rect 10491 22925 10503 22928
rect 10445 22919 10503 22925
rect 10721 22925 10733 22928
rect 10767 22925 10779 22959
rect 10721 22919 10779 22925
rect 12006 22916 12012 22968
rect 12064 22956 12070 22968
rect 12558 22956 12564 22968
rect 12064 22928 12564 22956
rect 12064 22916 12070 22928
rect 12558 22916 12564 22928
rect 12616 22916 12622 22968
rect 13021 22959 13079 22965
rect 13021 22925 13033 22959
rect 13067 22956 13079 22959
rect 13478 22956 13484 22968
rect 13067 22928 13484 22956
rect 13067 22925 13079 22928
rect 13021 22919 13079 22925
rect 13478 22916 13484 22928
rect 13536 22956 13542 22968
rect 13573 22959 13631 22965
rect 13573 22956 13585 22959
rect 13536 22928 13585 22956
rect 13536 22916 13542 22928
rect 13573 22925 13585 22928
rect 13619 22925 13631 22959
rect 13573 22919 13631 22925
rect 15870 22916 15876 22968
rect 15928 22956 15934 22968
rect 16057 22959 16115 22965
rect 16057 22956 16069 22959
rect 15928 22928 16069 22956
rect 15928 22916 15934 22928
rect 16057 22925 16069 22928
rect 16103 22956 16115 22959
rect 16146 22956 16152 22968
rect 16103 22928 16152 22956
rect 16103 22925 16115 22928
rect 16057 22919 16115 22925
rect 16146 22916 16152 22928
rect 16204 22956 16210 22968
rect 16885 22959 16943 22965
rect 16885 22956 16897 22959
rect 16204 22928 16897 22956
rect 16204 22916 16210 22928
rect 16885 22925 16897 22928
rect 16931 22956 16943 22959
rect 17897 22959 17955 22965
rect 17897 22956 17909 22959
rect 16931 22928 17909 22956
rect 16931 22925 16943 22928
rect 16885 22919 16943 22925
rect 17897 22925 17909 22928
rect 17943 22956 17955 22959
rect 18078 22956 18084 22968
rect 17943 22928 18084 22956
rect 17943 22925 17955 22928
rect 17897 22919 17955 22925
rect 18078 22916 18084 22928
rect 18136 22956 18142 22968
rect 18538 22956 18544 22968
rect 18136 22928 18544 22956
rect 18136 22916 18142 22928
rect 18538 22916 18544 22928
rect 18596 22916 18602 22968
rect 18630 22916 18636 22968
rect 18688 22956 18694 22968
rect 18688 22928 18781 22956
rect 18688 22916 18694 22928
rect 23230 22916 23236 22968
rect 23288 22956 23294 22968
rect 23846 22956 23874 22996
rect 24150 22984 24156 22996
rect 24208 22984 24214 23036
rect 24426 22984 24432 23036
rect 24484 23024 24490 23036
rect 26177 23027 26235 23033
rect 26177 23024 26189 23027
rect 24484 22996 26189 23024
rect 24484 22984 24490 22996
rect 26177 22993 26189 22996
rect 26223 22993 26235 23027
rect 26177 22987 26235 22993
rect 23288 22928 23874 22956
rect 23288 22916 23294 22928
rect 1886 22888 1892 22900
rect 1847 22860 1892 22888
rect 1886 22848 1892 22860
rect 1944 22848 1950 22900
rect 5198 22848 5204 22900
rect 5256 22888 5262 22900
rect 5477 22891 5535 22897
rect 5477 22888 5489 22891
rect 5256 22860 5489 22888
rect 5256 22848 5262 22860
rect 5477 22857 5489 22860
rect 5523 22857 5535 22891
rect 5477 22851 5535 22857
rect 8878 22848 8884 22900
rect 8936 22888 8942 22900
rect 9341 22891 9399 22897
rect 9341 22888 9353 22891
rect 8936 22860 9353 22888
rect 8936 22848 8942 22860
rect 9341 22857 9353 22860
rect 9387 22888 9399 22891
rect 9617 22891 9675 22897
rect 9617 22888 9629 22891
rect 9387 22860 9629 22888
rect 9387 22857 9399 22860
rect 9341 22851 9399 22857
rect 9617 22857 9629 22860
rect 9663 22857 9675 22891
rect 9617 22851 9675 22857
rect 10629 22891 10687 22897
rect 10629 22857 10641 22891
rect 10675 22888 10687 22891
rect 10905 22891 10963 22897
rect 10905 22888 10917 22891
rect 10675 22860 10917 22888
rect 10675 22857 10687 22860
rect 10629 22851 10687 22857
rect 10905 22857 10917 22860
rect 10951 22888 10963 22891
rect 10994 22888 11000 22900
rect 10951 22860 11000 22888
rect 10951 22857 10963 22860
rect 10905 22851 10963 22857
rect 10994 22848 11000 22860
rect 11052 22848 11058 22900
rect 11917 22891 11975 22897
rect 11917 22857 11929 22891
rect 11963 22888 11975 22891
rect 13110 22888 13116 22900
rect 11963 22860 13116 22888
rect 11963 22857 11975 22860
rect 11917 22851 11975 22857
rect 13110 22848 13116 22860
rect 13168 22848 13174 22900
rect 16422 22888 16428 22900
rect 16335 22860 16428 22888
rect 16422 22848 16428 22860
rect 16480 22888 16486 22900
rect 16517 22891 16575 22897
rect 16517 22888 16529 22891
rect 16480 22860 16529 22888
rect 16480 22848 16486 22860
rect 16517 22857 16529 22860
rect 16563 22857 16575 22891
rect 16517 22851 16575 22857
rect 18173 22891 18231 22897
rect 18173 22857 18185 22891
rect 18219 22888 18231 22891
rect 18648 22888 18676 22916
rect 19277 22891 19335 22897
rect 19277 22888 19289 22891
rect 18219 22860 19289 22888
rect 18219 22857 18231 22860
rect 18173 22851 18231 22857
rect 19277 22857 19289 22860
rect 19323 22888 19335 22891
rect 21666 22888 21672 22900
rect 19323 22860 21672 22888
rect 19323 22857 19335 22860
rect 19277 22851 19335 22857
rect 21666 22848 21672 22860
rect 21724 22848 21730 22900
rect 24061 22891 24119 22897
rect 24061 22857 24073 22891
rect 24107 22888 24119 22891
rect 24426 22888 24432 22900
rect 24107 22860 24432 22888
rect 24107 22857 24119 22860
rect 24061 22851 24119 22857
rect 24426 22848 24432 22860
rect 24484 22848 24490 22900
rect 24702 22848 24708 22900
rect 24760 22888 24766 22900
rect 24760 22860 24932 22888
rect 24760 22848 24766 22860
rect 1904 22820 1932 22848
rect 2165 22823 2223 22829
rect 2165 22820 2177 22823
rect 1904 22792 2177 22820
rect 2165 22789 2177 22792
rect 2211 22820 2223 22823
rect 2349 22823 2407 22829
rect 2349 22820 2361 22823
rect 2211 22792 2361 22820
rect 2211 22789 2223 22792
rect 2165 22783 2223 22789
rect 2349 22789 2361 22792
rect 2395 22789 2407 22823
rect 12006 22820 12012 22832
rect 11967 22792 12012 22820
rect 2349 22783 2407 22789
rect 12006 22780 12012 22792
rect 12064 22780 12070 22832
rect 12282 22820 12288 22832
rect 12243 22792 12288 22820
rect 12282 22780 12288 22792
rect 12340 22780 12346 22832
rect 15962 22820 15968 22832
rect 15923 22792 15968 22820
rect 15962 22780 15968 22792
rect 16020 22780 16026 22832
rect 20838 22820 20844 22832
rect 20799 22792 20844 22820
rect 20838 22780 20844 22792
rect 20896 22780 20902 22832
rect 23877 22823 23935 22829
rect 23877 22789 23889 22823
rect 23923 22820 23935 22823
rect 24720 22820 24748 22848
rect 23923 22792 24748 22820
rect 23923 22789 23935 22792
rect 23877 22783 23935 22789
rect 400 22730 27264 22752
rect 400 22678 18870 22730
rect 18922 22678 18934 22730
rect 18986 22678 18998 22730
rect 19050 22678 19062 22730
rect 19114 22678 19126 22730
rect 19178 22678 27264 22730
rect 400 22656 27264 22678
rect 1337 22619 1395 22625
rect 1337 22585 1349 22619
rect 1383 22616 1395 22619
rect 1794 22616 1800 22628
rect 1383 22588 1800 22616
rect 1383 22585 1395 22588
rect 1337 22579 1395 22585
rect 1794 22576 1800 22588
rect 1852 22576 1858 22628
rect 2162 22616 2168 22628
rect 1904 22588 2168 22616
rect 1904 22557 1932 22588
rect 2162 22576 2168 22588
rect 2220 22576 2226 22628
rect 18538 22616 18544 22628
rect 18499 22588 18544 22616
rect 18538 22576 18544 22588
rect 18596 22576 18602 22628
rect 24242 22616 24248 22628
rect 24203 22588 24248 22616
rect 24242 22576 24248 22588
rect 24300 22576 24306 22628
rect 1061 22551 1119 22557
rect 1061 22517 1073 22551
rect 1107 22548 1119 22551
rect 1889 22551 1947 22557
rect 1889 22548 1901 22551
rect 1107 22520 1901 22548
rect 1107 22517 1119 22520
rect 1061 22511 1119 22517
rect 1889 22517 1901 22520
rect 1935 22517 1947 22551
rect 5198 22548 5204 22560
rect 5159 22520 5204 22548
rect 1889 22511 1947 22517
rect 5198 22508 5204 22520
rect 5256 22508 5262 22560
rect 17710 22548 17716 22560
rect 16348 22520 17716 22548
rect 16348 22492 16376 22520
rect 17710 22508 17716 22520
rect 17768 22508 17774 22560
rect 24702 22548 24708 22560
rect 24663 22520 24708 22548
rect 24702 22508 24708 22520
rect 24760 22508 24766 22560
rect 4189 22483 4247 22489
rect 4189 22449 4201 22483
rect 4235 22480 4247 22483
rect 4278 22480 4284 22492
rect 4235 22452 4284 22480
rect 4235 22449 4247 22452
rect 4189 22443 4247 22449
rect 4278 22440 4284 22452
rect 4336 22440 4342 22492
rect 4373 22483 4431 22489
rect 4373 22449 4385 22483
rect 4419 22480 4431 22483
rect 4922 22480 4928 22492
rect 4419 22452 4928 22480
rect 4419 22449 4431 22452
rect 4373 22443 4431 22449
rect 4922 22440 4928 22452
rect 4980 22480 4986 22492
rect 5017 22483 5075 22489
rect 5017 22480 5029 22483
rect 4980 22452 5029 22480
rect 4980 22440 4986 22452
rect 5017 22449 5029 22452
rect 5063 22449 5075 22483
rect 10994 22480 11000 22492
rect 10955 22452 11000 22480
rect 5017 22443 5075 22449
rect 10994 22440 11000 22452
rect 11052 22440 11058 22492
rect 11362 22440 11368 22492
rect 11420 22480 11426 22492
rect 11825 22483 11883 22489
rect 11825 22480 11837 22483
rect 11420 22452 11837 22480
rect 11420 22440 11426 22452
rect 11825 22449 11837 22452
rect 11871 22480 11883 22483
rect 12006 22480 12012 22492
rect 11871 22452 12012 22480
rect 11871 22449 11883 22452
rect 11825 22443 11883 22449
rect 12006 22440 12012 22452
rect 12064 22440 12070 22492
rect 12742 22480 12748 22492
rect 12703 22452 12748 22480
rect 12742 22440 12748 22452
rect 12800 22440 12806 22492
rect 16330 22480 16336 22492
rect 16291 22452 16336 22480
rect 16330 22440 16336 22452
rect 16388 22440 16394 22492
rect 16882 22480 16888 22492
rect 16843 22452 16888 22480
rect 16882 22440 16888 22452
rect 16940 22440 16946 22492
rect 20194 22480 20200 22492
rect 20155 22452 20200 22480
rect 20194 22440 20200 22452
rect 20252 22440 20258 22492
rect 20838 22440 20844 22492
rect 20896 22480 20902 22492
rect 21761 22483 21819 22489
rect 21761 22480 21773 22483
rect 20896 22452 21773 22480
rect 20896 22440 20902 22452
rect 21761 22449 21773 22452
rect 21807 22480 21819 22483
rect 22770 22480 22776 22492
rect 21807 22452 22776 22480
rect 21807 22449 21819 22452
rect 21761 22443 21819 22449
rect 22770 22440 22776 22452
rect 22828 22440 22834 22492
rect 24426 22480 24432 22492
rect 24387 22452 24432 22480
rect 24426 22440 24432 22452
rect 24484 22440 24490 22492
rect 1242 22372 1248 22424
rect 1300 22412 1306 22424
rect 1429 22415 1487 22421
rect 1429 22412 1441 22415
rect 1300 22384 1441 22412
rect 1300 22372 1306 22384
rect 1429 22381 1441 22384
rect 1475 22381 1487 22415
rect 1978 22412 1984 22424
rect 1939 22384 1984 22412
rect 1429 22375 1487 22381
rect 1978 22372 1984 22384
rect 2036 22372 2042 22424
rect 13389 22415 13447 22421
rect 13389 22381 13401 22415
rect 13435 22412 13447 22415
rect 13478 22412 13484 22424
rect 13435 22384 13484 22412
rect 13435 22381 13447 22384
rect 13389 22375 13447 22381
rect 13478 22372 13484 22384
rect 13536 22372 13542 22424
rect 16422 22412 16428 22424
rect 16383 22384 16428 22412
rect 16422 22372 16428 22384
rect 16480 22372 16486 22424
rect 16698 22372 16704 22424
rect 16756 22412 16762 22424
rect 16793 22415 16851 22421
rect 16793 22412 16805 22415
rect 16756 22384 16805 22412
rect 16756 22372 16762 22384
rect 16793 22381 16805 22384
rect 16839 22381 16851 22415
rect 20470 22412 20476 22424
rect 20431 22384 20476 22412
rect 16793 22375 16851 22381
rect 20470 22372 20476 22384
rect 20528 22372 20534 22424
rect 22402 22372 22408 22424
rect 22460 22412 22466 22424
rect 22681 22415 22739 22421
rect 22681 22412 22693 22415
rect 22460 22384 22693 22412
rect 22460 22372 22466 22384
rect 22681 22381 22693 22384
rect 22727 22412 22739 22415
rect 24242 22412 24248 22424
rect 22727 22384 24248 22412
rect 22727 22381 22739 22384
rect 22681 22375 22739 22381
rect 16514 22344 16520 22356
rect 16475 22316 16520 22344
rect 16514 22304 16520 22316
rect 16572 22304 16578 22356
rect 23417 22347 23475 22353
rect 23417 22313 23429 22347
rect 23463 22344 23475 22347
rect 23874 22344 23880 22356
rect 23463 22316 23880 22344
rect 23463 22313 23475 22316
rect 23417 22307 23475 22313
rect 23874 22304 23880 22316
rect 23932 22304 23938 22356
rect 4002 22276 4008 22288
rect 3963 22248 4008 22276
rect 4002 22236 4008 22248
rect 4060 22236 4066 22288
rect 7774 22276 7780 22288
rect 7735 22248 7780 22276
rect 7774 22236 7780 22248
rect 7832 22236 7838 22288
rect 10810 22276 10816 22288
rect 10771 22248 10816 22276
rect 10810 22236 10816 22248
rect 10868 22236 10874 22288
rect 15410 22276 15416 22288
rect 15371 22248 15416 22276
rect 15410 22236 15416 22248
rect 15468 22236 15474 22288
rect 19090 22276 19096 22288
rect 19051 22248 19096 22276
rect 19090 22236 19096 22248
rect 19148 22236 19154 22288
rect 21758 22276 21764 22288
rect 21719 22248 21764 22276
rect 21758 22236 21764 22248
rect 21816 22236 21822 22288
rect 22586 22236 22592 22288
rect 22644 22276 22650 22288
rect 22957 22279 23015 22285
rect 22957 22276 22969 22279
rect 22644 22248 22969 22276
rect 22644 22236 22650 22248
rect 22957 22245 22969 22248
rect 23003 22245 23015 22279
rect 22957 22239 23015 22245
rect 23230 22236 23236 22288
rect 23288 22276 23294 22288
rect 23509 22279 23567 22285
rect 23509 22276 23521 22279
rect 23288 22248 23521 22276
rect 23288 22236 23294 22248
rect 23509 22245 23521 22248
rect 23555 22245 23567 22279
rect 23509 22239 23567 22245
rect 23785 22279 23843 22285
rect 23785 22245 23797 22279
rect 23831 22276 23843 22279
rect 23984 22276 24012 22384
rect 24242 22372 24248 22384
rect 24300 22372 24306 22424
rect 23831 22248 24012 22276
rect 23831 22245 23843 22248
rect 23785 22239 23843 22245
rect 400 22186 27264 22208
rect 400 22134 3510 22186
rect 3562 22134 3574 22186
rect 3626 22134 3638 22186
rect 3690 22134 3702 22186
rect 3754 22134 3766 22186
rect 3818 22134 27264 22186
rect 400 22112 27264 22134
rect 4002 22072 4008 22084
rect 3963 22044 4008 22072
rect 4002 22032 4008 22044
rect 4060 22032 4066 22084
rect 5198 22032 5204 22084
rect 5256 22072 5262 22084
rect 5477 22075 5535 22081
rect 5477 22072 5489 22075
rect 5256 22044 5489 22072
rect 5256 22032 5262 22044
rect 5477 22041 5489 22044
rect 5523 22041 5535 22075
rect 5477 22035 5535 22041
rect 6394 22032 6400 22084
rect 6452 22072 6458 22084
rect 7501 22075 7559 22081
rect 7501 22072 7513 22075
rect 6452 22044 7513 22072
rect 6452 22032 6458 22044
rect 7501 22041 7513 22044
rect 7547 22072 7559 22075
rect 8326 22072 8332 22084
rect 7547 22044 8332 22072
rect 7547 22041 7559 22044
rect 7501 22035 7559 22041
rect 8326 22032 8332 22044
rect 8384 22032 8390 22084
rect 11362 22072 11368 22084
rect 11323 22044 11368 22072
rect 11362 22032 11368 22044
rect 11420 22032 11426 22084
rect 13110 22032 13116 22084
rect 13168 22072 13174 22084
rect 13573 22075 13631 22081
rect 13573 22072 13585 22075
rect 13168 22044 13585 22072
rect 13168 22032 13174 22044
rect 13573 22041 13585 22044
rect 13619 22072 13631 22075
rect 13941 22075 13999 22081
rect 13941 22072 13953 22075
rect 13619 22044 13953 22072
rect 13619 22041 13631 22044
rect 13573 22035 13631 22041
rect 13941 22041 13953 22044
rect 13987 22041 13999 22075
rect 13941 22035 13999 22041
rect 15229 22075 15287 22081
rect 15229 22041 15241 22075
rect 15275 22072 15287 22075
rect 16330 22072 16336 22084
rect 15275 22044 16336 22072
rect 15275 22041 15287 22044
rect 15229 22035 15287 22041
rect 16330 22032 16336 22044
rect 16388 22032 16394 22084
rect 16514 22072 16520 22084
rect 16475 22044 16520 22072
rect 16514 22032 16520 22044
rect 16572 22032 16578 22084
rect 19090 22032 19096 22084
rect 19148 22072 19154 22084
rect 21577 22075 21635 22081
rect 19148 22044 21252 22072
rect 19148 22032 19154 22044
rect 2162 21964 2168 22016
rect 2220 22004 2226 22016
rect 2257 22007 2315 22013
rect 2257 22004 2269 22007
rect 2220 21976 2269 22004
rect 2220 21964 2226 21976
rect 2257 21973 2269 21976
rect 2303 21973 2315 22007
rect 2257 21967 2315 21973
rect 3821 22007 3879 22013
rect 3821 21973 3833 22007
rect 3867 22004 3879 22007
rect 4278 22004 4284 22016
rect 3867 21976 4284 22004
rect 3867 21973 3879 21976
rect 3821 21967 3879 21973
rect 4278 21964 4284 21976
rect 4336 22004 4342 22016
rect 7317 22007 7375 22013
rect 4336 21976 4554 22004
rect 4336 21964 4342 21976
rect 969 21871 1027 21877
rect 969 21837 981 21871
rect 1015 21837 1027 21871
rect 2070 21868 2076 21880
rect 2031 21840 2076 21868
rect 969 21831 1027 21837
rect 877 21735 935 21741
rect 877 21701 889 21735
rect 923 21732 935 21735
rect 984 21732 1012 21831
rect 2070 21828 2076 21840
rect 2128 21828 2134 21880
rect 4189 21871 4247 21877
rect 4189 21837 4201 21871
rect 4235 21868 4247 21871
rect 4281 21871 4339 21877
rect 4281 21868 4293 21871
rect 4235 21840 4293 21868
rect 4235 21837 4247 21840
rect 4189 21831 4247 21837
rect 4281 21837 4293 21840
rect 4327 21837 4339 21871
rect 4526 21868 4554 21976
rect 7317 21973 7329 22007
rect 7363 22004 7375 22007
rect 7363 21976 8740 22004
rect 7363 21973 7375 21976
rect 7317 21967 7375 21973
rect 8712 21948 8740 21976
rect 10994 21964 11000 22016
rect 11052 22004 11058 22016
rect 12742 22004 12748 22016
rect 11052 21976 12748 22004
rect 11052 21964 11058 21976
rect 7406 21896 7412 21948
rect 7464 21936 7470 21948
rect 7869 21939 7927 21945
rect 7869 21936 7881 21939
rect 7464 21908 7881 21936
rect 7464 21896 7470 21908
rect 7869 21905 7881 21908
rect 7915 21905 7927 21939
rect 8694 21936 8700 21948
rect 8655 21908 8700 21936
rect 7869 21899 7927 21905
rect 8694 21896 8700 21908
rect 8752 21896 8758 21948
rect 10169 21939 10227 21945
rect 10169 21905 10181 21939
rect 10215 21936 10227 21939
rect 10810 21936 10816 21948
rect 10215 21908 10816 21936
rect 10215 21905 10227 21908
rect 10169 21899 10227 21905
rect 10810 21896 10816 21908
rect 10868 21936 10874 21948
rect 11089 21939 11147 21945
rect 11089 21936 11101 21939
rect 10868 21908 11101 21936
rect 10868 21896 10874 21908
rect 11089 21905 11101 21908
rect 11135 21905 11147 21939
rect 11089 21899 11147 21905
rect 5201 21871 5259 21877
rect 5201 21868 5213 21871
rect 4526 21840 5213 21868
rect 4281 21831 4339 21837
rect 5201 21837 5213 21840
rect 5247 21837 5259 21871
rect 5201 21831 5259 21837
rect 1242 21732 1248 21744
rect 923 21704 1248 21732
rect 923 21701 935 21704
rect 877 21695 935 21701
rect 1242 21692 1248 21704
rect 1300 21692 1306 21744
rect 4296 21732 4324 21831
rect 5750 21828 5756 21880
rect 5808 21868 5814 21880
rect 6213 21871 6271 21877
rect 6213 21868 6225 21871
rect 5808 21840 6225 21868
rect 5808 21828 5814 21840
rect 6213 21837 6225 21840
rect 6259 21868 6271 21871
rect 6489 21871 6547 21877
rect 6489 21868 6501 21871
rect 6259 21840 6501 21868
rect 6259 21837 6271 21840
rect 6213 21831 6271 21837
rect 6489 21837 6501 21840
rect 6535 21837 6547 21871
rect 7774 21868 7780 21880
rect 7735 21840 7780 21868
rect 6489 21831 6547 21837
rect 7774 21828 7780 21840
rect 7832 21828 7838 21880
rect 8326 21828 8332 21880
rect 8384 21868 8390 21880
rect 8574 21871 8632 21877
rect 8574 21868 8586 21871
rect 8384 21840 8586 21868
rect 8384 21828 8390 21840
rect 8574 21837 8586 21840
rect 8620 21837 8632 21871
rect 8574 21831 8632 21837
rect 10261 21871 10319 21877
rect 10261 21837 10273 21871
rect 10307 21868 10319 21871
rect 10997 21871 11055 21877
rect 10997 21868 11009 21871
rect 10307 21840 11009 21868
rect 10307 21837 10319 21840
rect 10261 21831 10319 21837
rect 10997 21837 11009 21840
rect 11043 21868 11055 21871
rect 11549 21871 11607 21877
rect 11549 21868 11561 21871
rect 11043 21840 11561 21868
rect 11043 21837 11055 21840
rect 10997 21831 11055 21837
rect 11549 21837 11561 21840
rect 11595 21868 11607 21871
rect 11730 21868 11736 21880
rect 11595 21840 11736 21868
rect 11595 21837 11607 21840
rect 11549 21831 11607 21837
rect 11730 21828 11736 21840
rect 11788 21828 11794 21880
rect 12668 21877 12696 21976
rect 12742 21964 12748 21976
rect 12800 22004 12806 22016
rect 13205 22007 13263 22013
rect 13205 22004 13217 22007
rect 12800 21976 13217 22004
rect 12800 21964 12806 21976
rect 13205 21973 13217 21976
rect 13251 22004 13263 22007
rect 13297 22007 13355 22013
rect 13297 22004 13309 22007
rect 13251 21976 13309 22004
rect 13251 21973 13263 21976
rect 13205 21967 13263 21973
rect 13297 21973 13309 21976
rect 13343 21973 13355 22007
rect 15410 22004 15416 22016
rect 15371 21976 15416 22004
rect 13297 21967 13355 21973
rect 15410 21964 15416 21976
rect 15468 21964 15474 22016
rect 16422 21964 16428 22016
rect 16480 22004 16486 22016
rect 16701 22007 16759 22013
rect 16701 22004 16713 22007
rect 16480 21976 16713 22004
rect 16480 21964 16486 21976
rect 16701 21973 16713 21976
rect 16747 22004 16759 22007
rect 16747 21976 17388 22004
rect 16747 21973 16759 21976
rect 16701 21967 16759 21973
rect 13021 21939 13079 21945
rect 13021 21905 13033 21939
rect 13067 21936 13079 21939
rect 13478 21936 13484 21948
rect 13067 21908 13484 21936
rect 13067 21905 13079 21908
rect 13021 21899 13079 21905
rect 13478 21896 13484 21908
rect 13536 21896 13542 21948
rect 14861 21939 14919 21945
rect 14861 21905 14873 21939
rect 14907 21936 14919 21939
rect 15962 21936 15968 21948
rect 14907 21908 15968 21936
rect 14907 21905 14919 21908
rect 14861 21899 14919 21905
rect 15962 21896 15968 21908
rect 16020 21936 16026 21948
rect 17360 21945 17388 21976
rect 16149 21939 16207 21945
rect 16149 21936 16161 21939
rect 16020 21908 16161 21936
rect 16020 21896 16026 21908
rect 16149 21905 16161 21908
rect 16195 21905 16207 21939
rect 16149 21899 16207 21905
rect 17345 21939 17403 21945
rect 17345 21905 17357 21939
rect 17391 21936 17403 21939
rect 17989 21939 18047 21945
rect 17989 21936 18001 21939
rect 17391 21908 18001 21936
rect 17391 21905 17403 21908
rect 17345 21899 17403 21905
rect 17989 21905 18001 21908
rect 18035 21905 18047 21939
rect 17989 21899 18047 21905
rect 18817 21939 18875 21945
rect 18817 21905 18829 21939
rect 18863 21936 18875 21939
rect 21224 21936 21252 22044
rect 21577 22041 21589 22075
rect 21623 22072 21635 22075
rect 22770 22072 22776 22084
rect 21623 22044 22776 22072
rect 21623 22041 21635 22044
rect 21577 22035 21635 22041
rect 22770 22032 22776 22044
rect 22828 22032 22834 22084
rect 22402 22004 22408 22016
rect 22363 21976 22408 22004
rect 22402 21964 22408 21976
rect 22460 21964 22466 22016
rect 23230 21936 23236 21948
rect 18863 21908 20516 21936
rect 21224 21908 23236 21936
rect 18863 21905 18875 21908
rect 18817 21899 18875 21905
rect 20488 21880 20516 21908
rect 23230 21896 23236 21908
rect 23288 21896 23294 21948
rect 24242 21896 24248 21948
rect 24300 21936 24306 21948
rect 25257 21939 25315 21945
rect 25257 21936 25269 21939
rect 24300 21908 25269 21936
rect 24300 21896 24306 21908
rect 25257 21905 25269 21908
rect 25303 21905 25315 21939
rect 25257 21899 25315 21905
rect 12653 21871 12711 21877
rect 12653 21837 12665 21871
rect 12699 21837 12711 21871
rect 12653 21831 12711 21837
rect 15045 21871 15103 21877
rect 15045 21837 15057 21871
rect 15091 21868 15103 21871
rect 15321 21871 15379 21877
rect 15321 21868 15333 21871
rect 15091 21840 15333 21868
rect 15091 21837 15103 21840
rect 15045 21831 15103 21837
rect 15321 21837 15333 21840
rect 15367 21837 15379 21871
rect 15870 21868 15876 21880
rect 15831 21840 15876 21868
rect 15321 21831 15379 21837
rect 4922 21800 4928 21812
rect 4883 21772 4928 21800
rect 4922 21760 4928 21772
rect 4980 21800 4986 21812
rect 5293 21803 5351 21809
rect 5293 21800 5305 21803
rect 4980 21772 5305 21800
rect 4980 21760 4986 21772
rect 5293 21769 5305 21772
rect 5339 21769 5351 21803
rect 5293 21763 5351 21769
rect 9985 21803 10043 21809
rect 9985 21769 9997 21803
rect 10031 21800 10043 21803
rect 10721 21803 10779 21809
rect 10721 21800 10733 21803
rect 10031 21772 10733 21800
rect 10031 21769 10043 21772
rect 9985 21763 10043 21769
rect 10721 21769 10733 21772
rect 10767 21800 10779 21803
rect 12377 21803 12435 21809
rect 12377 21800 12389 21803
rect 10767 21772 12389 21800
rect 10767 21769 10779 21772
rect 10721 21763 10779 21769
rect 12377 21769 12389 21772
rect 12423 21769 12435 21803
rect 13481 21803 13539 21809
rect 13481 21800 13493 21803
rect 12377 21763 12435 21769
rect 12760 21772 13493 21800
rect 4554 21732 4560 21744
rect 4296 21704 4560 21732
rect 4554 21692 4560 21704
rect 4612 21692 4618 21744
rect 6026 21692 6032 21744
rect 6084 21732 6090 21744
rect 6305 21735 6363 21741
rect 6305 21732 6317 21735
rect 6084 21704 6317 21732
rect 6084 21692 6090 21704
rect 6305 21701 6317 21704
rect 6351 21732 6363 21735
rect 6673 21735 6731 21741
rect 6673 21732 6685 21735
rect 6351 21704 6685 21732
rect 6351 21701 6363 21704
rect 6305 21695 6363 21701
rect 6673 21701 6685 21704
rect 6719 21701 6731 21735
rect 12392 21732 12420 21763
rect 12760 21741 12788 21772
rect 13481 21769 13493 21772
rect 13527 21800 13539 21803
rect 13757 21803 13815 21809
rect 13757 21800 13769 21803
rect 13527 21772 13769 21800
rect 13527 21769 13539 21772
rect 13481 21763 13539 21769
rect 13757 21769 13769 21772
rect 13803 21769 13815 21803
rect 15336 21800 15364 21831
rect 15870 21828 15876 21840
rect 15928 21828 15934 21880
rect 16698 21828 16704 21880
rect 16756 21868 16762 21880
rect 17437 21871 17495 21877
rect 17437 21868 17449 21871
rect 16756 21840 17449 21868
rect 16756 21828 16762 21840
rect 17437 21837 17449 21840
rect 17483 21868 17495 21871
rect 18173 21871 18231 21877
rect 18173 21868 18185 21871
rect 17483 21840 18185 21868
rect 17483 21837 17495 21840
rect 17437 21831 17495 21837
rect 18173 21837 18185 21840
rect 18219 21837 18231 21871
rect 19090 21868 19096 21880
rect 18173 21831 18231 21837
rect 18924 21840 19096 21868
rect 17069 21803 17127 21809
rect 17069 21800 17081 21803
rect 15336 21772 17081 21800
rect 13757 21763 13815 21769
rect 17069 21769 17081 21772
rect 17115 21800 17127 21803
rect 17158 21800 17164 21812
rect 17115 21772 17164 21800
rect 17115 21769 17127 21772
rect 17069 21763 17127 21769
rect 17158 21760 17164 21772
rect 17216 21800 17222 21812
rect 17897 21803 17955 21809
rect 17897 21800 17909 21803
rect 17216 21772 17909 21800
rect 17216 21760 17222 21772
rect 17897 21769 17909 21772
rect 17943 21769 17955 21803
rect 17897 21763 17955 21769
rect 12745 21735 12803 21741
rect 12745 21732 12757 21735
rect 12392 21704 12757 21732
rect 6673 21695 6731 21701
rect 12745 21701 12757 21704
rect 12791 21701 12803 21735
rect 12745 21695 12803 21701
rect 15962 21692 15968 21744
rect 16020 21732 16026 21744
rect 17342 21732 17348 21744
rect 16020 21704 17348 21732
rect 16020 21692 16026 21704
rect 17342 21692 17348 21704
rect 17400 21732 17406 21744
rect 18924 21732 18952 21840
rect 19090 21828 19096 21840
rect 19148 21828 19154 21880
rect 20470 21828 20476 21880
rect 20528 21828 20534 21880
rect 19001 21803 19059 21809
rect 19001 21769 19013 21803
rect 19047 21800 19059 21803
rect 19366 21800 19372 21812
rect 19047 21772 19372 21800
rect 19047 21769 19059 21772
rect 19001 21763 19059 21769
rect 19366 21760 19372 21772
rect 19424 21760 19430 21812
rect 21117 21803 21175 21809
rect 21117 21769 21129 21803
rect 21163 21769 21175 21803
rect 23138 21800 23144 21812
rect 23051 21772 23144 21800
rect 21117 21763 21175 21769
rect 17400 21704 18952 21732
rect 17400 21692 17406 21704
rect 20102 21692 20108 21744
rect 20160 21732 20166 21744
rect 21132 21732 21160 21763
rect 23138 21760 23144 21772
rect 23196 21800 23202 21812
rect 23509 21803 23567 21809
rect 23509 21800 23521 21803
rect 23196 21772 23521 21800
rect 23196 21760 23202 21772
rect 23509 21769 23521 21772
rect 23555 21769 23567 21803
rect 23509 21763 23567 21769
rect 24518 21760 24524 21812
rect 24576 21760 24582 21812
rect 21758 21732 21764 21744
rect 20160 21704 21160 21732
rect 21719 21704 21764 21732
rect 20160 21692 20166 21704
rect 21758 21692 21764 21704
rect 21816 21692 21822 21744
rect 22586 21732 22592 21744
rect 22547 21704 22592 21732
rect 22586 21692 22592 21704
rect 22644 21692 22650 21744
rect 23874 21692 23880 21744
rect 23932 21732 23938 21744
rect 24536 21732 24564 21760
rect 23932 21704 24564 21732
rect 23932 21692 23938 21704
rect 400 21642 27264 21664
rect 400 21590 18870 21642
rect 18922 21590 18934 21642
rect 18986 21590 18998 21642
rect 19050 21590 19062 21642
rect 19114 21590 19126 21642
rect 19178 21590 27264 21642
rect 400 21568 27264 21590
rect 1705 21531 1763 21537
rect 1705 21497 1717 21531
rect 1751 21528 1763 21531
rect 1978 21528 1984 21540
rect 1751 21500 1984 21528
rect 1751 21497 1763 21500
rect 1705 21491 1763 21497
rect 1978 21488 1984 21500
rect 2036 21488 2042 21540
rect 4278 21528 4284 21540
rect 4239 21500 4284 21528
rect 4278 21488 4284 21500
rect 4336 21488 4342 21540
rect 7406 21488 7412 21540
rect 7464 21528 7470 21540
rect 7685 21531 7743 21537
rect 7685 21528 7697 21531
rect 7464 21500 7697 21528
rect 7464 21488 7470 21500
rect 7685 21497 7697 21500
rect 7731 21497 7743 21531
rect 7685 21491 7743 21497
rect 10905 21531 10963 21537
rect 10905 21497 10917 21531
rect 10951 21528 10963 21531
rect 10994 21528 11000 21540
rect 10951 21500 11000 21528
rect 10951 21497 10963 21500
rect 10905 21491 10963 21497
rect 10994 21488 11000 21500
rect 11052 21488 11058 21540
rect 15413 21531 15471 21537
rect 15413 21497 15425 21531
rect 15459 21528 15471 21531
rect 15870 21528 15876 21540
rect 15459 21500 15876 21528
rect 15459 21497 15471 21500
rect 15413 21491 15471 21497
rect 15870 21488 15876 21500
rect 15928 21488 15934 21540
rect 16149 21531 16207 21537
rect 16149 21497 16161 21531
rect 16195 21528 16207 21531
rect 16882 21528 16888 21540
rect 16195 21500 16888 21528
rect 16195 21497 16207 21500
rect 16149 21491 16207 21497
rect 16882 21488 16888 21500
rect 16940 21488 16946 21540
rect 20470 21528 20476 21540
rect 20431 21500 20476 21528
rect 20470 21488 20476 21500
rect 20528 21488 20534 21540
rect 24337 21531 24395 21537
rect 24337 21528 24349 21531
rect 20948 21500 24349 21528
rect 1061 21463 1119 21469
rect 1061 21429 1073 21463
rect 1107 21460 1119 21463
rect 2070 21460 2076 21472
rect 1107 21432 2076 21460
rect 1107 21429 1119 21432
rect 1061 21423 1119 21429
rect 2070 21420 2076 21432
rect 2128 21420 2134 21472
rect 4922 21420 4928 21472
rect 4980 21460 4986 21472
rect 5017 21463 5075 21469
rect 5017 21460 5029 21463
rect 4980 21432 5029 21460
rect 4980 21420 4986 21432
rect 5017 21429 5029 21432
rect 5063 21429 5075 21463
rect 5017 21423 5075 21429
rect 11914 21420 11920 21472
rect 11972 21460 11978 21472
rect 12009 21463 12067 21469
rect 12009 21460 12021 21463
rect 11972 21432 12021 21460
rect 11972 21420 11978 21432
rect 12009 21429 12021 21432
rect 12055 21429 12067 21463
rect 12009 21423 12067 21429
rect 15965 21463 16023 21469
rect 15965 21429 15977 21463
rect 16011 21460 16023 21463
rect 16011 21432 16744 21460
rect 16011 21429 16023 21432
rect 15965 21423 16023 21429
rect 16716 21404 16744 21432
rect 20194 21420 20200 21472
rect 20252 21460 20258 21472
rect 20289 21463 20347 21469
rect 20289 21460 20301 21463
rect 20252 21432 20301 21460
rect 20252 21420 20258 21432
rect 20289 21429 20301 21432
rect 20335 21460 20347 21463
rect 20948 21460 20976 21500
rect 24337 21497 24349 21500
rect 24383 21528 24395 21531
rect 24426 21528 24432 21540
rect 24383 21500 24432 21528
rect 24383 21497 24395 21500
rect 24337 21491 24395 21497
rect 24426 21488 24432 21500
rect 24484 21488 24490 21540
rect 24702 21528 24708 21540
rect 24663 21500 24708 21528
rect 24702 21488 24708 21500
rect 24760 21488 24766 21540
rect 20335 21432 20976 21460
rect 22681 21463 22739 21469
rect 20335 21429 20347 21432
rect 20289 21423 20347 21429
rect 22681 21429 22693 21463
rect 22727 21460 22739 21463
rect 22770 21460 22776 21472
rect 22727 21432 22776 21460
rect 22727 21429 22739 21432
rect 22681 21423 22739 21429
rect 22770 21420 22776 21432
rect 22828 21460 22834 21472
rect 23138 21460 23144 21472
rect 22828 21432 23144 21460
rect 22828 21420 22834 21432
rect 23138 21420 23144 21432
rect 23196 21420 23202 21472
rect 1886 21392 1892 21404
rect 1847 21364 1892 21392
rect 1886 21352 1892 21364
rect 1944 21352 1950 21404
rect 4002 21352 4008 21404
rect 4060 21392 4066 21404
rect 4738 21392 4744 21404
rect 4060 21364 4744 21392
rect 4060 21352 4066 21364
rect 4738 21352 4744 21364
rect 4796 21392 4802 21404
rect 5109 21395 5167 21401
rect 5109 21392 5121 21395
rect 4796 21364 5121 21392
rect 4796 21352 4802 21364
rect 5109 21361 5121 21364
rect 5155 21361 5167 21395
rect 5109 21355 5167 21361
rect 7682 21352 7688 21404
rect 7740 21392 7746 21404
rect 9246 21392 9252 21404
rect 7740 21364 9252 21392
rect 7740 21352 7746 21364
rect 9246 21352 9252 21364
rect 9304 21352 9310 21404
rect 9430 21392 9436 21404
rect 9391 21364 9436 21392
rect 9430 21352 9436 21364
rect 9488 21352 9494 21404
rect 11822 21352 11828 21404
rect 11880 21392 11886 21404
rect 12745 21395 12803 21401
rect 12745 21392 12757 21395
rect 11880 21364 12757 21392
rect 11880 21352 11886 21364
rect 12745 21361 12757 21364
rect 12791 21392 12803 21395
rect 13294 21392 13300 21404
rect 12791 21364 13300 21392
rect 12791 21361 12803 21364
rect 12745 21355 12803 21361
rect 13294 21352 13300 21364
rect 13352 21352 13358 21404
rect 16422 21392 16428 21404
rect 16383 21364 16428 21392
rect 16422 21352 16428 21364
rect 16480 21352 16486 21404
rect 16698 21392 16704 21404
rect 16659 21364 16704 21392
rect 16698 21352 16704 21364
rect 16756 21352 16762 21404
rect 17158 21392 17164 21404
rect 17119 21364 17164 21392
rect 17158 21352 17164 21364
rect 17216 21352 17222 21404
rect 17253 21395 17311 21401
rect 17253 21361 17265 21395
rect 17299 21361 17311 21395
rect 21298 21392 21304 21404
rect 21259 21364 21304 21392
rect 17253 21355 17311 21361
rect 4554 21284 4560 21336
rect 4612 21324 4618 21336
rect 11912 21327 11970 21333
rect 11912 21324 11924 21327
rect 4612 21296 4657 21324
rect 9540 21296 11924 21324
rect 4612 21284 4618 21296
rect 9540 21200 9568 21296
rect 11912 21293 11924 21296
rect 11958 21293 11970 21327
rect 11912 21287 11970 21293
rect 11932 21256 11960 21287
rect 12098 21284 12104 21336
rect 12156 21324 12162 21336
rect 12837 21327 12895 21333
rect 12837 21324 12849 21327
rect 12156 21296 12849 21324
rect 12156 21284 12162 21296
rect 12837 21293 12849 21296
rect 12883 21324 12895 21327
rect 12883 21296 14214 21324
rect 12883 21293 12895 21296
rect 12837 21287 12895 21293
rect 12190 21256 12196 21268
rect 11932 21228 12196 21256
rect 12190 21216 12196 21228
rect 12248 21216 12254 21268
rect 1242 21148 1248 21200
rect 1300 21188 1306 21200
rect 1429 21191 1487 21197
rect 1429 21188 1441 21191
rect 1300 21160 1441 21188
rect 1300 21148 1306 21160
rect 1429 21157 1441 21160
rect 1475 21157 1487 21191
rect 9522 21188 9528 21200
rect 9483 21160 9528 21188
rect 1429 21151 1487 21157
rect 9522 21148 9528 21160
rect 9580 21148 9586 21200
rect 13570 21188 13576 21200
rect 13531 21160 13576 21188
rect 13570 21148 13576 21160
rect 13628 21148 13634 21200
rect 14186 21188 14214 21296
rect 16790 21284 16796 21336
rect 16848 21324 16854 21336
rect 17268 21324 17296 21355
rect 21298 21352 21304 21364
rect 21356 21352 21362 21404
rect 21666 21392 21672 21404
rect 21627 21364 21672 21392
rect 21666 21352 21672 21364
rect 21724 21352 21730 21404
rect 22586 21352 22592 21404
rect 22644 21392 22650 21404
rect 23325 21395 23383 21401
rect 23325 21392 23337 21395
rect 22644 21364 23337 21392
rect 22644 21352 22650 21364
rect 23325 21361 23337 21364
rect 23371 21392 23383 21395
rect 23506 21392 23512 21404
rect 23371 21364 23512 21392
rect 23371 21361 23383 21364
rect 23325 21355 23383 21361
rect 23506 21352 23512 21364
rect 23564 21352 23570 21404
rect 23690 21392 23696 21404
rect 23651 21364 23696 21392
rect 23690 21352 23696 21364
rect 23748 21352 23754 21404
rect 21206 21324 21212 21336
rect 16848 21296 17296 21324
rect 21167 21296 21212 21324
rect 16848 21284 16854 21296
rect 21206 21284 21212 21296
rect 21264 21284 21270 21336
rect 21758 21324 21764 21336
rect 21671 21296 21764 21324
rect 21758 21284 21764 21296
rect 21816 21284 21822 21336
rect 23138 21284 23144 21336
rect 23196 21324 23202 21336
rect 23233 21327 23291 21333
rect 23233 21324 23245 21327
rect 23196 21296 23245 21324
rect 23196 21284 23202 21296
rect 23233 21293 23245 21296
rect 23279 21324 23291 21327
rect 23414 21324 23420 21336
rect 23279 21296 23420 21324
rect 23279 21293 23291 21296
rect 23233 21287 23291 21293
rect 23414 21284 23420 21296
rect 23472 21284 23478 21336
rect 23785 21327 23843 21333
rect 23785 21293 23797 21327
rect 23831 21293 23843 21327
rect 23785 21287 23843 21293
rect 16885 21259 16943 21265
rect 16885 21225 16897 21259
rect 16931 21256 16943 21259
rect 16974 21256 16980 21268
rect 16931 21228 16980 21256
rect 16931 21225 16943 21228
rect 16885 21219 16943 21225
rect 16974 21216 16980 21228
rect 17032 21216 17038 21268
rect 21776 21256 21804 21284
rect 23322 21256 23328 21268
rect 21776 21228 23328 21256
rect 23322 21216 23328 21228
rect 23380 21256 23386 21268
rect 23800 21256 23828 21287
rect 23380 21228 23828 21256
rect 23380 21216 23386 21228
rect 18262 21188 18268 21200
rect 14186 21160 18268 21188
rect 18262 21148 18268 21160
rect 18320 21148 18326 21200
rect 19185 21191 19243 21197
rect 19185 21157 19197 21191
rect 19231 21188 19243 21191
rect 20102 21188 20108 21200
rect 19231 21160 20108 21188
rect 19231 21157 19243 21160
rect 19185 21151 19243 21157
rect 20102 21148 20108 21160
rect 20160 21148 20166 21200
rect 20746 21188 20752 21200
rect 20707 21160 20752 21188
rect 20746 21148 20752 21160
rect 20804 21148 20810 21200
rect 24337 21191 24395 21197
rect 24337 21157 24349 21191
rect 24383 21188 24395 21191
rect 24521 21191 24579 21197
rect 24521 21188 24533 21191
rect 24383 21160 24533 21188
rect 24383 21157 24395 21160
rect 24337 21151 24395 21157
rect 24521 21157 24533 21160
rect 24567 21188 24579 21191
rect 24610 21188 24616 21200
rect 24567 21160 24616 21188
rect 24567 21157 24579 21160
rect 24521 21151 24579 21157
rect 24610 21148 24616 21160
rect 24668 21148 24674 21200
rect 400 21098 27264 21120
rect 400 21046 3510 21098
rect 3562 21046 3574 21098
rect 3626 21046 3638 21098
rect 3690 21046 3702 21098
rect 3754 21046 3766 21098
rect 3818 21046 27264 21098
rect 400 21024 27264 21046
rect 1886 20984 1892 20996
rect 1847 20956 1892 20984
rect 1886 20944 1892 20956
rect 1944 20944 1950 20996
rect 1978 20944 1984 20996
rect 2036 20984 2042 20996
rect 2073 20987 2131 20993
rect 2073 20984 2085 20987
rect 2036 20956 2085 20984
rect 2036 20944 2042 20956
rect 2073 20953 2085 20956
rect 2119 20953 2131 20987
rect 4738 20984 4744 20996
rect 4699 20956 4744 20984
rect 2073 20947 2131 20953
rect 4738 20944 4744 20956
rect 4796 20944 4802 20996
rect 4922 20984 4928 20996
rect 4883 20956 4928 20984
rect 4922 20944 4928 20956
rect 4980 20944 4986 20996
rect 9246 20944 9252 20996
rect 9304 20984 9310 20996
rect 9433 20987 9491 20993
rect 9433 20984 9445 20987
rect 9304 20956 9445 20984
rect 9304 20944 9310 20956
rect 9433 20953 9445 20956
rect 9479 20953 9491 20987
rect 9433 20947 9491 20953
rect 9522 20944 9528 20996
rect 9580 20984 9586 20996
rect 9617 20987 9675 20993
rect 9617 20984 9629 20987
rect 9580 20956 9629 20984
rect 9580 20944 9586 20956
rect 9617 20953 9629 20956
rect 9663 20953 9675 20987
rect 12190 20984 12196 20996
rect 12151 20956 12196 20984
rect 9617 20947 9675 20953
rect 12190 20944 12196 20956
rect 12248 20944 12254 20996
rect 13294 20984 13300 20996
rect 13255 20956 13300 20984
rect 13294 20944 13300 20956
rect 13352 20944 13358 20996
rect 16333 20987 16391 20993
rect 16333 20953 16345 20987
rect 16379 20984 16391 20987
rect 16422 20984 16428 20996
rect 16379 20956 16428 20984
rect 16379 20953 16391 20956
rect 16333 20947 16391 20953
rect 16422 20944 16428 20956
rect 16480 20944 16486 20996
rect 16701 20987 16759 20993
rect 16701 20953 16713 20987
rect 16747 20984 16759 20987
rect 17158 20984 17164 20996
rect 16747 20956 17164 20984
rect 16747 20953 16759 20956
rect 16701 20947 16759 20953
rect 17158 20944 17164 20956
rect 17216 20944 17222 20996
rect 19366 20944 19372 20996
rect 19424 20984 19430 20996
rect 19921 20987 19979 20993
rect 19921 20984 19933 20987
rect 19424 20956 19933 20984
rect 19424 20944 19430 20956
rect 19921 20953 19933 20956
rect 19967 20984 19979 20987
rect 20289 20987 20347 20993
rect 20289 20984 20301 20987
rect 19967 20956 20301 20984
rect 19967 20953 19979 20956
rect 19921 20947 19979 20953
rect 20289 20953 20301 20956
rect 20335 20953 20347 20987
rect 20289 20947 20347 20953
rect 21117 20987 21175 20993
rect 21117 20953 21129 20987
rect 21163 20984 21175 20987
rect 21758 20984 21764 20996
rect 21163 20956 21764 20984
rect 21163 20953 21175 20956
rect 21117 20947 21175 20953
rect 21758 20944 21764 20956
rect 21816 20944 21822 20996
rect 22770 20984 22776 20996
rect 22731 20956 22776 20984
rect 22770 20944 22776 20956
rect 22828 20944 22834 20996
rect 23506 20984 23512 20996
rect 23467 20956 23512 20984
rect 23506 20944 23512 20956
rect 23564 20944 23570 20996
rect 12098 20916 12104 20928
rect 12059 20888 12104 20916
rect 12098 20876 12104 20888
rect 12156 20876 12162 20928
rect 16974 20916 16980 20928
rect 16935 20888 16980 20916
rect 16974 20876 16980 20888
rect 17032 20876 17038 20928
rect 4554 20808 4560 20860
rect 4612 20848 4618 20860
rect 4649 20851 4707 20857
rect 4649 20848 4661 20851
rect 4612 20820 4661 20848
rect 4612 20808 4618 20820
rect 4649 20817 4661 20820
rect 4695 20848 4707 20851
rect 10166 20848 10172 20860
rect 4695 20820 10172 20848
rect 4695 20817 4707 20820
rect 4649 20811 4707 20817
rect 10166 20808 10172 20820
rect 10224 20808 10230 20860
rect 13205 20851 13263 20857
rect 13205 20817 13217 20851
rect 13251 20848 13263 20851
rect 16517 20851 16575 20857
rect 13251 20820 14536 20848
rect 13251 20817 13263 20820
rect 13205 20811 13263 20817
rect 7593 20783 7651 20789
rect 7593 20749 7605 20783
rect 7639 20780 7651 20783
rect 13570 20780 13576 20792
rect 7639 20752 8372 20780
rect 13531 20752 13576 20780
rect 7639 20749 7651 20752
rect 7593 20743 7651 20749
rect 7038 20672 7044 20724
rect 7096 20712 7102 20724
rect 7409 20715 7467 20721
rect 7409 20712 7421 20715
rect 7096 20684 7421 20712
rect 7096 20672 7102 20684
rect 7409 20681 7421 20684
rect 7455 20712 7467 20715
rect 8237 20715 8295 20721
rect 8237 20712 8249 20715
rect 7455 20684 8249 20712
rect 7455 20681 7467 20684
rect 7409 20675 7467 20681
rect 8237 20681 8249 20684
rect 8283 20681 8295 20715
rect 8237 20675 8295 20681
rect 6210 20604 6216 20656
rect 6268 20644 6274 20656
rect 7317 20647 7375 20653
rect 7317 20644 7329 20647
rect 6268 20616 7329 20644
rect 6268 20604 6274 20616
rect 7317 20613 7329 20616
rect 7363 20644 7375 20647
rect 7685 20647 7743 20653
rect 7685 20644 7697 20647
rect 7363 20616 7697 20644
rect 7363 20613 7375 20616
rect 7317 20607 7375 20613
rect 7685 20613 7697 20616
rect 7731 20613 7743 20647
rect 7685 20607 7743 20613
rect 8145 20647 8203 20653
rect 8145 20613 8157 20647
rect 8191 20644 8203 20647
rect 8344 20644 8372 20752
rect 13570 20740 13576 20752
rect 13628 20740 13634 20792
rect 14508 20789 14536 20820
rect 16517 20817 16529 20851
rect 16563 20848 16575 20851
rect 16698 20848 16704 20860
rect 16563 20820 16704 20848
rect 16563 20817 16575 20820
rect 16517 20811 16575 20817
rect 16698 20808 16704 20820
rect 16756 20808 16762 20860
rect 24518 20808 24524 20860
rect 24576 20848 24582 20860
rect 24889 20851 24947 20857
rect 24889 20848 24901 20851
rect 24576 20820 24901 20848
rect 24576 20808 24582 20820
rect 24889 20817 24901 20820
rect 24935 20848 24947 20851
rect 25349 20851 25407 20857
rect 25349 20848 25361 20851
rect 24935 20820 25361 20848
rect 24935 20817 24947 20820
rect 24889 20811 24947 20817
rect 25349 20817 25361 20820
rect 25395 20817 25407 20851
rect 25349 20811 25407 20817
rect 14401 20783 14459 20789
rect 14401 20780 14413 20783
rect 14186 20752 14413 20780
rect 9341 20715 9399 20721
rect 9341 20681 9353 20715
rect 9387 20712 9399 20715
rect 9522 20712 9528 20724
rect 9387 20684 9528 20712
rect 9387 20681 9399 20684
rect 9341 20675 9399 20681
rect 9356 20644 9384 20675
rect 9522 20672 9528 20684
rect 9580 20672 9586 20724
rect 11914 20672 11920 20724
rect 11972 20712 11978 20724
rect 12377 20715 12435 20721
rect 12377 20712 12389 20715
rect 11972 20684 12389 20712
rect 11972 20672 11978 20684
rect 12377 20681 12389 20684
rect 12423 20681 12435 20715
rect 12377 20675 12435 20681
rect 13021 20715 13079 20721
rect 13021 20681 13033 20715
rect 13067 20712 13079 20715
rect 13665 20715 13723 20721
rect 13665 20712 13677 20715
rect 13067 20684 13677 20712
rect 13067 20681 13079 20684
rect 13021 20675 13079 20681
rect 13665 20681 13677 20684
rect 13711 20712 13723 20715
rect 13754 20712 13760 20724
rect 13711 20684 13760 20712
rect 13711 20681 13723 20684
rect 13665 20675 13723 20681
rect 13754 20672 13760 20684
rect 13812 20672 13818 20724
rect 11822 20644 11828 20656
rect 8191 20616 9384 20644
rect 11783 20616 11828 20644
rect 8191 20613 8203 20616
rect 8145 20607 8203 20613
rect 11822 20604 11828 20616
rect 11880 20604 11886 20656
rect 13294 20604 13300 20656
rect 13352 20644 13358 20656
rect 14186 20644 14214 20752
rect 14401 20749 14413 20752
rect 14447 20749 14459 20783
rect 14401 20743 14459 20749
rect 14493 20783 14551 20789
rect 14493 20749 14505 20783
rect 14539 20749 14551 20783
rect 14493 20743 14551 20749
rect 20105 20783 20163 20789
rect 20105 20749 20117 20783
rect 20151 20780 20163 20783
rect 20565 20783 20623 20789
rect 20565 20780 20577 20783
rect 20151 20752 20577 20780
rect 20151 20749 20163 20752
rect 20105 20743 20163 20749
rect 20565 20749 20577 20752
rect 20611 20780 20623 20783
rect 20746 20780 20752 20792
rect 20611 20752 20752 20780
rect 20611 20749 20623 20752
rect 20565 20743 20623 20749
rect 14508 20712 14536 20743
rect 20746 20740 20752 20752
rect 20804 20780 20810 20792
rect 21393 20783 21451 20789
rect 21393 20780 21405 20783
rect 20804 20752 21405 20780
rect 20804 20740 20810 20752
rect 21393 20749 21405 20752
rect 21439 20749 21451 20783
rect 24610 20780 24616 20792
rect 24523 20752 24616 20780
rect 21393 20743 21451 20749
rect 24610 20740 24616 20752
rect 24668 20780 24674 20792
rect 24668 20752 25208 20780
rect 24668 20740 24674 20752
rect 20286 20712 20292 20724
rect 14508 20684 20292 20712
rect 20286 20672 20292 20684
rect 20344 20672 20350 20724
rect 20933 20715 20991 20721
rect 20933 20681 20945 20715
rect 20979 20712 20991 20715
rect 21666 20712 21672 20724
rect 20979 20684 21672 20712
rect 20979 20681 20991 20684
rect 20933 20675 20991 20681
rect 21666 20672 21672 20684
rect 21724 20712 21730 20724
rect 22034 20712 22040 20724
rect 21724 20684 22040 20712
rect 21724 20672 21730 20684
rect 22034 20672 22040 20684
rect 22092 20672 22098 20724
rect 23049 20715 23107 20721
rect 23049 20681 23061 20715
rect 23095 20712 23107 20715
rect 23690 20712 23696 20724
rect 23095 20684 23696 20712
rect 23095 20681 23107 20684
rect 23049 20675 23107 20681
rect 23690 20672 23696 20684
rect 23748 20712 23754 20724
rect 24150 20712 24156 20724
rect 23748 20684 24156 20712
rect 23748 20672 23754 20684
rect 24150 20672 24156 20684
rect 24208 20672 24214 20724
rect 25180 20656 25208 20752
rect 16790 20644 16796 20656
rect 13352 20616 14214 20644
rect 16751 20616 16796 20644
rect 13352 20604 13358 20616
rect 16790 20604 16796 20616
rect 16848 20604 16854 20656
rect 18354 20604 18360 20656
rect 18412 20644 18418 20656
rect 20657 20647 20715 20653
rect 20657 20644 20669 20647
rect 18412 20616 20669 20644
rect 18412 20604 18418 20616
rect 20657 20613 20669 20616
rect 20703 20644 20715 20647
rect 21206 20644 21212 20656
rect 20703 20616 21212 20644
rect 20703 20613 20715 20616
rect 20657 20607 20715 20613
rect 21206 20604 21212 20616
rect 21264 20604 21270 20656
rect 21301 20647 21359 20653
rect 21301 20613 21313 20647
rect 21347 20644 21359 20647
rect 21390 20644 21396 20656
rect 21347 20616 21396 20644
rect 21347 20613 21359 20616
rect 21301 20607 21359 20613
rect 21390 20604 21396 20616
rect 21448 20604 21454 20656
rect 23138 20644 23144 20656
rect 23099 20616 23144 20644
rect 23138 20604 23144 20616
rect 23196 20604 23202 20656
rect 23322 20644 23328 20656
rect 23283 20616 23328 20644
rect 23322 20604 23328 20616
rect 23380 20604 23386 20656
rect 25162 20644 25168 20656
rect 25123 20616 25168 20644
rect 25162 20604 25168 20616
rect 25220 20604 25226 20656
rect 400 20554 27264 20576
rect 400 20502 18870 20554
rect 18922 20502 18934 20554
rect 18986 20502 18998 20554
rect 19050 20502 19062 20554
rect 19114 20502 19126 20554
rect 19178 20502 27264 20554
rect 400 20480 27264 20502
rect 6121 20443 6179 20449
rect 6121 20409 6133 20443
rect 6167 20440 6179 20443
rect 6394 20440 6400 20452
rect 6167 20412 6400 20440
rect 6167 20409 6179 20412
rect 6121 20403 6179 20409
rect 6394 20400 6400 20412
rect 6452 20440 6458 20452
rect 7774 20440 7780 20452
rect 6452 20412 7780 20440
rect 6452 20400 6458 20412
rect 7774 20400 7780 20412
rect 7832 20400 7838 20452
rect 8142 20440 8148 20452
rect 8055 20412 8148 20440
rect 8142 20400 8148 20412
rect 8200 20440 8206 20452
rect 11086 20440 11092 20452
rect 8200 20412 11092 20440
rect 8200 20400 8206 20412
rect 11086 20400 11092 20412
rect 11144 20400 11150 20452
rect 23230 20400 23236 20452
rect 23288 20440 23294 20452
rect 23785 20443 23843 20449
rect 23785 20440 23797 20443
rect 23288 20412 23797 20440
rect 23288 20400 23294 20412
rect 23785 20409 23797 20412
rect 23831 20409 23843 20443
rect 23785 20403 23843 20409
rect 9985 20375 10043 20381
rect 4526 20344 7452 20372
rect 4526 20316 4554 20344
rect 877 20307 935 20313
rect 877 20273 889 20307
rect 923 20304 935 20307
rect 1242 20304 1248 20316
rect 923 20276 1248 20304
rect 923 20273 935 20276
rect 877 20267 935 20273
rect 1242 20264 1248 20276
rect 1300 20264 1306 20316
rect 1518 20264 1524 20316
rect 1576 20304 1582 20316
rect 1613 20307 1671 20313
rect 1613 20304 1625 20307
rect 1576 20276 1625 20304
rect 1576 20264 1582 20276
rect 1613 20273 1625 20276
rect 1659 20273 1671 20307
rect 1613 20267 1671 20273
rect 4097 20307 4155 20313
rect 4097 20273 4109 20307
rect 4143 20304 4155 20307
rect 4281 20307 4339 20313
rect 4143 20276 4232 20304
rect 4143 20273 4155 20276
rect 4097 20267 4155 20273
rect 782 20236 788 20248
rect 743 20208 788 20236
rect 782 20196 788 20208
rect 840 20196 846 20248
rect 966 20196 972 20248
rect 1024 20236 1030 20248
rect 1705 20239 1763 20245
rect 1705 20236 1717 20239
rect 1024 20208 1717 20236
rect 1024 20196 1030 20208
rect 1705 20205 1717 20208
rect 1751 20205 1763 20239
rect 4204 20236 4232 20276
rect 4281 20273 4293 20307
rect 4327 20304 4339 20307
rect 4526 20304 4560 20316
rect 4327 20276 4560 20304
rect 4327 20273 4339 20276
rect 4281 20267 4339 20273
rect 4554 20264 4560 20276
rect 4612 20264 4618 20316
rect 5474 20304 5480 20316
rect 5435 20276 5480 20304
rect 5474 20264 5480 20276
rect 5532 20264 5538 20316
rect 7038 20304 7044 20316
rect 6999 20276 7044 20304
rect 7038 20264 7044 20276
rect 7096 20264 7102 20316
rect 5624 20239 5682 20245
rect 4204 20208 4554 20236
rect 1705 20199 1763 20205
rect 4370 20100 4376 20112
rect 4331 20072 4376 20100
rect 4370 20060 4376 20072
rect 4428 20060 4434 20112
rect 4526 20100 4554 20208
rect 5624 20205 5636 20239
rect 5670 20236 5682 20239
rect 5750 20236 5756 20248
rect 5670 20208 5756 20236
rect 5670 20205 5682 20208
rect 5624 20199 5682 20205
rect 5750 20196 5756 20208
rect 5808 20196 5814 20248
rect 5845 20239 5903 20245
rect 5845 20205 5857 20239
rect 5891 20236 5903 20239
rect 5934 20236 5940 20248
rect 5891 20208 5940 20236
rect 5891 20205 5903 20208
rect 5845 20199 5903 20205
rect 5934 20196 5940 20208
rect 5992 20196 5998 20248
rect 7424 20245 7452 20344
rect 9985 20341 9997 20375
rect 10031 20372 10043 20375
rect 10258 20372 10264 20384
rect 10031 20344 10264 20372
rect 10031 20341 10043 20344
rect 9985 20335 10043 20341
rect 10258 20332 10264 20344
rect 10316 20372 10322 20384
rect 13570 20372 13576 20384
rect 10316 20344 13576 20372
rect 10316 20332 10322 20344
rect 13570 20332 13576 20344
rect 13628 20332 13634 20384
rect 15410 20332 15416 20384
rect 15468 20372 15474 20384
rect 15468 20344 16100 20372
rect 15468 20332 15474 20344
rect 9430 20304 9436 20316
rect 9391 20276 9436 20304
rect 9430 20264 9436 20276
rect 9488 20264 9494 20316
rect 9617 20307 9675 20313
rect 9617 20273 9629 20307
rect 9663 20273 9675 20307
rect 13478 20304 13484 20316
rect 13439 20276 13484 20304
rect 9617 20267 9675 20273
rect 7409 20239 7467 20245
rect 7409 20205 7421 20239
rect 7455 20205 7467 20239
rect 7682 20236 7688 20248
rect 7643 20208 7688 20236
rect 7409 20199 7467 20205
rect 7682 20196 7688 20208
rect 7740 20196 7746 20248
rect 9338 20196 9344 20248
rect 9396 20236 9402 20248
rect 9632 20236 9660 20267
rect 13478 20264 13484 20276
rect 13536 20264 13542 20316
rect 16072 20313 16100 20344
rect 16422 20332 16428 20384
rect 16480 20332 16486 20384
rect 21758 20372 21764 20384
rect 21671 20344 21764 20372
rect 21758 20332 21764 20344
rect 21816 20372 21822 20384
rect 22402 20372 22408 20384
rect 21816 20344 22408 20372
rect 21816 20332 21822 20344
rect 22402 20332 22408 20344
rect 22460 20332 22466 20384
rect 16057 20307 16115 20313
rect 16057 20273 16069 20307
rect 16103 20273 16115 20307
rect 16790 20304 16796 20316
rect 16703 20276 16796 20304
rect 16057 20267 16115 20273
rect 16790 20264 16796 20276
rect 16848 20304 16854 20316
rect 17986 20304 17992 20316
rect 16848 20276 17992 20304
rect 16848 20264 16854 20276
rect 17986 20264 17992 20276
rect 18044 20264 18050 20316
rect 20102 20264 20108 20316
rect 20160 20304 20166 20316
rect 20197 20307 20255 20313
rect 20197 20304 20209 20307
rect 20160 20276 20209 20304
rect 20160 20264 20166 20276
rect 20197 20273 20209 20276
rect 20243 20304 20255 20307
rect 21853 20307 21911 20313
rect 21853 20304 21865 20307
rect 20243 20276 21865 20304
rect 20243 20273 20255 20276
rect 20197 20267 20255 20273
rect 21853 20273 21865 20276
rect 21899 20304 21911 20307
rect 22126 20304 22132 20316
rect 21899 20276 22132 20304
rect 21899 20273 21911 20276
rect 21853 20267 21911 20273
rect 22126 20264 22132 20276
rect 22184 20264 22190 20316
rect 9396 20208 9660 20236
rect 9396 20196 9402 20208
rect 7314 20168 7320 20180
rect 5584 20140 7320 20168
rect 5584 20112 5612 20140
rect 7314 20128 7320 20140
rect 7372 20128 7378 20180
rect 13662 20168 13668 20180
rect 13623 20140 13668 20168
rect 13662 20128 13668 20140
rect 13720 20128 13726 20180
rect 4646 20100 4652 20112
rect 4526 20072 4652 20100
rect 4646 20060 4652 20072
rect 4704 20100 4710 20112
rect 5566 20100 5572 20112
rect 4704 20072 5572 20100
rect 4704 20060 4710 20072
rect 5566 20060 5572 20072
rect 5624 20060 5630 20112
rect 5753 20103 5811 20109
rect 5753 20069 5765 20103
rect 5799 20100 5811 20103
rect 6210 20100 6216 20112
rect 5799 20072 6216 20100
rect 5799 20069 5811 20072
rect 5753 20063 5811 20069
rect 6210 20060 6216 20072
rect 6268 20060 6274 20112
rect 6854 20060 6860 20112
rect 6912 20100 6918 20112
rect 7179 20103 7237 20109
rect 7179 20100 7191 20103
rect 6912 20072 7191 20100
rect 6912 20060 6918 20072
rect 7179 20069 7191 20072
rect 7225 20069 7237 20103
rect 7866 20100 7872 20112
rect 7827 20072 7872 20100
rect 7179 20063 7237 20069
rect 7866 20060 7872 20072
rect 7924 20060 7930 20112
rect 20473 20103 20531 20109
rect 20473 20069 20485 20103
rect 20519 20100 20531 20103
rect 20930 20100 20936 20112
rect 20519 20072 20936 20100
rect 20519 20069 20531 20072
rect 20473 20063 20531 20069
rect 20930 20060 20936 20072
rect 20988 20060 20994 20112
rect 21577 20103 21635 20109
rect 21577 20069 21589 20103
rect 21623 20100 21635 20103
rect 21666 20100 21672 20112
rect 21623 20072 21672 20100
rect 21623 20069 21635 20072
rect 21577 20063 21635 20069
rect 21666 20060 21672 20072
rect 21724 20060 21730 20112
rect 22034 20100 22040 20112
rect 21995 20072 22040 20100
rect 22034 20060 22040 20072
rect 22092 20060 22098 20112
rect 400 20010 27264 20032
rect 400 19958 3510 20010
rect 3562 19958 3574 20010
rect 3626 19958 3638 20010
rect 3690 19958 3702 20010
rect 3754 19958 3766 20010
rect 3818 19958 27264 20010
rect 400 19936 27264 19958
rect 874 19896 880 19908
rect 835 19868 880 19896
rect 874 19856 880 19868
rect 932 19856 938 19908
rect 1242 19896 1248 19908
rect 1203 19868 1248 19896
rect 1242 19856 1248 19868
rect 1300 19856 1306 19908
rect 1705 19899 1763 19905
rect 1705 19865 1717 19899
rect 1751 19896 1763 19899
rect 2070 19896 2076 19908
rect 1751 19868 2076 19896
rect 1751 19865 1763 19868
rect 1705 19859 1763 19865
rect 2070 19856 2076 19868
rect 2128 19856 2134 19908
rect 5474 19896 5480 19908
rect 4526 19868 5480 19896
rect 782 19788 788 19840
rect 840 19828 846 19840
rect 1061 19831 1119 19837
rect 1061 19828 1073 19831
rect 840 19800 1073 19828
rect 840 19788 846 19800
rect 1061 19797 1073 19800
rect 1107 19797 1119 19831
rect 1061 19791 1119 19797
rect 4370 19720 4376 19772
rect 4428 19760 4434 19772
rect 4526 19760 4554 19868
rect 5474 19856 5480 19868
rect 5532 19856 5538 19908
rect 6210 19896 6216 19908
rect 6171 19868 6216 19896
rect 6210 19856 6216 19868
rect 6268 19856 6274 19908
rect 6394 19896 6400 19908
rect 6355 19868 6400 19896
rect 6394 19856 6400 19868
rect 6452 19856 6458 19908
rect 6765 19899 6823 19905
rect 6765 19865 6777 19899
rect 6811 19896 6823 19899
rect 7038 19896 7044 19908
rect 6811 19868 7044 19896
rect 6811 19865 6823 19868
rect 6765 19859 6823 19865
rect 7038 19856 7044 19868
rect 7096 19856 7102 19908
rect 7314 19896 7320 19908
rect 7275 19868 7320 19896
rect 7314 19856 7320 19868
rect 7372 19856 7378 19908
rect 7685 19899 7743 19905
rect 7685 19865 7697 19899
rect 7731 19896 7743 19899
rect 8513 19899 8571 19905
rect 8513 19896 8525 19899
rect 7731 19868 8525 19896
rect 7731 19865 7743 19868
rect 7685 19859 7743 19865
rect 8513 19865 8525 19868
rect 8559 19896 8571 19899
rect 8697 19899 8755 19905
rect 8697 19896 8709 19899
rect 8559 19868 8709 19896
rect 8559 19865 8571 19868
rect 8513 19859 8571 19865
rect 8697 19865 8709 19868
rect 8743 19896 8755 19899
rect 9249 19899 9307 19905
rect 9249 19896 9261 19899
rect 8743 19868 9261 19896
rect 8743 19865 8755 19868
rect 8697 19859 8755 19865
rect 9249 19865 9261 19868
rect 9295 19865 9307 19899
rect 9249 19859 9307 19865
rect 9430 19856 9436 19908
rect 9488 19896 9494 19908
rect 9985 19899 10043 19905
rect 9985 19896 9997 19899
rect 9488 19868 9997 19896
rect 9488 19856 9494 19868
rect 9985 19865 9997 19868
rect 10031 19865 10043 19899
rect 10258 19896 10264 19908
rect 10219 19868 10264 19896
rect 9985 19859 10043 19865
rect 10258 19856 10264 19868
rect 10316 19856 10322 19908
rect 13478 19896 13484 19908
rect 13439 19868 13484 19896
rect 13478 19856 13484 19868
rect 13536 19856 13542 19908
rect 15410 19856 15416 19908
rect 15468 19896 15474 19908
rect 15597 19899 15655 19905
rect 15597 19896 15609 19899
rect 15468 19868 15609 19896
rect 15468 19856 15474 19868
rect 15597 19865 15609 19868
rect 15643 19865 15655 19899
rect 15597 19859 15655 19865
rect 15873 19899 15931 19905
rect 15873 19865 15885 19899
rect 15919 19896 15931 19899
rect 16422 19896 16428 19908
rect 15919 19868 16428 19896
rect 15919 19865 15931 19868
rect 15873 19859 15931 19865
rect 16422 19856 16428 19868
rect 16480 19856 16486 19908
rect 19921 19899 19979 19905
rect 19921 19865 19933 19899
rect 19967 19896 19979 19899
rect 20473 19899 20531 19905
rect 20473 19896 20485 19899
rect 19967 19868 20485 19896
rect 19967 19865 19979 19868
rect 19921 19859 19979 19865
rect 20473 19865 20485 19868
rect 20519 19896 20531 19899
rect 20654 19896 20660 19908
rect 20519 19868 20660 19896
rect 20519 19865 20531 19868
rect 20473 19859 20531 19865
rect 20654 19856 20660 19868
rect 20712 19856 20718 19908
rect 20838 19856 20844 19908
rect 20896 19896 20902 19908
rect 21025 19899 21083 19905
rect 21025 19896 21037 19899
rect 20896 19868 21037 19896
rect 20896 19856 20902 19868
rect 21025 19865 21037 19868
rect 21071 19865 21083 19899
rect 21758 19896 21764 19908
rect 21719 19868 21764 19896
rect 21025 19859 21083 19865
rect 21758 19856 21764 19868
rect 21816 19856 21822 19908
rect 22126 19896 22132 19908
rect 22087 19868 22132 19896
rect 22126 19856 22132 19868
rect 22184 19856 22190 19908
rect 5014 19788 5020 19840
rect 5072 19828 5078 19840
rect 6489 19831 6547 19837
rect 6489 19828 6501 19831
rect 5072 19800 6501 19828
rect 5072 19788 5078 19800
rect 6489 19797 6501 19800
rect 6535 19828 6547 19831
rect 7547 19831 7605 19837
rect 7547 19828 7559 19831
rect 6535 19800 7559 19828
rect 6535 19797 6547 19800
rect 6489 19791 6547 19797
rect 7547 19797 7559 19800
rect 7593 19797 7605 19831
rect 7547 19791 7605 19797
rect 8329 19831 8387 19837
rect 8329 19797 8341 19831
rect 8375 19828 8387 19831
rect 9448 19828 9476 19856
rect 8375 19800 9476 19828
rect 15505 19831 15563 19837
rect 8375 19797 8387 19800
rect 8329 19791 8387 19797
rect 15505 19797 15517 19831
rect 15551 19828 15563 19831
rect 16790 19828 16796 19840
rect 15551 19800 16796 19828
rect 15551 19797 15563 19800
rect 15505 19791 15563 19797
rect 4428 19720 4554 19760
rect 5198 19720 5204 19772
rect 5256 19760 5262 19772
rect 7777 19763 7835 19769
rect 7777 19760 7789 19763
rect 5256 19732 7789 19760
rect 5256 19720 5262 19732
rect 7777 19729 7789 19732
rect 7823 19760 7835 19763
rect 7866 19760 7872 19772
rect 7823 19732 7872 19760
rect 7823 19729 7835 19732
rect 7777 19723 7835 19729
rect 7866 19720 7872 19732
rect 7924 19720 7930 19772
rect 8142 19760 8148 19772
rect 8103 19732 8148 19760
rect 8142 19720 8148 19732
rect 8200 19720 8206 19772
rect 4388 19706 4554 19720
rect 1613 19627 1671 19633
rect 1613 19593 1625 19627
rect 1659 19593 1671 19627
rect 1613 19587 1671 19593
rect 506 19516 512 19568
rect 564 19556 570 19568
rect 693 19559 751 19565
rect 693 19556 705 19559
rect 564 19528 705 19556
rect 564 19516 570 19528
rect 693 19525 705 19528
rect 739 19556 751 19559
rect 1518 19556 1524 19568
rect 739 19528 1524 19556
rect 739 19525 751 19528
rect 693 19519 751 19525
rect 1518 19516 1524 19528
rect 1576 19516 1582 19568
rect 1628 19556 1656 19587
rect 1702 19584 1708 19636
rect 1760 19624 1766 19636
rect 4388 19624 4416 19706
rect 5934 19652 5940 19704
rect 5992 19692 5998 19704
rect 6854 19692 6860 19704
rect 5992 19664 6860 19692
rect 5992 19652 5998 19664
rect 6854 19652 6860 19664
rect 6912 19652 6918 19704
rect 7409 19695 7467 19701
rect 7409 19661 7421 19695
rect 7455 19692 7467 19695
rect 8050 19692 8056 19704
rect 7455 19664 8056 19692
rect 7455 19661 7467 19664
rect 7409 19655 7467 19661
rect 8050 19652 8056 19664
rect 8108 19692 8114 19704
rect 8344 19692 8372 19791
rect 16790 19788 16796 19800
rect 16848 19788 16854 19840
rect 16974 19788 16980 19840
rect 17032 19828 17038 19840
rect 20013 19831 20071 19837
rect 20013 19828 20025 19831
rect 17032 19800 20025 19828
rect 17032 19788 17038 19800
rect 20013 19797 20025 19800
rect 20059 19797 20071 19831
rect 20013 19791 20071 19797
rect 18078 19720 18084 19772
rect 18136 19760 18142 19772
rect 18357 19763 18415 19769
rect 18357 19760 18369 19763
rect 18136 19732 18369 19760
rect 18136 19720 18142 19732
rect 18357 19729 18369 19732
rect 18403 19760 18415 19763
rect 18403 19732 19320 19760
rect 18403 19729 18415 19732
rect 18357 19723 18415 19729
rect 9157 19695 9215 19701
rect 9157 19692 9169 19695
rect 8108 19664 8372 19692
rect 8436 19664 9169 19692
rect 8108 19652 8114 19664
rect 4557 19627 4615 19633
rect 4557 19624 4569 19627
rect 1760 19596 4569 19624
rect 1760 19584 1766 19596
rect 4557 19593 4569 19596
rect 4603 19593 4615 19627
rect 5750 19624 5756 19636
rect 5663 19596 5756 19624
rect 4557 19587 4615 19593
rect 5750 19584 5756 19596
rect 5808 19624 5814 19636
rect 6578 19624 6584 19636
rect 5808 19596 6584 19624
rect 5808 19584 5814 19596
rect 6578 19584 6584 19596
rect 6636 19624 6642 19636
rect 8436 19624 8464 19664
rect 9157 19661 9169 19664
rect 9203 19692 9215 19695
rect 9617 19695 9675 19701
rect 9617 19692 9629 19695
rect 9203 19664 9629 19692
rect 9203 19661 9215 19664
rect 9157 19655 9215 19661
rect 9617 19661 9629 19664
rect 9663 19661 9675 19695
rect 9617 19655 9675 19661
rect 18449 19695 18507 19701
rect 18449 19661 18461 19695
rect 18495 19692 18507 19695
rect 18722 19692 18728 19704
rect 18495 19664 18728 19692
rect 18495 19661 18507 19664
rect 18449 19655 18507 19661
rect 18722 19652 18728 19664
rect 18780 19692 18786 19704
rect 19185 19695 19243 19701
rect 19185 19692 19197 19695
rect 18780 19664 19197 19692
rect 18780 19652 18786 19664
rect 19185 19661 19197 19664
rect 19231 19661 19243 19695
rect 19185 19655 19243 19661
rect 6636 19596 8464 19624
rect 8881 19627 8939 19633
rect 6636 19584 6642 19596
rect 8881 19593 8893 19627
rect 8927 19624 8939 19627
rect 8973 19627 9031 19633
rect 8973 19624 8985 19627
rect 8927 19596 8985 19624
rect 8927 19593 8939 19596
rect 8881 19587 8939 19593
rect 8973 19593 8985 19596
rect 9019 19624 9031 19627
rect 9338 19624 9344 19636
rect 9019 19596 9344 19624
rect 9019 19593 9031 19596
rect 8973 19587 9031 19593
rect 9338 19584 9344 19596
rect 9396 19624 9402 19636
rect 9801 19627 9859 19633
rect 9801 19624 9813 19627
rect 9396 19596 9813 19624
rect 9396 19584 9402 19596
rect 9801 19593 9813 19596
rect 9847 19593 9859 19627
rect 18909 19627 18967 19633
rect 18909 19624 18921 19627
rect 9801 19587 9859 19593
rect 18188 19596 18921 19624
rect 18188 19568 18216 19596
rect 18909 19593 18921 19596
rect 18955 19593 18967 19627
rect 18909 19587 18967 19593
rect 19093 19627 19151 19633
rect 19093 19593 19105 19627
rect 19139 19624 19151 19627
rect 19292 19624 19320 19732
rect 20028 19692 20056 19791
rect 20197 19763 20255 19769
rect 20197 19729 20209 19763
rect 20243 19760 20255 19763
rect 20470 19760 20476 19772
rect 20243 19732 20476 19760
rect 20243 19729 20255 19732
rect 20197 19723 20255 19729
rect 20470 19720 20476 19732
rect 20528 19760 20534 19772
rect 20856 19760 20884 19856
rect 21669 19831 21727 19837
rect 21669 19797 21681 19831
rect 21715 19828 21727 19831
rect 22034 19828 22040 19840
rect 21715 19800 22040 19828
rect 21715 19797 21727 19800
rect 21669 19791 21727 19797
rect 22034 19788 22040 19800
rect 22092 19788 22098 19840
rect 20528 19732 20884 19760
rect 20528 19720 20534 19732
rect 23230 19720 23236 19772
rect 23288 19760 23294 19772
rect 23785 19763 23843 19769
rect 23785 19760 23797 19763
rect 23288 19732 23797 19760
rect 23288 19720 23294 19732
rect 23785 19729 23797 19732
rect 23831 19729 23843 19763
rect 23785 19723 23843 19729
rect 20286 19692 20292 19704
rect 20028 19664 20292 19692
rect 20286 19652 20292 19664
rect 20344 19652 20350 19704
rect 20930 19692 20936 19704
rect 20843 19664 20936 19692
rect 20930 19652 20936 19664
rect 20988 19692 20994 19704
rect 21850 19692 21856 19704
rect 20988 19664 21856 19692
rect 20988 19652 20994 19664
rect 21850 19652 21856 19664
rect 21908 19652 21914 19704
rect 19366 19624 19372 19636
rect 19139 19596 19372 19624
rect 19139 19593 19151 19596
rect 19093 19587 19151 19593
rect 19366 19584 19372 19596
rect 19424 19624 19430 19636
rect 20948 19624 20976 19652
rect 19424 19596 20976 19624
rect 19424 19584 19430 19596
rect 21666 19584 21672 19636
rect 21724 19624 21730 19636
rect 22037 19627 22095 19633
rect 22037 19624 22049 19627
rect 21724 19596 22049 19624
rect 21724 19584 21730 19596
rect 22037 19593 22049 19596
rect 22083 19624 22095 19627
rect 23509 19627 23567 19633
rect 22083 19596 23276 19624
rect 22083 19593 22095 19596
rect 22037 19587 22095 19593
rect 23248 19568 23276 19596
rect 23509 19593 23521 19627
rect 23555 19624 23567 19627
rect 23555 19596 23920 19624
rect 23555 19593 23567 19596
rect 23509 19587 23567 19593
rect 1981 19559 2039 19565
rect 1981 19556 1993 19559
rect 1628 19528 1993 19556
rect 1981 19525 1993 19528
rect 2027 19556 2039 19559
rect 2254 19556 2260 19568
rect 2027 19528 2260 19556
rect 2027 19525 2039 19528
rect 1981 19519 2039 19525
rect 2254 19516 2260 19528
rect 2312 19516 2318 19568
rect 4186 19556 4192 19568
rect 4147 19528 4192 19556
rect 4186 19516 4192 19528
rect 4244 19516 4250 19568
rect 4281 19559 4339 19565
rect 4281 19525 4293 19559
rect 4327 19556 4339 19559
rect 4462 19556 4468 19568
rect 4327 19528 4468 19556
rect 4327 19525 4339 19528
rect 4281 19519 4339 19525
rect 4462 19516 4468 19528
rect 4520 19556 4526 19568
rect 4646 19556 4652 19568
rect 4520 19528 4652 19556
rect 4520 19516 4526 19528
rect 4646 19516 4652 19528
rect 4704 19516 4710 19568
rect 5934 19556 5940 19568
rect 5895 19528 5940 19556
rect 5934 19516 5940 19528
rect 5992 19516 5998 19568
rect 7130 19556 7136 19568
rect 7091 19528 7136 19556
rect 7130 19516 7136 19528
rect 7188 19516 7194 19568
rect 13662 19556 13668 19568
rect 13575 19528 13668 19556
rect 13662 19516 13668 19528
rect 13720 19556 13726 19568
rect 14122 19556 14128 19568
rect 13720 19528 14128 19556
rect 13720 19516 13726 19528
rect 14122 19516 14128 19528
rect 14180 19516 14186 19568
rect 18170 19556 18176 19568
rect 18131 19528 18176 19556
rect 18170 19516 18176 19528
rect 18228 19516 18234 19568
rect 23230 19556 23236 19568
rect 23191 19528 23236 19556
rect 23230 19516 23236 19528
rect 23288 19516 23294 19568
rect 23693 19559 23751 19565
rect 23693 19525 23705 19559
rect 23739 19556 23751 19559
rect 23782 19556 23788 19568
rect 23739 19528 23788 19556
rect 23739 19525 23751 19528
rect 23693 19519 23751 19525
rect 23782 19516 23788 19528
rect 23840 19516 23846 19568
rect 23892 19556 23920 19596
rect 23966 19584 23972 19636
rect 24024 19624 24030 19636
rect 24061 19627 24119 19633
rect 24061 19624 24073 19627
rect 24024 19596 24073 19624
rect 24024 19584 24030 19596
rect 24061 19593 24073 19596
rect 24107 19593 24119 19627
rect 25806 19624 25812 19636
rect 24061 19587 24119 19593
rect 24536 19556 24564 19624
rect 25767 19596 25812 19624
rect 25806 19584 25812 19596
rect 25864 19584 25870 19636
rect 24978 19556 24984 19568
rect 23892 19528 24984 19556
rect 24978 19516 24984 19528
rect 25036 19516 25042 19568
rect 400 19466 27264 19488
rect 400 19414 18870 19466
rect 18922 19414 18934 19466
rect 18986 19414 18998 19466
rect 19050 19414 19062 19466
rect 19114 19414 19126 19466
rect 19178 19414 27264 19466
rect 400 19392 27264 19414
rect 1334 19352 1340 19364
rect 1247 19324 1340 19352
rect 1334 19312 1340 19324
rect 1392 19352 1398 19364
rect 1702 19352 1708 19364
rect 1392 19324 1708 19352
rect 1392 19312 1398 19324
rect 1702 19312 1708 19324
rect 1760 19312 1766 19364
rect 7133 19355 7191 19361
rect 7133 19321 7145 19355
rect 7179 19352 7191 19355
rect 7682 19352 7688 19364
rect 7179 19324 7688 19352
rect 7179 19321 7191 19324
rect 7133 19315 7191 19321
rect 7682 19312 7688 19324
rect 7740 19312 7746 19364
rect 19645 19355 19703 19361
rect 19645 19321 19657 19355
rect 19691 19352 19703 19355
rect 20102 19352 20108 19364
rect 19691 19324 20108 19352
rect 19691 19321 19703 19324
rect 19645 19315 19703 19321
rect 20102 19312 20108 19324
rect 20160 19352 20166 19364
rect 20197 19355 20255 19361
rect 20197 19352 20209 19355
rect 20160 19324 20209 19352
rect 20160 19312 20166 19324
rect 20197 19321 20209 19324
rect 20243 19321 20255 19355
rect 20197 19315 20255 19321
rect 23049 19355 23107 19361
rect 23049 19321 23061 19355
rect 23095 19352 23107 19355
rect 23138 19352 23144 19364
rect 23095 19324 23144 19352
rect 23095 19321 23107 19324
rect 23049 19315 23107 19321
rect 23138 19312 23144 19324
rect 23196 19352 23202 19364
rect 23506 19352 23512 19364
rect 23196 19324 23512 19352
rect 23196 19312 23202 19324
rect 23506 19312 23512 19324
rect 23564 19312 23570 19364
rect 4554 19244 4560 19296
rect 4612 19284 4618 19296
rect 4649 19287 4707 19293
rect 4649 19284 4661 19287
rect 4612 19256 4661 19284
rect 4612 19244 4618 19256
rect 4649 19253 4661 19256
rect 4695 19284 4707 19287
rect 6210 19284 6216 19296
rect 4695 19256 6216 19284
rect 4695 19253 4707 19256
rect 4649 19247 4707 19253
rect 6210 19244 6216 19256
rect 6268 19244 6274 19296
rect 7038 19244 7044 19296
rect 7096 19284 7102 19296
rect 8053 19287 8111 19293
rect 8053 19284 8065 19287
rect 7096 19256 8065 19284
rect 7096 19244 7102 19256
rect 8053 19253 8065 19256
rect 8099 19253 8111 19287
rect 8053 19247 8111 19253
rect 17437 19287 17495 19293
rect 17437 19253 17449 19287
rect 17483 19284 17495 19287
rect 17483 19256 18768 19284
rect 17483 19253 17495 19256
rect 17437 19247 17495 19253
rect 18740 19228 18768 19256
rect 22402 19244 22408 19296
rect 22460 19284 22466 19296
rect 23417 19287 23475 19293
rect 23417 19284 23429 19287
rect 22460 19256 23429 19284
rect 22460 19244 22466 19256
rect 23417 19253 23429 19256
rect 23463 19284 23475 19287
rect 24058 19284 24064 19296
rect 23463 19256 24064 19284
rect 23463 19253 23475 19256
rect 23417 19247 23475 19253
rect 24058 19244 24064 19256
rect 24116 19244 24122 19296
rect 26174 19284 26180 19296
rect 26100 19256 26180 19284
rect 4738 19176 4744 19228
rect 4796 19216 4802 19228
rect 4833 19219 4891 19225
rect 4833 19216 4845 19219
rect 4796 19188 4845 19216
rect 4796 19176 4802 19188
rect 4833 19185 4845 19188
rect 4879 19185 4891 19219
rect 7590 19216 7596 19228
rect 7551 19188 7596 19216
rect 4833 19179 4891 19185
rect 7590 19176 7596 19188
rect 7648 19176 7654 19228
rect 9982 19176 9988 19228
rect 10040 19216 10046 19228
rect 10445 19219 10503 19225
rect 10445 19216 10457 19219
rect 10040 19188 10457 19216
rect 10040 19176 10046 19188
rect 10445 19185 10457 19188
rect 10491 19185 10503 19219
rect 11086 19216 11092 19228
rect 11047 19188 11092 19216
rect 10445 19179 10503 19185
rect 11086 19176 11092 19188
rect 11144 19216 11150 19228
rect 11822 19216 11828 19228
rect 11144 19188 11828 19216
rect 11144 19176 11150 19188
rect 11822 19176 11828 19188
rect 11880 19176 11886 19228
rect 12653 19219 12711 19225
rect 12653 19185 12665 19219
rect 12699 19216 12711 19219
rect 12926 19216 12932 19228
rect 12699 19188 12932 19216
rect 12699 19185 12711 19188
rect 12653 19179 12711 19185
rect 12926 19176 12932 19188
rect 12984 19176 12990 19228
rect 13478 19216 13484 19228
rect 13439 19188 13484 19216
rect 13478 19176 13484 19188
rect 13536 19176 13542 19228
rect 18357 19219 18415 19225
rect 18357 19185 18369 19219
rect 18403 19216 18415 19219
rect 18538 19216 18544 19228
rect 18403 19188 18544 19216
rect 18403 19185 18415 19188
rect 18357 19179 18415 19185
rect 18538 19176 18544 19188
rect 18596 19176 18602 19228
rect 18722 19216 18728 19228
rect 18683 19188 18728 19216
rect 18722 19176 18728 19188
rect 18780 19176 18786 19228
rect 18909 19219 18967 19225
rect 18909 19185 18921 19219
rect 18955 19216 18967 19219
rect 19366 19216 19372 19228
rect 18955 19188 19372 19216
rect 18955 19185 18967 19188
rect 18909 19179 18967 19185
rect 19366 19176 19372 19188
rect 19424 19176 19430 19228
rect 22218 19216 22224 19228
rect 22179 19188 22224 19216
rect 22218 19176 22224 19188
rect 22276 19176 22282 19228
rect 23322 19176 23328 19228
rect 23380 19216 23386 19228
rect 26100 19225 26128 19256
rect 26174 19244 26180 19256
rect 26232 19244 26238 19296
rect 23509 19219 23567 19225
rect 23509 19216 23521 19219
rect 23380 19188 23521 19216
rect 23380 19176 23386 19188
rect 23509 19185 23521 19188
rect 23555 19185 23567 19219
rect 23509 19179 23567 19185
rect 26085 19219 26143 19225
rect 26085 19185 26097 19219
rect 26131 19185 26143 19219
rect 26085 19179 26143 19185
rect 7498 19148 7504 19160
rect 7411 19120 7504 19148
rect 7498 19108 7504 19120
rect 7556 19148 7562 19160
rect 8970 19148 8976 19160
rect 7556 19120 8976 19148
rect 7556 19108 7562 19120
rect 8970 19108 8976 19120
rect 9028 19148 9034 19160
rect 10721 19151 10779 19157
rect 9028 19120 10580 19148
rect 9028 19108 9034 19120
rect 10166 19040 10172 19092
rect 10224 19080 10230 19092
rect 10445 19083 10503 19089
rect 10445 19080 10457 19083
rect 10224 19052 10457 19080
rect 10224 19040 10230 19052
rect 10445 19049 10457 19052
rect 10491 19049 10503 19083
rect 10552 19080 10580 19120
rect 10721 19117 10733 19151
rect 10767 19148 10779 19151
rect 10810 19148 10816 19160
rect 10767 19120 10816 19148
rect 10767 19117 10779 19120
rect 10721 19111 10779 19117
rect 10810 19108 10816 19120
rect 10868 19108 10874 19160
rect 10994 19148 11000 19160
rect 10955 19120 11000 19148
rect 10994 19108 11000 19120
rect 11052 19108 11058 19160
rect 12742 19108 12748 19160
rect 12800 19148 12806 19160
rect 13570 19148 13576 19160
rect 12800 19120 12845 19148
rect 13531 19120 13576 19148
rect 12800 19108 12806 19120
rect 13570 19108 13576 19120
rect 13628 19108 13634 19160
rect 18170 19148 18176 19160
rect 18131 19120 18176 19148
rect 18170 19108 18176 19120
rect 18228 19108 18234 19160
rect 21390 19148 21396 19160
rect 21351 19120 21396 19148
rect 21390 19108 21396 19120
rect 21448 19108 21454 19160
rect 21850 19108 21856 19160
rect 21908 19148 21914 19160
rect 21945 19151 22003 19157
rect 21945 19148 21957 19151
rect 21908 19120 21957 19148
rect 21908 19108 21914 19120
rect 21945 19117 21957 19120
rect 21991 19117 22003 19151
rect 22402 19148 22408 19160
rect 22363 19120 22408 19148
rect 21945 19111 22003 19117
rect 22402 19108 22408 19120
rect 22460 19108 22466 19160
rect 11012 19080 11040 19108
rect 10552 19052 11040 19080
rect 10445 19043 10503 19049
rect 16330 19040 16336 19092
rect 16388 19080 16394 19092
rect 17621 19083 17679 19089
rect 17621 19080 17633 19083
rect 16388 19052 17633 19080
rect 16388 19040 16394 19052
rect 17621 19049 17633 19052
rect 17667 19080 17679 19083
rect 17894 19080 17900 19092
rect 17667 19052 17900 19080
rect 17667 19049 17679 19052
rect 17621 19043 17679 19049
rect 17894 19040 17900 19052
rect 17952 19040 17958 19092
rect 19274 19040 19280 19092
rect 19332 19080 19338 19092
rect 19918 19080 19924 19092
rect 19332 19052 19924 19080
rect 19332 19040 19338 19052
rect 19918 19040 19924 19052
rect 19976 19040 19982 19092
rect 4925 19015 4983 19021
rect 4925 18981 4937 19015
rect 4971 19012 4983 19015
rect 5014 19012 5020 19024
rect 4971 18984 5020 19012
rect 4971 18981 4983 18984
rect 4925 18975 4983 18981
rect 5014 18972 5020 18984
rect 5072 18972 5078 19024
rect 13846 19012 13852 19024
rect 13807 18984 13852 19012
rect 13846 18972 13852 18984
rect 13904 18972 13910 19024
rect 17986 19012 17992 19024
rect 17947 18984 17992 19012
rect 17986 18972 17992 18984
rect 18044 18972 18050 19024
rect 23230 19012 23236 19024
rect 23191 18984 23236 19012
rect 23230 18972 23236 18984
rect 23288 18972 23294 19024
rect 23598 18972 23604 19024
rect 23656 19012 23662 19024
rect 23693 19015 23751 19021
rect 23693 19012 23705 19015
rect 23656 18984 23705 19012
rect 23656 18972 23662 18984
rect 23693 18981 23705 18984
rect 23739 18981 23751 19015
rect 26082 19012 26088 19024
rect 26043 18984 26088 19012
rect 23693 18975 23751 18981
rect 26082 18972 26088 18984
rect 26140 18972 26146 19024
rect 400 18922 27264 18944
rect 400 18870 3510 18922
rect 3562 18870 3574 18922
rect 3626 18870 3638 18922
rect 3690 18870 3702 18922
rect 3754 18870 3766 18922
rect 3818 18870 27264 18922
rect 400 18848 27264 18870
rect 782 18768 788 18820
rect 840 18808 846 18820
rect 1702 18808 1708 18820
rect 840 18780 1708 18808
rect 840 18768 846 18780
rect 1702 18768 1708 18780
rect 1760 18808 1766 18820
rect 2993 18811 3051 18817
rect 2993 18808 3005 18811
rect 1760 18780 3005 18808
rect 1760 18768 1766 18780
rect 2993 18777 3005 18780
rect 3039 18808 3051 18811
rect 3453 18811 3511 18817
rect 3453 18808 3465 18811
rect 3039 18780 3465 18808
rect 3039 18777 3051 18780
rect 2993 18771 3051 18777
rect 3453 18777 3465 18780
rect 3499 18777 3511 18811
rect 3453 18771 3511 18777
rect 4373 18811 4431 18817
rect 4373 18777 4385 18811
rect 4419 18808 4431 18811
rect 4554 18808 4560 18820
rect 4419 18780 4560 18808
rect 4419 18777 4431 18780
rect 4373 18771 4431 18777
rect 4554 18768 4560 18780
rect 4612 18808 4618 18820
rect 6949 18811 7007 18817
rect 4612 18780 4657 18808
rect 4612 18768 4618 18780
rect 6949 18777 6961 18811
rect 6995 18808 7007 18811
rect 7038 18808 7044 18820
rect 6995 18780 7044 18808
rect 6995 18777 7007 18780
rect 6949 18771 7007 18777
rect 7038 18768 7044 18780
rect 7096 18768 7102 18820
rect 7133 18811 7191 18817
rect 7133 18777 7145 18811
rect 7179 18808 7191 18811
rect 7685 18811 7743 18817
rect 7685 18808 7697 18811
rect 7179 18780 7697 18808
rect 7179 18777 7191 18780
rect 7133 18771 7191 18777
rect 7685 18777 7697 18780
rect 7731 18808 7743 18811
rect 8789 18811 8847 18817
rect 8789 18808 8801 18811
rect 7731 18780 8801 18808
rect 7731 18777 7743 18780
rect 7685 18771 7743 18777
rect 8789 18777 8801 18780
rect 8835 18808 8847 18811
rect 8835 18780 9016 18808
rect 8835 18777 8847 18780
rect 8789 18771 8847 18777
rect 874 18632 880 18684
rect 932 18672 938 18684
rect 2257 18675 2315 18681
rect 2257 18672 2269 18675
rect 932 18644 2269 18672
rect 932 18632 938 18644
rect 2257 18641 2269 18644
rect 2303 18641 2315 18675
rect 4572 18672 4600 18768
rect 4738 18700 4744 18752
rect 4796 18740 4802 18752
rect 5477 18743 5535 18749
rect 5477 18740 5489 18743
rect 4796 18712 5489 18740
rect 4796 18700 4802 18712
rect 5477 18709 5489 18712
rect 5523 18709 5535 18743
rect 5477 18703 5535 18709
rect 7317 18743 7375 18749
rect 7317 18709 7329 18743
rect 7363 18740 7375 18743
rect 7498 18740 7504 18752
rect 7363 18712 7504 18740
rect 7363 18709 7375 18712
rect 7317 18703 7375 18709
rect 7498 18700 7504 18712
rect 7556 18700 7562 18752
rect 8050 18740 8056 18752
rect 8011 18712 8056 18740
rect 8050 18700 8056 18712
rect 8108 18700 8114 18752
rect 8326 18740 8332 18752
rect 8287 18712 8332 18740
rect 8326 18700 8332 18712
rect 8384 18700 8390 18752
rect 4572 18644 4692 18672
rect 2257 18635 2315 18641
rect 1334 18604 1340 18616
rect 1295 18576 1340 18604
rect 1334 18564 1340 18576
rect 1392 18564 1398 18616
rect 2165 18607 2223 18613
rect 2165 18604 2177 18607
rect 2075 18576 2177 18604
rect 2165 18573 2177 18576
rect 2211 18573 2223 18607
rect 3358 18604 3364 18616
rect 3319 18576 3364 18604
rect 2165 18567 2223 18573
rect 506 18496 512 18548
rect 564 18536 570 18548
rect 1061 18539 1119 18545
rect 1061 18536 1073 18539
rect 564 18508 1073 18536
rect 564 18496 570 18508
rect 1061 18505 1073 18508
rect 1107 18505 1119 18539
rect 1061 18499 1119 18505
rect 874 18468 880 18480
rect 835 18440 880 18468
rect 874 18428 880 18440
rect 932 18428 938 18480
rect 1076 18468 1104 18499
rect 1242 18496 1248 18548
rect 1300 18536 1306 18548
rect 1429 18539 1487 18545
rect 1429 18536 1441 18539
rect 1300 18508 1441 18536
rect 1300 18496 1306 18508
rect 1429 18505 1441 18508
rect 1475 18505 1487 18539
rect 1429 18499 1487 18505
rect 2180 18468 2208 18567
rect 3358 18564 3364 18576
rect 3416 18604 3422 18616
rect 4664 18613 4692 18644
rect 4756 18644 5520 18672
rect 3821 18607 3879 18613
rect 3821 18604 3833 18607
rect 3416 18576 3833 18604
rect 3416 18564 3422 18576
rect 3821 18573 3833 18576
rect 3867 18604 3879 18607
rect 4649 18607 4707 18613
rect 3867 18576 4554 18604
rect 3867 18573 3879 18576
rect 3821 18567 3879 18573
rect 3177 18539 3235 18545
rect 3177 18505 3189 18539
rect 3223 18536 3235 18539
rect 4526 18536 4554 18576
rect 4649 18573 4661 18607
rect 4695 18573 4707 18607
rect 4649 18567 4707 18573
rect 4756 18536 4784 18644
rect 4833 18607 4891 18613
rect 4833 18573 4845 18607
rect 4879 18604 4891 18607
rect 5492 18604 5520 18644
rect 6302 18632 6308 18684
rect 6360 18672 6366 18684
rect 7038 18672 7044 18684
rect 6360 18644 7044 18672
rect 6360 18632 6366 18644
rect 7038 18632 7044 18644
rect 7096 18632 7102 18684
rect 7777 18675 7835 18681
rect 7777 18641 7789 18675
rect 7823 18672 7835 18675
rect 8344 18672 8372 18700
rect 7823 18644 8372 18672
rect 7823 18641 7835 18644
rect 7777 18635 7835 18641
rect 7498 18604 7504 18616
rect 4879 18576 5428 18604
rect 5492 18576 7504 18604
rect 4879 18573 4891 18576
rect 4833 18567 4891 18573
rect 3223 18508 4140 18536
rect 4526 18508 4784 18536
rect 3223 18505 3235 18508
rect 3177 18499 3235 18505
rect 4112 18477 4140 18508
rect 1076 18440 2208 18468
rect 4097 18471 4155 18477
rect 4097 18437 4109 18471
rect 4143 18468 4155 18471
rect 4462 18468 4468 18480
rect 4143 18440 4468 18468
rect 4143 18437 4155 18440
rect 4097 18431 4155 18437
rect 4462 18428 4468 18440
rect 4520 18428 4526 18480
rect 4922 18468 4928 18480
rect 4883 18440 4928 18468
rect 4922 18428 4928 18440
rect 4980 18428 4986 18480
rect 5400 18477 5428 18576
rect 7498 18564 7504 18576
rect 7556 18613 7562 18616
rect 7556 18607 7614 18613
rect 7556 18573 7568 18607
rect 7602 18573 7614 18607
rect 7556 18567 7614 18573
rect 7556 18564 7562 18567
rect 5566 18496 5572 18548
rect 5624 18536 5630 18548
rect 6765 18539 6823 18545
rect 6765 18536 6777 18539
rect 5624 18508 6777 18536
rect 5624 18496 5630 18508
rect 6765 18505 6777 18508
rect 6811 18536 6823 18539
rect 7409 18539 7467 18545
rect 7409 18536 7421 18539
rect 6811 18508 7421 18536
rect 6811 18505 6823 18508
rect 6765 18499 6823 18505
rect 7409 18505 7421 18508
rect 7455 18505 7467 18539
rect 8344 18536 8372 18644
rect 8988 18613 9016 18780
rect 9154 18768 9160 18820
rect 9212 18808 9218 18820
rect 9249 18811 9307 18817
rect 9249 18808 9261 18811
rect 9212 18780 9261 18808
rect 9212 18768 9218 18780
rect 9249 18777 9261 18780
rect 9295 18777 9307 18811
rect 9249 18771 9307 18777
rect 10353 18811 10411 18817
rect 10353 18777 10365 18811
rect 10399 18808 10411 18811
rect 10994 18808 11000 18820
rect 10399 18780 11000 18808
rect 10399 18777 10411 18780
rect 10353 18771 10411 18777
rect 10994 18768 11000 18780
rect 11052 18768 11058 18820
rect 12837 18811 12895 18817
rect 12837 18777 12849 18811
rect 12883 18808 12895 18811
rect 13570 18808 13576 18820
rect 12883 18780 13576 18808
rect 12883 18777 12895 18780
rect 12837 18771 12895 18777
rect 13570 18768 13576 18780
rect 13628 18768 13634 18820
rect 18170 18768 18176 18820
rect 18228 18808 18234 18820
rect 19369 18811 19427 18817
rect 19369 18808 19381 18811
rect 18228 18780 19381 18808
rect 18228 18768 18234 18780
rect 19369 18777 19381 18780
rect 19415 18808 19427 18811
rect 19415 18780 19780 18808
rect 19415 18777 19427 18780
rect 19369 18771 19427 18777
rect 15778 18700 15784 18752
rect 15836 18740 15842 18752
rect 17161 18743 17219 18749
rect 17161 18740 17173 18743
rect 15836 18712 17173 18740
rect 15836 18700 15842 18712
rect 17161 18709 17173 18712
rect 17207 18740 17219 18743
rect 17713 18743 17771 18749
rect 17713 18740 17725 18743
rect 17207 18712 17725 18740
rect 17207 18709 17219 18712
rect 17161 18703 17219 18709
rect 17713 18709 17725 18712
rect 17759 18709 17771 18743
rect 17713 18703 17771 18709
rect 17986 18700 17992 18752
rect 18044 18740 18050 18752
rect 19001 18743 19059 18749
rect 19001 18740 19013 18743
rect 18044 18712 19013 18740
rect 18044 18700 18050 18712
rect 19001 18709 19013 18712
rect 19047 18709 19059 18743
rect 19274 18740 19280 18752
rect 19187 18712 19280 18740
rect 19001 18703 19059 18709
rect 19274 18700 19280 18712
rect 19332 18740 19338 18752
rect 19645 18743 19703 18749
rect 19645 18740 19657 18743
rect 19332 18712 19657 18740
rect 19332 18700 19338 18712
rect 19645 18709 19657 18712
rect 19691 18709 19703 18743
rect 19645 18703 19703 18709
rect 9522 18632 9528 18684
rect 9580 18672 9586 18684
rect 10813 18675 10871 18681
rect 10813 18672 10825 18675
rect 9580 18644 10825 18672
rect 9580 18632 9586 18644
rect 10813 18641 10825 18644
rect 10859 18672 10871 18675
rect 11273 18675 11331 18681
rect 11273 18672 11285 18675
rect 10859 18644 11285 18672
rect 10859 18641 10871 18644
rect 10813 18635 10871 18641
rect 11273 18641 11285 18644
rect 11319 18641 11331 18675
rect 14217 18675 14275 18681
rect 14217 18672 14229 18675
rect 11273 18635 11331 18641
rect 13220 18644 14229 18672
rect 8973 18607 9031 18613
rect 8973 18573 8985 18607
rect 9019 18604 9031 18607
rect 9062 18604 9068 18616
rect 9019 18576 9068 18604
rect 9019 18573 9031 18576
rect 8973 18567 9031 18573
rect 9062 18564 9068 18576
rect 9120 18564 9126 18616
rect 9157 18607 9215 18613
rect 9157 18573 9169 18607
rect 9203 18604 9215 18607
rect 9617 18607 9675 18613
rect 9617 18604 9629 18607
rect 9203 18576 9629 18604
rect 9203 18573 9215 18576
rect 9157 18567 9215 18573
rect 9617 18573 9629 18576
rect 9663 18604 9675 18607
rect 10721 18607 10779 18613
rect 9663 18576 10074 18604
rect 9663 18573 9675 18576
rect 9617 18567 9675 18573
rect 9172 18536 9200 18567
rect 8344 18508 9200 18536
rect 10046 18536 10074 18576
rect 10721 18573 10733 18607
rect 10767 18604 10779 18607
rect 11089 18607 11147 18613
rect 11089 18604 11101 18607
rect 10767 18576 11101 18604
rect 10767 18573 10779 18576
rect 10721 18567 10779 18573
rect 11089 18573 11101 18576
rect 11135 18604 11147 18607
rect 12006 18604 12012 18616
rect 11135 18576 12012 18604
rect 11135 18573 11147 18576
rect 11089 18567 11147 18573
rect 12006 18564 12012 18576
rect 12064 18564 12070 18616
rect 12469 18607 12527 18613
rect 12469 18573 12481 18607
rect 12515 18604 12527 18607
rect 12742 18604 12748 18616
rect 12515 18576 12748 18604
rect 12515 18573 12527 18576
rect 12469 18567 12527 18573
rect 12742 18564 12748 18576
rect 12800 18604 12806 18616
rect 13110 18604 13116 18616
rect 12800 18576 13116 18604
rect 12800 18564 12806 18576
rect 13110 18564 13116 18576
rect 13168 18604 13174 18616
rect 13220 18613 13248 18644
rect 14217 18641 14229 18644
rect 14263 18641 14275 18675
rect 14217 18635 14275 18641
rect 16977 18675 17035 18681
rect 16977 18641 16989 18675
rect 17023 18672 17035 18675
rect 18633 18675 18691 18681
rect 17023 18644 18032 18672
rect 17023 18641 17035 18644
rect 16977 18635 17035 18641
rect 13205 18607 13263 18613
rect 13205 18604 13217 18607
rect 13168 18576 13217 18604
rect 13168 18564 13174 18576
rect 13205 18573 13217 18576
rect 13251 18573 13263 18607
rect 13846 18604 13852 18616
rect 13807 18576 13852 18604
rect 13205 18567 13263 18573
rect 13846 18564 13852 18576
rect 13904 18564 13910 18616
rect 15502 18564 15508 18616
rect 15560 18604 15566 18616
rect 15597 18607 15655 18613
rect 15597 18604 15609 18607
rect 15560 18576 15609 18604
rect 15560 18564 15566 18576
rect 15597 18573 15609 18576
rect 15643 18604 15655 18607
rect 16149 18607 16207 18613
rect 16149 18604 16161 18607
rect 15643 18576 16161 18604
rect 15643 18573 15655 18576
rect 15597 18567 15655 18573
rect 16149 18573 16161 18576
rect 16195 18573 16207 18607
rect 17894 18604 17900 18616
rect 17855 18576 17900 18604
rect 16149 18567 16207 18573
rect 17894 18564 17900 18576
rect 17952 18564 17958 18616
rect 18004 18613 18032 18644
rect 18633 18641 18645 18675
rect 18679 18672 18691 18675
rect 18722 18672 18728 18684
rect 18679 18644 18728 18672
rect 18679 18641 18691 18644
rect 18633 18635 18691 18641
rect 18722 18632 18728 18644
rect 18780 18632 18786 18684
rect 17989 18607 18047 18613
rect 17989 18573 18001 18607
rect 18035 18604 18047 18607
rect 18078 18604 18084 18616
rect 18035 18576 18084 18604
rect 18035 18573 18047 18576
rect 17989 18567 18047 18573
rect 18078 18564 18084 18576
rect 18136 18564 18142 18616
rect 18354 18604 18360 18616
rect 18267 18576 18360 18604
rect 18354 18564 18360 18576
rect 18412 18564 18418 18616
rect 19752 18613 19780 18780
rect 21390 18768 21396 18820
rect 21448 18808 21454 18820
rect 21945 18811 22003 18817
rect 21945 18808 21957 18811
rect 21448 18780 21957 18808
rect 21448 18768 21454 18780
rect 21945 18777 21957 18780
rect 21991 18777 22003 18811
rect 21945 18771 22003 18777
rect 22218 18768 22224 18820
rect 22276 18808 22282 18820
rect 22589 18811 22647 18817
rect 22589 18808 22601 18811
rect 22276 18780 22601 18808
rect 22276 18768 22282 18780
rect 22589 18777 22601 18780
rect 22635 18808 22647 18811
rect 24150 18808 24156 18820
rect 22635 18780 24156 18808
rect 22635 18777 22647 18780
rect 22589 18771 22647 18777
rect 24150 18768 24156 18780
rect 24208 18768 24214 18820
rect 24978 18808 24984 18820
rect 24939 18780 24984 18808
rect 24978 18768 24984 18780
rect 25036 18808 25042 18820
rect 25901 18811 25959 18817
rect 25036 18780 25392 18808
rect 25036 18768 25042 18780
rect 21485 18743 21543 18749
rect 21485 18709 21497 18743
rect 21531 18740 21543 18743
rect 22402 18740 22408 18752
rect 21531 18712 22408 18740
rect 21531 18709 21543 18712
rect 21485 18703 21543 18709
rect 22402 18700 22408 18712
rect 22460 18740 22466 18752
rect 22773 18743 22831 18749
rect 22773 18740 22785 18743
rect 22460 18712 22785 18740
rect 22460 18700 22466 18712
rect 22773 18709 22785 18712
rect 22819 18740 22831 18743
rect 22819 18712 23874 18740
rect 22819 18709 22831 18712
rect 22773 18703 22831 18709
rect 21850 18672 21856 18684
rect 21811 18644 21856 18672
rect 21850 18632 21856 18644
rect 21908 18632 21914 18684
rect 22221 18675 22279 18681
rect 22221 18641 22233 18675
rect 22267 18672 22279 18675
rect 22957 18675 23015 18681
rect 22957 18672 22969 18675
rect 22267 18644 22969 18672
rect 22267 18641 22279 18644
rect 22221 18635 22279 18641
rect 22957 18641 22969 18644
rect 23003 18672 23015 18675
rect 23414 18672 23420 18684
rect 23003 18644 23420 18672
rect 23003 18641 23015 18644
rect 22957 18635 23015 18641
rect 23414 18632 23420 18644
rect 23472 18632 23478 18684
rect 23506 18632 23512 18684
rect 23564 18672 23570 18684
rect 23564 18644 23609 18672
rect 23564 18632 23570 18644
rect 19737 18607 19795 18613
rect 19737 18573 19749 18607
rect 19783 18573 19795 18607
rect 20102 18604 20108 18616
rect 20063 18576 20108 18604
rect 19737 18567 19795 18573
rect 20102 18564 20108 18576
rect 20160 18564 20166 18616
rect 20378 18604 20384 18616
rect 20339 18576 20384 18604
rect 20378 18564 20384 18576
rect 20436 18564 20442 18616
rect 23598 18604 23604 18616
rect 22420 18576 23604 18604
rect 10169 18539 10227 18545
rect 10169 18536 10181 18539
rect 10046 18508 10181 18536
rect 7409 18499 7467 18505
rect 10169 18505 10181 18508
rect 10215 18536 10227 18539
rect 10994 18536 11000 18548
rect 10215 18508 11000 18536
rect 10215 18505 10227 18508
rect 10169 18499 10227 18505
rect 10994 18496 11000 18508
rect 11052 18496 11058 18548
rect 13478 18536 13484 18548
rect 12576 18508 13484 18536
rect 5385 18471 5443 18477
rect 5385 18437 5397 18471
rect 5431 18468 5443 18471
rect 6302 18468 6308 18480
rect 5431 18440 6308 18468
rect 5431 18437 5443 18440
rect 5385 18431 5443 18437
rect 6302 18428 6308 18440
rect 6360 18428 6366 18480
rect 8697 18471 8755 18477
rect 8697 18437 8709 18471
rect 8743 18468 8755 18471
rect 9154 18468 9160 18480
rect 8743 18440 9160 18468
rect 8743 18437 8755 18440
rect 8697 18431 8755 18437
rect 9154 18428 9160 18440
rect 9212 18428 9218 18480
rect 9982 18468 9988 18480
rect 9943 18440 9988 18468
rect 9982 18428 9988 18440
rect 10040 18428 10046 18480
rect 10810 18428 10816 18480
rect 10868 18468 10874 18480
rect 10905 18471 10963 18477
rect 10905 18468 10917 18471
rect 10868 18440 10917 18468
rect 10868 18428 10874 18440
rect 10905 18437 10917 18440
rect 10951 18437 10963 18471
rect 10905 18431 10963 18437
rect 12190 18428 12196 18480
rect 12248 18468 12254 18480
rect 12576 18477 12604 18508
rect 13478 18496 13484 18508
rect 13536 18496 13542 18548
rect 14122 18536 14128 18548
rect 14083 18508 14128 18536
rect 14122 18496 14128 18508
rect 14180 18496 14186 18548
rect 15870 18536 15876 18548
rect 15831 18508 15876 18536
rect 15870 18496 15876 18508
rect 15928 18536 15934 18548
rect 16238 18536 16244 18548
rect 15928 18508 16244 18536
rect 15928 18496 15934 18508
rect 16238 18496 16244 18508
rect 16296 18536 16302 18548
rect 16333 18539 16391 18545
rect 16333 18536 16345 18539
rect 16296 18508 16345 18536
rect 16296 18496 16302 18508
rect 16333 18505 16345 18508
rect 16379 18505 16391 18539
rect 16333 18499 16391 18505
rect 16793 18539 16851 18545
rect 16793 18505 16805 18539
rect 16839 18536 16851 18539
rect 18372 18536 18400 18564
rect 16839 18508 18400 18536
rect 21669 18539 21727 18545
rect 16839 18505 16851 18508
rect 16793 18499 16851 18505
rect 21669 18505 21681 18539
rect 21715 18536 21727 18539
rect 22218 18536 22224 18548
rect 21715 18508 22224 18536
rect 21715 18505 21727 18508
rect 21669 18499 21727 18505
rect 22218 18496 22224 18508
rect 22276 18496 22282 18548
rect 22420 18480 22448 18576
rect 23598 18564 23604 18576
rect 23656 18564 23662 18616
rect 23846 18604 23874 18712
rect 25364 18681 25392 18780
rect 25901 18777 25913 18811
rect 25947 18808 25959 18811
rect 26174 18808 26180 18820
rect 25947 18780 26180 18808
rect 25947 18777 25959 18780
rect 25901 18771 25959 18777
rect 26174 18768 26180 18780
rect 26232 18768 26238 18820
rect 25349 18675 25407 18681
rect 25349 18641 25361 18675
rect 25395 18641 25407 18675
rect 25349 18635 25407 18641
rect 23966 18604 23972 18616
rect 23846 18576 23972 18604
rect 23966 18564 23972 18576
rect 24024 18564 24030 18616
rect 24150 18604 24156 18616
rect 24111 18576 24156 18604
rect 24150 18564 24156 18576
rect 24208 18564 24214 18616
rect 25162 18604 25168 18616
rect 25075 18576 25168 18604
rect 25162 18564 25168 18576
rect 25220 18604 25226 18616
rect 25220 18576 26036 18604
rect 25220 18564 25226 18576
rect 26008 18480 26036 18576
rect 12561 18471 12619 18477
rect 12561 18468 12573 18471
rect 12248 18440 12573 18468
rect 12248 18428 12254 18440
rect 12561 18437 12573 18440
rect 12607 18437 12619 18471
rect 12926 18468 12932 18480
rect 12887 18440 12932 18468
rect 12561 18431 12619 18437
rect 12926 18428 12932 18440
rect 12984 18428 12990 18480
rect 18538 18428 18544 18480
rect 18596 18468 18602 18480
rect 18817 18471 18875 18477
rect 18817 18468 18829 18471
rect 18596 18440 18829 18468
rect 18596 18428 18602 18440
rect 18817 18437 18829 18440
rect 18863 18437 18875 18471
rect 22402 18468 22408 18480
rect 22363 18440 22408 18468
rect 18817 18431 18875 18437
rect 22402 18428 22408 18440
rect 22460 18428 22466 18480
rect 24058 18428 24064 18480
rect 24116 18468 24122 18480
rect 24245 18471 24303 18477
rect 24245 18468 24257 18471
rect 24116 18440 24257 18468
rect 24116 18428 24122 18440
rect 24245 18437 24257 18440
rect 24291 18437 24303 18471
rect 25990 18468 25996 18480
rect 25951 18440 25996 18468
rect 24245 18431 24303 18437
rect 25990 18428 25996 18440
rect 26048 18428 26054 18480
rect 26174 18468 26180 18480
rect 26135 18440 26180 18468
rect 26174 18428 26180 18440
rect 26232 18428 26238 18480
rect 400 18378 27264 18400
rect 400 18326 18870 18378
rect 18922 18326 18934 18378
rect 18986 18326 18998 18378
rect 19050 18326 19062 18378
rect 19114 18326 19126 18378
rect 19178 18326 27264 18378
rect 400 18304 27264 18326
rect 3910 18224 3916 18276
rect 3968 18264 3974 18276
rect 4922 18264 4928 18276
rect 3968 18236 4928 18264
rect 3968 18224 3974 18236
rect 4922 18224 4928 18236
rect 4980 18224 4986 18276
rect 6578 18264 6584 18276
rect 6539 18236 6584 18264
rect 6578 18224 6584 18236
rect 6636 18224 6642 18276
rect 7869 18267 7927 18273
rect 7869 18233 7881 18267
rect 7915 18264 7927 18267
rect 8050 18264 8056 18276
rect 7915 18236 8056 18264
rect 7915 18233 7927 18236
rect 7869 18227 7927 18233
rect 8050 18224 8056 18236
rect 8108 18224 8114 18276
rect 10166 18264 10172 18276
rect 10127 18236 10172 18264
rect 10166 18224 10172 18236
rect 10224 18224 10230 18276
rect 18170 18264 18176 18276
rect 18131 18236 18176 18264
rect 18170 18224 18176 18236
rect 18228 18224 18234 18276
rect 19645 18267 19703 18273
rect 19645 18233 19657 18267
rect 19691 18264 19703 18267
rect 20378 18264 20384 18276
rect 19691 18236 20384 18264
rect 19691 18233 19703 18236
rect 19645 18227 19703 18233
rect 13573 18199 13631 18205
rect 13573 18165 13585 18199
rect 13619 18196 13631 18199
rect 13846 18196 13852 18208
rect 13619 18168 13852 18196
rect 13619 18165 13631 18168
rect 13573 18159 13631 18165
rect 13846 18156 13852 18168
rect 13904 18156 13910 18208
rect 15778 18196 15784 18208
rect 15739 18168 15784 18196
rect 15778 18156 15784 18168
rect 15836 18156 15842 18208
rect 16238 18156 16244 18208
rect 16296 18156 16302 18208
rect 17989 18199 18047 18205
rect 17989 18165 18001 18199
rect 18035 18196 18047 18199
rect 18722 18196 18728 18208
rect 18035 18168 18728 18196
rect 18035 18165 18047 18168
rect 17989 18159 18047 18165
rect 18722 18156 18728 18168
rect 18780 18156 18786 18208
rect 4094 18128 4100 18140
rect 4055 18100 4100 18128
rect 4094 18088 4100 18100
rect 4152 18088 4158 18140
rect 6302 18128 6308 18140
rect 6263 18100 6308 18128
rect 6302 18088 6308 18100
rect 6360 18088 6366 18140
rect 6489 18131 6547 18137
rect 6489 18097 6501 18131
rect 6535 18128 6547 18131
rect 7406 18128 7412 18140
rect 6535 18100 7412 18128
rect 6535 18097 6547 18100
rect 6489 18091 6547 18097
rect 4186 18020 4192 18072
rect 4244 18060 4250 18072
rect 4465 18063 4523 18069
rect 4465 18060 4477 18063
rect 4244 18032 4477 18060
rect 4244 18020 4250 18032
rect 4465 18029 4477 18032
rect 4511 18060 4523 18063
rect 4922 18060 4928 18072
rect 4511 18032 4928 18060
rect 4511 18029 4523 18032
rect 4465 18023 4523 18029
rect 4922 18020 4928 18032
rect 4980 18020 4986 18072
rect 6210 18020 6216 18072
rect 6268 18060 6274 18072
rect 6504 18060 6532 18091
rect 7406 18088 7412 18100
rect 7464 18088 7470 18140
rect 9154 18088 9160 18140
rect 9212 18128 9218 18140
rect 9249 18131 9307 18137
rect 9249 18128 9261 18131
rect 9212 18100 9261 18128
rect 9212 18088 9218 18100
rect 9249 18097 9261 18100
rect 9295 18097 9307 18131
rect 9430 18128 9436 18140
rect 9391 18100 9436 18128
rect 9249 18091 9307 18097
rect 9430 18088 9436 18100
rect 9488 18088 9494 18140
rect 10994 18128 11000 18140
rect 10955 18100 11000 18128
rect 10994 18088 11000 18100
rect 11052 18088 11058 18140
rect 13110 18128 13116 18140
rect 13071 18100 13116 18128
rect 13110 18088 13116 18100
rect 13168 18088 13174 18140
rect 17529 18131 17587 18137
rect 17529 18097 17541 18131
rect 17575 18128 17587 18131
rect 18630 18128 18636 18140
rect 17575 18100 18636 18128
rect 17575 18097 17587 18100
rect 17529 18091 17587 18097
rect 18630 18088 18636 18100
rect 18688 18128 18694 18140
rect 19660 18128 19688 18227
rect 20378 18224 20384 18236
rect 20436 18224 20442 18276
rect 22402 18224 22408 18276
rect 22460 18264 22466 18276
rect 22957 18267 23015 18273
rect 22957 18264 22969 18267
rect 22460 18236 22969 18264
rect 22460 18224 22466 18236
rect 22957 18233 22969 18236
rect 23003 18233 23015 18267
rect 23322 18264 23328 18276
rect 23283 18236 23328 18264
rect 22957 18227 23015 18233
rect 23322 18224 23328 18236
rect 23380 18224 23386 18276
rect 20197 18199 20255 18205
rect 20197 18165 20209 18199
rect 20243 18196 20255 18199
rect 20286 18196 20292 18208
rect 20243 18168 20292 18196
rect 20243 18165 20255 18168
rect 20197 18159 20255 18165
rect 20286 18156 20292 18168
rect 20344 18156 20350 18208
rect 23782 18196 23788 18208
rect 23743 18168 23788 18196
rect 23782 18156 23788 18168
rect 23840 18156 23846 18208
rect 18688 18100 19688 18128
rect 20381 18131 20439 18137
rect 18688 18088 18694 18100
rect 20381 18097 20393 18131
rect 20427 18128 20439 18131
rect 20470 18128 20476 18140
rect 20427 18100 20476 18128
rect 20427 18097 20439 18100
rect 20381 18091 20439 18097
rect 20470 18088 20476 18100
rect 20528 18088 20534 18140
rect 23414 18128 23420 18140
rect 23375 18100 23420 18128
rect 23414 18088 23420 18100
rect 23472 18088 23478 18140
rect 6268 18032 6532 18060
rect 6268 18020 6274 18032
rect 6854 18020 6860 18072
rect 6912 18060 6918 18072
rect 7498 18060 7504 18072
rect 6912 18032 7504 18060
rect 6912 18020 6918 18032
rect 7498 18020 7504 18032
rect 7556 18060 7562 18072
rect 8786 18060 8792 18072
rect 7556 18032 8792 18060
rect 7556 18020 7562 18032
rect 8786 18020 8792 18032
rect 8844 18020 8850 18072
rect 13662 18060 13668 18072
rect 13623 18032 13668 18060
rect 13662 18020 13668 18032
rect 13720 18020 13726 18072
rect 15505 18063 15563 18069
rect 15505 18029 15517 18063
rect 15551 18029 15563 18063
rect 15505 18023 15563 18029
rect 17805 18063 17863 18069
rect 17805 18029 17817 18063
rect 17851 18060 17863 18063
rect 18078 18060 18084 18072
rect 17851 18032 18084 18060
rect 17851 18029 17863 18032
rect 17805 18023 17863 18029
rect 12926 17992 12932 18004
rect 4572 17964 12932 17992
rect 4572 17936 4600 17964
rect 12926 17952 12932 17964
rect 12984 17952 12990 18004
rect 506 17884 512 17936
rect 564 17924 570 17936
rect 693 17927 751 17933
rect 693 17924 705 17927
rect 564 17896 705 17924
rect 564 17884 570 17896
rect 693 17893 705 17896
rect 739 17893 751 17927
rect 693 17887 751 17893
rect 782 17884 788 17936
rect 840 17924 846 17936
rect 877 17927 935 17933
rect 877 17924 889 17927
rect 840 17896 889 17924
rect 840 17884 846 17896
rect 877 17893 889 17896
rect 923 17893 935 17927
rect 877 17887 935 17893
rect 1058 17884 1064 17936
rect 1116 17924 1122 17936
rect 1242 17924 1248 17936
rect 1116 17896 1248 17924
rect 1116 17884 1122 17896
rect 1242 17884 1248 17896
rect 1300 17884 1306 17936
rect 4186 17884 4192 17936
rect 4244 17933 4250 17936
rect 4244 17927 4293 17933
rect 4244 17893 4247 17927
rect 4281 17893 4293 17927
rect 4244 17887 4293 17893
rect 4373 17927 4431 17933
rect 4373 17893 4385 17927
rect 4419 17924 4431 17927
rect 4462 17924 4468 17936
rect 4419 17896 4468 17924
rect 4419 17893 4431 17896
rect 4373 17887 4431 17893
rect 4244 17884 4250 17887
rect 4462 17884 4468 17896
rect 4520 17884 4526 17936
rect 4554 17884 4560 17936
rect 4612 17924 4618 17936
rect 4612 17896 4657 17924
rect 4612 17884 4618 17896
rect 5014 17884 5020 17936
rect 5072 17924 5078 17936
rect 5109 17927 5167 17933
rect 5109 17924 5121 17927
rect 5072 17896 5121 17924
rect 5072 17884 5078 17896
rect 5109 17893 5121 17896
rect 5155 17893 5167 17927
rect 7590 17924 7596 17936
rect 7551 17896 7596 17924
rect 5109 17887 5167 17893
rect 7590 17884 7596 17896
rect 7648 17884 7654 17936
rect 9338 17884 9344 17936
rect 9396 17924 9402 17936
rect 9525 17927 9583 17933
rect 9525 17924 9537 17927
rect 9396 17896 9537 17924
rect 9396 17884 9402 17896
rect 9525 17893 9537 17896
rect 9571 17893 9583 17927
rect 10810 17924 10816 17936
rect 10771 17896 10816 17924
rect 9525 17887 9583 17893
rect 10810 17884 10816 17896
rect 10868 17884 10874 17936
rect 13849 17927 13907 17933
rect 13849 17893 13861 17927
rect 13895 17924 13907 17927
rect 14122 17924 14128 17936
rect 13895 17896 14128 17924
rect 13895 17893 13907 17896
rect 13849 17887 13907 17893
rect 14122 17884 14128 17896
rect 14180 17884 14186 17936
rect 15520 17924 15548 18023
rect 18078 18020 18084 18032
rect 18136 18020 18142 18072
rect 20746 18060 20752 18072
rect 20707 18032 20752 18060
rect 20746 18020 20752 18032
rect 20804 18020 20810 18072
rect 23230 18020 23236 18072
rect 23288 18060 23294 18072
rect 23288 18032 23874 18060
rect 23288 18020 23294 18032
rect 15962 17924 15968 17936
rect 15520 17896 15968 17924
rect 15962 17884 15968 17896
rect 16020 17884 16026 17936
rect 23846 17924 23874 18032
rect 23969 17927 24027 17933
rect 23969 17924 23981 17927
rect 23846 17896 23981 17924
rect 23969 17893 23981 17896
rect 24015 17924 24027 17927
rect 24426 17924 24432 17936
rect 24015 17896 24432 17924
rect 24015 17893 24027 17896
rect 23969 17887 24027 17893
rect 24426 17884 24432 17896
rect 24484 17884 24490 17936
rect 400 17834 27264 17856
rect 400 17782 3510 17834
rect 3562 17782 3574 17834
rect 3626 17782 3638 17834
rect 3690 17782 3702 17834
rect 3754 17782 3766 17834
rect 3818 17782 27264 17834
rect 400 17760 27264 17782
rect 4189 17723 4247 17729
rect 4189 17689 4201 17723
rect 4235 17720 4247 17723
rect 4922 17720 4928 17732
rect 4235 17692 4928 17720
rect 4235 17689 4247 17692
rect 4189 17683 4247 17689
rect 4922 17680 4928 17692
rect 4980 17680 4986 17732
rect 5566 17720 5572 17732
rect 5527 17692 5572 17720
rect 5566 17680 5572 17692
rect 5624 17680 5630 17732
rect 5753 17723 5811 17729
rect 5753 17689 5765 17723
rect 5799 17720 5811 17723
rect 6578 17720 6584 17732
rect 5799 17692 6584 17720
rect 5799 17689 5811 17692
rect 5753 17683 5811 17689
rect 5385 17655 5443 17661
rect 5385 17652 5397 17655
rect 4848 17624 5397 17652
rect 782 17584 788 17596
rect 743 17556 788 17584
rect 782 17544 788 17556
rect 840 17544 846 17596
rect 877 17587 935 17593
rect 877 17553 889 17587
rect 923 17584 935 17587
rect 966 17584 972 17596
rect 923 17556 972 17584
rect 923 17553 935 17556
rect 877 17547 935 17553
rect 966 17544 972 17556
rect 1024 17544 1030 17596
rect 3266 17544 3272 17596
rect 3324 17584 3330 17596
rect 4281 17587 4339 17593
rect 4281 17584 4293 17587
rect 3324 17556 4293 17584
rect 3324 17544 3330 17556
rect 4281 17553 4293 17556
rect 4327 17584 4339 17587
rect 4462 17584 4468 17596
rect 4327 17556 4468 17584
rect 4327 17553 4339 17556
rect 4281 17547 4339 17553
rect 4462 17544 4468 17556
rect 4520 17544 4526 17596
rect 506 17476 512 17528
rect 564 17516 570 17528
rect 1613 17519 1671 17525
rect 1613 17516 1625 17519
rect 564 17488 1625 17516
rect 564 17476 570 17488
rect 1613 17485 1625 17488
rect 1659 17485 1671 17519
rect 1613 17479 1671 17485
rect 1705 17519 1763 17525
rect 1705 17485 1717 17519
rect 1751 17485 1763 17519
rect 1705 17479 1763 17485
rect 3453 17519 3511 17525
rect 3453 17485 3465 17519
rect 3499 17516 3511 17519
rect 4002 17516 4008 17528
rect 3499 17488 4008 17516
rect 3499 17485 3511 17488
rect 3453 17479 3511 17485
rect 690 17408 696 17460
rect 748 17448 754 17460
rect 1720 17448 1748 17479
rect 4002 17476 4008 17488
rect 4060 17516 4066 17528
rect 4738 17516 4744 17528
rect 4060 17488 4744 17516
rect 4060 17476 4066 17488
rect 4738 17476 4744 17488
rect 4796 17476 4802 17528
rect 4848 17525 4876 17624
rect 5385 17621 5397 17624
rect 5431 17652 5443 17655
rect 5768 17652 5796 17683
rect 6578 17680 6584 17692
rect 6636 17680 6642 17732
rect 6854 17720 6860 17732
rect 6815 17692 6860 17720
rect 6854 17680 6860 17692
rect 6912 17680 6918 17732
rect 7314 17680 7320 17732
rect 7372 17720 7378 17732
rect 7777 17723 7835 17729
rect 7777 17720 7789 17723
rect 7372 17692 7789 17720
rect 7372 17680 7378 17692
rect 7777 17689 7789 17692
rect 7823 17720 7835 17723
rect 8421 17723 8479 17729
rect 8421 17720 8433 17723
rect 7823 17692 8433 17720
rect 7823 17689 7835 17692
rect 7777 17683 7835 17689
rect 8421 17689 8433 17692
rect 8467 17689 8479 17723
rect 9798 17720 9804 17732
rect 9759 17692 9804 17720
rect 8421 17683 8479 17689
rect 9798 17680 9804 17692
rect 9856 17680 9862 17732
rect 13110 17720 13116 17732
rect 13071 17692 13116 17720
rect 13110 17680 13116 17692
rect 13168 17680 13174 17732
rect 13573 17723 13631 17729
rect 13573 17689 13585 17723
rect 13619 17720 13631 17723
rect 13846 17720 13852 17732
rect 13619 17692 13852 17720
rect 13619 17689 13631 17692
rect 13573 17683 13631 17689
rect 13846 17680 13852 17692
rect 13904 17680 13910 17732
rect 15781 17723 15839 17729
rect 15781 17689 15793 17723
rect 15827 17720 15839 17723
rect 15870 17720 15876 17732
rect 15827 17692 15876 17720
rect 15827 17689 15839 17692
rect 15781 17683 15839 17689
rect 15870 17680 15876 17692
rect 15928 17680 15934 17732
rect 18449 17723 18507 17729
rect 18449 17689 18461 17723
rect 18495 17720 18507 17723
rect 18722 17720 18728 17732
rect 18495 17692 18728 17720
rect 18495 17689 18507 17692
rect 18449 17683 18507 17689
rect 18722 17680 18728 17692
rect 18780 17680 18786 17732
rect 20289 17723 20347 17729
rect 20289 17689 20301 17723
rect 20335 17720 20347 17723
rect 20470 17720 20476 17732
rect 20335 17692 20476 17720
rect 20335 17689 20347 17692
rect 20289 17683 20347 17689
rect 20470 17680 20476 17692
rect 20528 17680 20534 17732
rect 23414 17680 23420 17732
rect 23472 17720 23478 17732
rect 23785 17723 23843 17729
rect 23785 17720 23797 17723
rect 23472 17692 23797 17720
rect 23472 17680 23478 17692
rect 23785 17689 23797 17692
rect 23831 17689 23843 17723
rect 23785 17683 23843 17689
rect 23966 17680 23972 17732
rect 24024 17720 24030 17732
rect 24245 17723 24303 17729
rect 24245 17720 24257 17723
rect 24024 17692 24257 17720
rect 24024 17680 24030 17692
rect 24245 17689 24257 17692
rect 24291 17720 24303 17723
rect 24613 17723 24671 17729
rect 24613 17720 24625 17723
rect 24291 17692 24625 17720
rect 24291 17689 24303 17692
rect 24245 17683 24303 17689
rect 24613 17689 24625 17692
rect 24659 17689 24671 17723
rect 24613 17683 24671 17689
rect 24889 17723 24947 17729
rect 24889 17689 24901 17723
rect 24935 17720 24947 17723
rect 25806 17720 25812 17732
rect 24935 17692 25812 17720
rect 24935 17689 24947 17692
rect 24889 17683 24947 17689
rect 5431 17624 5796 17652
rect 5431 17621 5443 17624
rect 5385 17615 5443 17621
rect 6394 17612 6400 17664
rect 6452 17652 6458 17664
rect 6872 17652 6900 17680
rect 6452 17624 6900 17652
rect 13389 17655 13447 17661
rect 6452 17612 6458 17624
rect 13389 17621 13401 17655
rect 13435 17652 13447 17655
rect 13662 17652 13668 17664
rect 13435 17624 13668 17652
rect 13435 17621 13447 17624
rect 13389 17615 13447 17621
rect 13662 17612 13668 17624
rect 13720 17652 13726 17664
rect 13941 17655 13999 17661
rect 13941 17652 13953 17655
rect 13720 17624 13953 17652
rect 13720 17612 13726 17624
rect 13941 17621 13953 17624
rect 13987 17652 13999 17655
rect 14217 17655 14275 17661
rect 14217 17652 14229 17655
rect 13987 17624 14229 17652
rect 13987 17621 13999 17624
rect 13941 17615 13999 17621
rect 14217 17621 14229 17624
rect 14263 17621 14275 17655
rect 14217 17615 14275 17621
rect 16149 17655 16207 17661
rect 16149 17621 16161 17655
rect 16195 17652 16207 17655
rect 18630 17652 18636 17664
rect 16195 17624 18636 17652
rect 16195 17621 16207 17624
rect 16149 17615 16207 17621
rect 18630 17612 18636 17624
rect 18688 17612 18694 17664
rect 24150 17652 24156 17664
rect 23616 17624 24156 17652
rect 5937 17587 5995 17593
rect 5937 17553 5949 17587
rect 5983 17584 5995 17587
rect 10169 17587 10227 17593
rect 10169 17584 10181 17587
rect 5983 17556 6716 17584
rect 5983 17553 5995 17556
rect 5937 17547 5995 17553
rect 4833 17519 4891 17525
rect 4833 17485 4845 17519
rect 4879 17485 4891 17519
rect 4833 17479 4891 17485
rect 4922 17476 4928 17528
rect 4980 17516 4986 17528
rect 5952 17516 5980 17547
rect 4980 17488 5980 17516
rect 6305 17519 6363 17525
rect 4980 17476 4986 17488
rect 6305 17485 6317 17519
rect 6351 17516 6363 17519
rect 6394 17516 6400 17528
rect 6351 17488 6400 17516
rect 6351 17485 6363 17488
rect 6305 17479 6363 17485
rect 6394 17476 6400 17488
rect 6452 17476 6458 17528
rect 6688 17525 6716 17556
rect 9724 17556 10181 17584
rect 6673 17519 6731 17525
rect 6673 17485 6685 17519
rect 6719 17516 6731 17519
rect 7130 17516 7136 17528
rect 6719 17488 7136 17516
rect 6719 17485 6731 17488
rect 6673 17479 6731 17485
rect 7130 17476 7136 17488
rect 7188 17516 7194 17528
rect 8050 17516 8056 17528
rect 7188 17488 8056 17516
rect 7188 17476 7194 17488
rect 8050 17476 8056 17488
rect 8108 17476 8114 17528
rect 8329 17519 8387 17525
rect 8329 17485 8341 17519
rect 8375 17516 8387 17519
rect 8375 17488 8924 17516
rect 8375 17485 8387 17488
rect 8329 17479 8387 17485
rect 748 17420 1748 17448
rect 3177 17451 3235 17457
rect 748 17408 754 17420
rect 3177 17417 3189 17451
rect 3223 17448 3235 17451
rect 3269 17451 3327 17457
rect 3269 17448 3281 17451
rect 3223 17420 3281 17448
rect 3223 17417 3235 17420
rect 3177 17411 3235 17417
rect 3269 17417 3281 17420
rect 3315 17448 3327 17451
rect 4649 17451 4707 17457
rect 4649 17448 4661 17451
rect 3315 17420 4661 17448
rect 3315 17417 3327 17420
rect 3269 17411 3327 17417
rect 4649 17417 4661 17420
rect 4695 17448 4707 17451
rect 5566 17448 5572 17460
rect 4695 17420 5572 17448
rect 4695 17417 4707 17420
rect 4649 17411 4707 17417
rect 5566 17408 5572 17420
rect 5624 17408 5630 17460
rect 6118 17448 6124 17460
rect 6031 17420 6124 17448
rect 6118 17408 6124 17420
rect 6176 17448 6182 17460
rect 6854 17448 6860 17460
rect 6176 17420 6860 17448
rect 6176 17408 6182 17420
rect 6854 17408 6860 17420
rect 6912 17448 6918 17460
rect 6949 17451 7007 17457
rect 6949 17448 6961 17451
rect 6912 17420 6961 17448
rect 6912 17408 6918 17420
rect 6949 17417 6961 17420
rect 6995 17417 7007 17451
rect 6949 17411 7007 17417
rect 8145 17451 8203 17457
rect 8145 17417 8157 17451
rect 8191 17417 8203 17451
rect 8145 17411 8203 17417
rect 2622 17340 2628 17392
rect 2680 17380 2686 17392
rect 2993 17383 3051 17389
rect 2993 17380 3005 17383
rect 2680 17352 3005 17380
rect 2680 17340 2686 17352
rect 2993 17349 3005 17352
rect 3039 17380 3051 17383
rect 3545 17383 3603 17389
rect 3545 17380 3557 17383
rect 3039 17352 3557 17380
rect 3039 17349 3051 17352
rect 2993 17343 3051 17349
rect 3545 17349 3557 17352
rect 3591 17349 3603 17383
rect 4002 17380 4008 17392
rect 3963 17352 4008 17380
rect 3545 17343 3603 17349
rect 4002 17340 4008 17352
rect 4060 17340 4066 17392
rect 4370 17340 4376 17392
rect 4428 17380 4434 17392
rect 4557 17383 4615 17389
rect 4557 17380 4569 17383
rect 4428 17352 4569 17380
rect 4428 17340 4434 17352
rect 4557 17349 4569 17352
rect 4603 17380 4615 17383
rect 4925 17383 4983 17389
rect 4925 17380 4937 17383
rect 4603 17352 4937 17380
rect 4603 17349 4615 17352
rect 4557 17343 4615 17349
rect 4925 17349 4937 17352
rect 4971 17349 4983 17383
rect 4925 17343 4983 17349
rect 7225 17383 7283 17389
rect 7225 17349 7237 17383
rect 7271 17380 7283 17383
rect 7406 17380 7412 17392
rect 7271 17352 7412 17380
rect 7271 17349 7283 17352
rect 7225 17343 7283 17349
rect 7406 17340 7412 17352
rect 7464 17340 7470 17392
rect 7958 17380 7964 17392
rect 7919 17352 7964 17380
rect 7958 17340 7964 17352
rect 8016 17380 8022 17392
rect 8160 17380 8188 17411
rect 8896 17389 8924 17488
rect 9246 17476 9252 17528
rect 9304 17516 9310 17528
rect 9724 17525 9752 17556
rect 10169 17553 10181 17556
rect 10215 17553 10227 17587
rect 10169 17547 10227 17553
rect 15597 17587 15655 17593
rect 15597 17553 15609 17587
rect 15643 17584 15655 17587
rect 15778 17584 15784 17596
rect 15643 17556 15784 17584
rect 15643 17553 15655 17556
rect 15597 17547 15655 17553
rect 15778 17544 15784 17556
rect 15836 17544 15842 17596
rect 20286 17544 20292 17596
rect 20344 17584 20350 17596
rect 20381 17587 20439 17593
rect 20381 17584 20393 17587
rect 20344 17556 20393 17584
rect 20344 17544 20350 17556
rect 20381 17553 20393 17556
rect 20427 17553 20439 17587
rect 20381 17547 20439 17553
rect 9709 17519 9767 17525
rect 9709 17516 9721 17519
rect 9304 17488 9721 17516
rect 9304 17476 9310 17488
rect 9709 17485 9721 17488
rect 9755 17485 9767 17519
rect 9709 17479 9767 17485
rect 9890 17476 9896 17528
rect 9948 17516 9954 17528
rect 10810 17516 10816 17528
rect 9948 17488 10816 17516
rect 9948 17476 9954 17488
rect 10810 17476 10816 17488
rect 10868 17516 10874 17528
rect 10905 17519 10963 17525
rect 10905 17516 10917 17519
rect 10868 17488 10917 17516
rect 10868 17476 10874 17488
rect 10905 17485 10917 17488
rect 10951 17485 10963 17519
rect 14122 17516 14128 17528
rect 14083 17488 14128 17516
rect 10905 17479 10963 17485
rect 14122 17476 14128 17488
rect 14180 17516 14186 17528
rect 14401 17519 14459 17525
rect 14401 17516 14413 17519
rect 14180 17488 14413 17516
rect 14180 17476 14186 17488
rect 14401 17485 14413 17488
rect 14447 17485 14459 17519
rect 14401 17479 14459 17485
rect 20105 17519 20163 17525
rect 20105 17485 20117 17519
rect 20151 17516 20163 17519
rect 20746 17516 20752 17528
rect 20151 17488 20752 17516
rect 20151 17485 20163 17488
rect 20105 17479 20163 17485
rect 20746 17476 20752 17488
rect 20804 17516 20810 17528
rect 21114 17516 21120 17528
rect 20804 17488 21120 17516
rect 20804 17476 20810 17488
rect 21114 17476 21120 17488
rect 21172 17476 21178 17528
rect 22773 17519 22831 17525
rect 22773 17485 22785 17519
rect 22819 17516 22831 17519
rect 23233 17519 23291 17525
rect 23233 17516 23245 17519
rect 22819 17488 23245 17516
rect 22819 17485 22831 17488
rect 22773 17479 22831 17485
rect 23233 17485 23245 17488
rect 23279 17516 23291 17519
rect 23506 17516 23512 17528
rect 23279 17488 23512 17516
rect 23279 17485 23291 17488
rect 23233 17479 23291 17485
rect 23506 17476 23512 17488
rect 23564 17476 23570 17528
rect 9154 17448 9160 17460
rect 9067 17420 9160 17448
rect 9154 17408 9160 17420
rect 9212 17448 9218 17460
rect 9525 17451 9583 17457
rect 9525 17448 9537 17451
rect 9212 17420 9537 17448
rect 9212 17408 9218 17420
rect 9525 17417 9537 17420
rect 9571 17448 9583 17451
rect 9982 17448 9988 17460
rect 9571 17420 9988 17448
rect 9571 17417 9583 17420
rect 9525 17411 9583 17417
rect 9982 17408 9988 17420
rect 10040 17448 10046 17460
rect 10353 17451 10411 17457
rect 10353 17448 10365 17451
rect 10040 17420 10365 17448
rect 10040 17408 10046 17420
rect 10353 17417 10365 17420
rect 10399 17417 10411 17451
rect 10353 17411 10411 17417
rect 13846 17408 13852 17460
rect 13904 17448 13910 17460
rect 14582 17448 14588 17460
rect 13904 17420 14588 17448
rect 13904 17408 13910 17420
rect 14582 17408 14588 17420
rect 14640 17408 14646 17460
rect 21022 17448 21028 17460
rect 20935 17420 21028 17448
rect 21022 17408 21028 17420
rect 21080 17448 21086 17460
rect 23616 17457 23644 17624
rect 24150 17612 24156 17624
rect 24208 17612 24214 17664
rect 23690 17476 23696 17528
rect 23748 17516 23754 17528
rect 24058 17516 24064 17528
rect 23748 17488 24064 17516
rect 23748 17476 23754 17488
rect 24058 17476 24064 17488
rect 24116 17476 24122 17528
rect 24426 17516 24432 17528
rect 24339 17488 24432 17516
rect 24426 17476 24432 17488
rect 24484 17516 24490 17528
rect 24904 17516 24932 17683
rect 25806 17680 25812 17692
rect 25864 17680 25870 17732
rect 24484 17488 24932 17516
rect 24484 17476 24490 17488
rect 21301 17451 21359 17457
rect 21301 17448 21313 17451
rect 21080 17420 21313 17448
rect 21080 17408 21086 17420
rect 21301 17417 21313 17420
rect 21347 17417 21359 17451
rect 21301 17411 21359 17417
rect 23325 17451 23383 17457
rect 23325 17417 23337 17451
rect 23371 17448 23383 17451
rect 23601 17451 23659 17457
rect 23601 17448 23613 17451
rect 23371 17420 23613 17448
rect 23371 17417 23383 17420
rect 23325 17411 23383 17417
rect 23601 17417 23613 17420
rect 23647 17417 23659 17451
rect 23601 17411 23659 17417
rect 8016 17352 8188 17380
rect 8881 17383 8939 17389
rect 8016 17340 8022 17352
rect 8881 17349 8893 17383
rect 8927 17380 8939 17383
rect 9341 17383 9399 17389
rect 9341 17380 9353 17383
rect 8927 17352 9353 17380
rect 8927 17349 8939 17352
rect 8881 17343 8939 17349
rect 9341 17349 9353 17352
rect 9387 17380 9399 17383
rect 9430 17380 9436 17392
rect 9387 17352 9436 17380
rect 9387 17349 9399 17352
rect 9341 17343 9399 17349
rect 9430 17340 9436 17352
rect 9488 17340 9494 17392
rect 10813 17383 10871 17389
rect 10813 17349 10825 17383
rect 10859 17380 10871 17383
rect 10994 17380 11000 17392
rect 10859 17352 11000 17380
rect 10859 17349 10871 17352
rect 10813 17343 10871 17349
rect 10994 17340 11000 17352
rect 11052 17380 11058 17392
rect 12190 17380 12196 17392
rect 11052 17352 12196 17380
rect 11052 17340 11058 17352
rect 12190 17340 12196 17352
rect 12248 17340 12254 17392
rect 15962 17380 15968 17392
rect 15923 17352 15968 17380
rect 15962 17340 15968 17352
rect 16020 17340 16026 17392
rect 23509 17383 23567 17389
rect 23509 17349 23521 17383
rect 23555 17380 23567 17383
rect 23782 17380 23788 17392
rect 23555 17352 23788 17380
rect 23555 17349 23567 17352
rect 23509 17343 23567 17349
rect 23782 17340 23788 17352
rect 23840 17340 23846 17392
rect 400 17290 27264 17312
rect 400 17238 18870 17290
rect 18922 17238 18934 17290
rect 18986 17238 18998 17290
rect 19050 17238 19062 17290
rect 19114 17238 19126 17290
rect 19178 17238 27264 17290
rect 400 17216 27264 17238
rect 966 17176 972 17188
rect 927 17148 972 17176
rect 966 17136 972 17148
rect 1024 17136 1030 17188
rect 2622 17176 2628 17188
rect 2583 17148 2628 17176
rect 2622 17136 2628 17148
rect 2680 17136 2686 17188
rect 4094 17136 4100 17188
rect 4152 17176 4158 17188
rect 4281 17179 4339 17185
rect 4281 17176 4293 17179
rect 4152 17148 4293 17176
rect 4152 17136 4158 17148
rect 4281 17145 4293 17148
rect 4327 17145 4339 17179
rect 4281 17139 4339 17145
rect 4554 17136 4560 17188
rect 4612 17176 4618 17188
rect 9338 17176 9344 17188
rect 4612 17148 4657 17176
rect 9299 17148 9344 17176
rect 4612 17136 4618 17148
rect 9338 17136 9344 17148
rect 9396 17136 9402 17188
rect 14582 17176 14588 17188
rect 14543 17148 14588 17176
rect 14582 17136 14588 17148
rect 14640 17136 14646 17188
rect 1702 17108 1708 17120
rect 1663 17080 1708 17108
rect 1702 17068 1708 17080
rect 1760 17068 1766 17120
rect 5477 17111 5535 17117
rect 5477 17077 5489 17111
rect 5523 17108 5535 17111
rect 5750 17108 5756 17120
rect 5523 17080 5756 17108
rect 5523 17077 5535 17080
rect 5477 17071 5535 17077
rect 5750 17068 5756 17080
rect 5808 17108 5814 17120
rect 5808 17080 7084 17108
rect 5808 17068 5814 17080
rect 5566 17000 5572 17052
rect 5624 17040 5630 17052
rect 5661 17043 5719 17049
rect 5661 17040 5673 17043
rect 5624 17012 5673 17040
rect 5624 17000 5630 17012
rect 5661 17009 5673 17012
rect 5707 17040 5719 17043
rect 6118 17040 6124 17052
rect 5707 17012 6124 17040
rect 5707 17009 5719 17012
rect 5661 17003 5719 17009
rect 6118 17000 6124 17012
rect 6176 17000 6182 17052
rect 6857 17043 6915 17049
rect 6857 17009 6869 17043
rect 6903 17040 6915 17043
rect 6946 17040 6952 17052
rect 6903 17012 6952 17040
rect 6903 17009 6915 17012
rect 6857 17003 6915 17009
rect 6946 17000 6952 17012
rect 7004 17000 7010 17052
rect 7056 17049 7084 17080
rect 20470 17068 20476 17120
rect 20528 17108 20534 17120
rect 21482 17108 21488 17120
rect 20528 17080 21488 17108
rect 20528 17068 20534 17080
rect 7041 17043 7099 17049
rect 7041 17009 7053 17043
rect 7087 17009 7099 17043
rect 7041 17003 7099 17009
rect 10258 17000 10264 17052
rect 10316 17040 10322 17052
rect 11549 17043 11607 17049
rect 11549 17040 11561 17043
rect 10316 17012 11561 17040
rect 10316 17000 10322 17012
rect 11549 17009 11561 17012
rect 11595 17009 11607 17043
rect 11549 17003 11607 17009
rect 12190 17000 12196 17052
rect 12248 17040 12254 17052
rect 12293 17043 12351 17049
rect 12293 17040 12305 17043
rect 12248 17012 12305 17040
rect 12248 17000 12254 17012
rect 12293 17009 12305 17012
rect 12339 17009 12351 17043
rect 12293 17003 12351 17009
rect 15134 17000 15140 17052
rect 15192 17040 15198 17052
rect 15781 17043 15839 17049
rect 15781 17040 15793 17043
rect 15192 17012 15793 17040
rect 15192 17000 15198 17012
rect 15781 17009 15793 17012
rect 15827 17009 15839 17043
rect 15781 17003 15839 17009
rect 16333 17043 16391 17049
rect 16333 17009 16345 17043
rect 16379 17040 16391 17043
rect 16422 17040 16428 17052
rect 16379 17012 16428 17040
rect 16379 17009 16391 17012
rect 16333 17003 16391 17009
rect 16422 17000 16428 17012
rect 16480 17000 16486 17052
rect 20654 17000 20660 17052
rect 20712 17040 20718 17052
rect 20948 17049 20976 17080
rect 21482 17068 21488 17080
rect 21540 17068 21546 17120
rect 20841 17043 20899 17049
rect 20841 17040 20853 17043
rect 20712 17012 20853 17040
rect 20712 17000 20718 17012
rect 20841 17009 20853 17012
rect 20887 17009 20899 17043
rect 20841 17003 20899 17009
rect 20933 17043 20991 17049
rect 20933 17009 20945 17043
rect 20979 17009 20991 17043
rect 21206 17040 21212 17052
rect 21167 17012 21212 17040
rect 20933 17003 20991 17009
rect 21206 17000 21212 17012
rect 21264 17000 21270 17052
rect 24334 17000 24340 17052
rect 24392 17040 24398 17052
rect 25809 17043 25867 17049
rect 25809 17040 25821 17043
rect 24392 17012 25821 17040
rect 24392 17000 24398 17012
rect 25809 17009 25821 17012
rect 25855 17040 25867 17043
rect 26450 17040 26456 17052
rect 25855 17012 26456 17040
rect 25855 17009 25867 17012
rect 25809 17003 25867 17009
rect 26450 17000 26456 17012
rect 26508 17000 26514 17052
rect 1242 16932 1248 16984
rect 1300 16972 1306 16984
rect 2073 16975 2131 16981
rect 2073 16972 2085 16975
rect 1300 16944 2085 16972
rect 1300 16932 1306 16944
rect 2073 16941 2085 16944
rect 2119 16972 2131 16975
rect 4097 16975 4155 16981
rect 4097 16972 4109 16975
rect 2119 16944 4109 16972
rect 2119 16941 2131 16944
rect 2073 16935 2131 16941
rect 4097 16941 4109 16944
rect 4143 16972 4155 16975
rect 4186 16972 4192 16984
rect 4143 16944 4192 16972
rect 4143 16941 4155 16944
rect 4097 16935 4155 16941
rect 4186 16932 4192 16944
rect 4244 16932 4250 16984
rect 7958 16932 7964 16984
rect 8016 16972 8022 16984
rect 9525 16975 9583 16981
rect 9525 16972 9537 16975
rect 8016 16944 9537 16972
rect 8016 16932 8022 16944
rect 9525 16941 9537 16944
rect 9571 16972 9583 16975
rect 9798 16972 9804 16984
rect 9571 16944 9804 16972
rect 9571 16941 9583 16944
rect 9525 16935 9583 16941
rect 9798 16932 9804 16944
rect 9856 16972 9862 16984
rect 10902 16972 10908 16984
rect 9856 16944 10908 16972
rect 9856 16932 9862 16944
rect 10902 16932 10908 16944
rect 10960 16972 10966 16984
rect 11457 16975 11515 16981
rect 11457 16972 11469 16975
rect 10960 16944 11469 16972
rect 10960 16932 10966 16944
rect 11457 16941 11469 16944
rect 11503 16941 11515 16975
rect 12374 16972 12380 16984
rect 12335 16944 12380 16972
rect 11457 16935 11515 16941
rect 12374 16932 12380 16944
rect 12432 16932 12438 16984
rect 16517 16975 16575 16981
rect 16517 16941 16529 16975
rect 16563 16972 16575 16975
rect 16698 16972 16704 16984
rect 16563 16944 16704 16972
rect 16563 16941 16575 16944
rect 16517 16935 16575 16941
rect 16698 16932 16704 16944
rect 16756 16932 16762 16984
rect 21114 16932 21120 16984
rect 21172 16972 21178 16984
rect 21301 16975 21359 16981
rect 21301 16972 21313 16975
rect 21172 16944 21313 16972
rect 21172 16932 21178 16944
rect 21301 16941 21313 16944
rect 21347 16941 21359 16975
rect 21301 16935 21359 16941
rect 782 16864 788 16916
rect 840 16904 846 16916
rect 2165 16907 2223 16913
rect 2165 16904 2177 16907
rect 840 16876 2177 16904
rect 840 16864 846 16876
rect 2165 16873 2177 16876
rect 2211 16873 2223 16907
rect 2165 16867 2223 16873
rect 2530 16864 2536 16916
rect 2588 16904 2594 16916
rect 6210 16904 6216 16916
rect 2588 16876 6216 16904
rect 2588 16864 2594 16876
rect 6210 16864 6216 16876
rect 6268 16864 6274 16916
rect 6302 16864 6308 16916
rect 6360 16904 6366 16916
rect 6397 16907 6455 16913
rect 6397 16904 6409 16907
rect 6360 16876 6409 16904
rect 6360 16864 6366 16876
rect 6397 16873 6409 16876
rect 6443 16904 6455 16907
rect 11546 16904 11552 16916
rect 6443 16876 11552 16904
rect 6443 16873 6455 16876
rect 6397 16867 6455 16873
rect 11546 16864 11552 16876
rect 11604 16864 11610 16916
rect 23049 16907 23107 16913
rect 23049 16873 23061 16907
rect 23095 16904 23107 16907
rect 23230 16904 23236 16916
rect 23095 16876 23236 16904
rect 23095 16873 23107 16876
rect 23049 16867 23107 16873
rect 23230 16864 23236 16876
rect 23288 16864 23294 16916
rect 690 16836 696 16848
rect 651 16808 696 16836
rect 690 16796 696 16808
rect 748 16796 754 16848
rect 1702 16796 1708 16848
rect 1760 16836 1766 16848
rect 1843 16839 1901 16845
rect 1843 16836 1855 16839
rect 1760 16808 1855 16836
rect 1760 16796 1766 16808
rect 1843 16805 1855 16808
rect 1889 16805 1901 16839
rect 1843 16799 1901 16805
rect 1981 16839 2039 16845
rect 1981 16805 1993 16839
rect 2027 16836 2039 16839
rect 2622 16836 2628 16848
rect 2027 16808 2628 16836
rect 2027 16805 2039 16808
rect 1981 16799 2039 16805
rect 2622 16796 2628 16808
rect 2680 16796 2686 16848
rect 5658 16796 5664 16848
rect 5716 16836 5722 16848
rect 5753 16839 5811 16845
rect 5753 16836 5765 16839
rect 5716 16808 5765 16836
rect 5716 16796 5722 16808
rect 5753 16805 5765 16808
rect 5799 16805 5811 16839
rect 5753 16799 5811 16805
rect 7133 16839 7191 16845
rect 7133 16805 7145 16839
rect 7179 16836 7191 16839
rect 7222 16836 7228 16848
rect 7179 16808 7228 16836
rect 7179 16805 7191 16808
rect 7133 16799 7191 16805
rect 7222 16796 7228 16808
rect 7280 16796 7286 16848
rect 8421 16839 8479 16845
rect 8421 16805 8433 16839
rect 8467 16836 8479 16839
rect 8602 16836 8608 16848
rect 8467 16808 8608 16836
rect 8467 16805 8479 16808
rect 8421 16799 8479 16805
rect 8602 16796 8608 16808
rect 8660 16796 8666 16848
rect 14674 16836 14680 16848
rect 14635 16808 14680 16836
rect 14674 16796 14680 16808
rect 14732 16796 14738 16848
rect 15410 16836 15416 16848
rect 15371 16808 15416 16836
rect 15410 16796 15416 16808
rect 15468 16796 15474 16848
rect 17802 16836 17808 16848
rect 17763 16808 17808 16836
rect 17802 16796 17808 16808
rect 17860 16796 17866 16848
rect 20286 16836 20292 16848
rect 20247 16808 20292 16836
rect 20286 16796 20292 16808
rect 20344 16796 20350 16848
rect 23138 16836 23144 16848
rect 23099 16808 23144 16836
rect 23138 16796 23144 16808
rect 23196 16796 23202 16848
rect 24978 16836 24984 16848
rect 24939 16808 24984 16836
rect 24978 16796 24984 16808
rect 25036 16796 25042 16848
rect 25993 16839 26051 16845
rect 25993 16805 26005 16839
rect 26039 16836 26051 16839
rect 26358 16836 26364 16848
rect 26039 16808 26364 16836
rect 26039 16805 26051 16808
rect 25993 16799 26051 16805
rect 26358 16796 26364 16808
rect 26416 16796 26422 16848
rect 400 16746 27264 16768
rect 400 16694 3510 16746
rect 3562 16694 3574 16746
rect 3626 16694 3638 16746
rect 3690 16694 3702 16746
rect 3754 16694 3766 16746
rect 3818 16694 27264 16746
rect 400 16672 27264 16694
rect 782 16592 788 16644
rect 840 16632 846 16644
rect 1153 16635 1211 16641
rect 1153 16632 1165 16635
rect 840 16604 1165 16632
rect 840 16592 846 16604
rect 1153 16601 1165 16604
rect 1199 16601 1211 16635
rect 1794 16632 1800 16644
rect 1755 16604 1800 16632
rect 1153 16595 1211 16601
rect 1794 16592 1800 16604
rect 1852 16592 1858 16644
rect 2257 16635 2315 16641
rect 2257 16601 2269 16635
rect 2303 16632 2315 16635
rect 2625 16635 2683 16641
rect 2625 16632 2637 16635
rect 2303 16604 2637 16632
rect 2303 16601 2315 16604
rect 2257 16595 2315 16601
rect 2625 16601 2637 16604
rect 2671 16632 2683 16635
rect 3266 16632 3272 16644
rect 2671 16604 3272 16632
rect 2671 16601 2683 16604
rect 2625 16595 2683 16601
rect 3266 16592 3272 16604
rect 3324 16592 3330 16644
rect 3545 16635 3603 16641
rect 3545 16601 3557 16635
rect 3591 16632 3603 16635
rect 4094 16632 4100 16644
rect 3591 16604 4100 16632
rect 3591 16601 3603 16604
rect 3545 16595 3603 16601
rect 4094 16592 4100 16604
rect 4152 16632 4158 16644
rect 4465 16635 4523 16641
rect 4465 16632 4477 16635
rect 4152 16604 4477 16632
rect 4152 16592 4158 16604
rect 4465 16601 4477 16604
rect 4511 16601 4523 16635
rect 5566 16632 5572 16644
rect 5527 16604 5572 16632
rect 4465 16595 4523 16601
rect 5566 16592 5572 16604
rect 5624 16592 5630 16644
rect 5658 16592 5664 16644
rect 5716 16632 5722 16644
rect 5845 16635 5903 16641
rect 5845 16632 5857 16635
rect 5716 16604 5857 16632
rect 5716 16592 5722 16604
rect 5845 16601 5857 16604
rect 5891 16601 5903 16635
rect 5845 16595 5903 16601
rect 6946 16592 6952 16644
rect 7004 16632 7010 16644
rect 7041 16635 7099 16641
rect 7041 16632 7053 16635
rect 7004 16604 7053 16632
rect 7004 16592 7010 16604
rect 7041 16601 7053 16604
rect 7087 16601 7099 16635
rect 7041 16595 7099 16601
rect 8970 16592 8976 16644
rect 9028 16632 9034 16644
rect 9157 16635 9215 16641
rect 9157 16632 9169 16635
rect 9028 16604 9169 16632
rect 9028 16592 9034 16604
rect 9157 16601 9169 16604
rect 9203 16601 9215 16635
rect 9157 16595 9215 16601
rect 11089 16635 11147 16641
rect 11089 16601 11101 16635
rect 11135 16632 11147 16635
rect 12374 16632 12380 16644
rect 11135 16604 12380 16632
rect 11135 16601 11147 16604
rect 11089 16595 11147 16601
rect 12374 16592 12380 16604
rect 12432 16592 12438 16644
rect 14582 16632 14588 16644
rect 14543 16604 14588 16632
rect 14582 16592 14588 16604
rect 14640 16592 14646 16644
rect 14674 16592 14680 16644
rect 14732 16632 14738 16644
rect 14769 16635 14827 16641
rect 14769 16632 14781 16635
rect 14732 16604 14781 16632
rect 14732 16592 14738 16604
rect 14769 16601 14781 16604
rect 14815 16601 14827 16635
rect 15134 16632 15140 16644
rect 15095 16604 15140 16632
rect 14769 16595 14827 16601
rect 15134 16592 15140 16604
rect 15192 16592 15198 16644
rect 20470 16632 20476 16644
rect 20431 16604 20476 16632
rect 20470 16592 20476 16604
rect 20528 16592 20534 16644
rect 20654 16632 20660 16644
rect 20615 16604 20660 16632
rect 20654 16592 20660 16604
rect 20712 16592 20718 16644
rect 20841 16635 20899 16641
rect 20841 16601 20853 16635
rect 20887 16632 20899 16635
rect 21114 16632 21120 16644
rect 20887 16604 21120 16632
rect 20887 16601 20899 16604
rect 20841 16595 20899 16601
rect 21114 16592 21120 16604
rect 21172 16592 21178 16644
rect 22773 16635 22831 16641
rect 22773 16601 22785 16635
rect 22819 16632 22831 16635
rect 24058 16632 24064 16644
rect 22819 16604 24064 16632
rect 22819 16601 22831 16604
rect 22773 16595 22831 16601
rect 24058 16592 24064 16604
rect 24116 16632 24122 16644
rect 24797 16635 24855 16641
rect 24797 16632 24809 16635
rect 24116 16604 24809 16632
rect 24116 16592 24122 16604
rect 24797 16601 24809 16604
rect 24843 16601 24855 16635
rect 26450 16632 26456 16644
rect 26411 16604 26456 16632
rect 24797 16595 24855 16601
rect 3910 16564 3916 16576
rect 3871 16536 3916 16564
rect 3910 16524 3916 16536
rect 3968 16524 3974 16576
rect 4278 16564 4284 16576
rect 4239 16536 4284 16564
rect 4278 16524 4284 16536
rect 4336 16524 4342 16576
rect 4925 16567 4983 16573
rect 4925 16533 4937 16567
rect 4971 16564 4983 16567
rect 5934 16564 5940 16576
rect 4971 16536 5940 16564
rect 4971 16533 4983 16536
rect 4925 16527 4983 16533
rect 2530 16505 2536 16508
rect 1889 16499 1947 16505
rect 1889 16465 1901 16499
rect 1935 16496 1947 16499
rect 2496 16499 2536 16505
rect 2496 16496 2508 16499
rect 1935 16468 2508 16496
rect 1935 16465 1947 16468
rect 1889 16459 1947 16465
rect 2496 16465 2508 16468
rect 2496 16459 2536 16465
rect 2530 16456 2536 16459
rect 2588 16456 2594 16508
rect 2717 16499 2775 16505
rect 2717 16465 2729 16499
rect 2763 16496 2775 16499
rect 3177 16499 3235 16505
rect 3177 16496 3189 16499
rect 2763 16468 3189 16496
rect 2763 16465 2775 16468
rect 2717 16459 2775 16465
rect 3177 16465 3189 16468
rect 3223 16496 3235 16499
rect 3358 16496 3364 16508
rect 3223 16468 3364 16496
rect 3223 16465 3235 16468
rect 3177 16459 3235 16465
rect 3358 16456 3364 16468
rect 3416 16456 3422 16508
rect 3729 16499 3787 16505
rect 3729 16465 3741 16499
rect 3775 16496 3787 16499
rect 4373 16499 4431 16505
rect 4373 16496 4385 16499
rect 3775 16468 4385 16496
rect 3775 16465 3787 16468
rect 3729 16459 3787 16465
rect 4373 16465 4385 16468
rect 4419 16465 4431 16499
rect 4373 16459 4431 16465
rect 1429 16431 1487 16437
rect 1429 16397 1441 16431
rect 1475 16428 1487 16431
rect 2349 16431 2407 16437
rect 2349 16428 2361 16431
rect 1475 16400 2361 16428
rect 1475 16397 1487 16400
rect 1429 16391 1487 16397
rect 2349 16397 2361 16400
rect 2395 16428 2407 16431
rect 2622 16428 2628 16440
rect 2395 16400 2628 16428
rect 2395 16397 2407 16400
rect 2349 16391 2407 16397
rect 2622 16388 2628 16400
rect 2680 16388 2686 16440
rect 3266 16388 3272 16440
rect 3324 16428 3330 16440
rect 3744 16428 3772 16459
rect 3324 16400 3772 16428
rect 3324 16388 3330 16400
rect 3910 16388 3916 16440
rect 3968 16428 3974 16440
rect 4005 16431 4063 16437
rect 4005 16428 4017 16431
rect 3968 16400 4017 16428
rect 3968 16388 3974 16400
rect 4005 16397 4017 16400
rect 4051 16397 4063 16431
rect 4005 16391 4063 16397
rect 4152 16431 4210 16437
rect 4152 16397 4164 16431
rect 4198 16428 4210 16431
rect 4940 16428 4968 16527
rect 5934 16524 5940 16536
rect 5992 16564 5998 16576
rect 7222 16564 7228 16576
rect 5992 16536 7228 16564
rect 5992 16524 5998 16536
rect 7222 16524 7228 16536
rect 7280 16524 7286 16576
rect 15045 16567 15103 16573
rect 15045 16533 15057 16567
rect 15091 16564 15103 16567
rect 15091 16536 16376 16564
rect 15091 16533 15103 16536
rect 15045 16527 15103 16533
rect 9062 16496 9068 16508
rect 9023 16468 9068 16496
rect 9062 16456 9068 16468
rect 9120 16456 9126 16508
rect 11178 16456 11184 16508
rect 11236 16496 11242 16508
rect 12745 16499 12803 16505
rect 12745 16496 12757 16499
rect 11236 16468 12757 16496
rect 11236 16456 11242 16468
rect 12745 16465 12757 16468
rect 12791 16465 12803 16499
rect 15410 16496 15416 16508
rect 15371 16468 15416 16496
rect 12745 16459 12803 16465
rect 15410 16456 15416 16468
rect 15468 16456 15474 16508
rect 16348 16505 16376 16536
rect 17802 16524 17808 16576
rect 17860 16564 17866 16576
rect 19001 16567 19059 16573
rect 19001 16564 19013 16567
rect 17860 16536 19013 16564
rect 17860 16524 17866 16536
rect 19001 16533 19013 16536
rect 19047 16533 19059 16567
rect 19001 16527 19059 16533
rect 20289 16567 20347 16573
rect 20289 16533 20301 16567
rect 20335 16564 20347 16567
rect 21025 16567 21083 16573
rect 21025 16564 21037 16567
rect 20335 16536 21037 16564
rect 20335 16533 20347 16536
rect 20289 16527 20347 16533
rect 21025 16533 21037 16536
rect 21071 16564 21083 16567
rect 21206 16564 21212 16576
rect 21071 16536 21212 16564
rect 21071 16533 21083 16536
rect 21025 16527 21083 16533
rect 21206 16524 21212 16536
rect 21264 16564 21270 16576
rect 21577 16567 21635 16573
rect 21577 16564 21589 16567
rect 21264 16536 21589 16564
rect 21264 16524 21270 16536
rect 21577 16533 21589 16536
rect 21623 16533 21635 16567
rect 23138 16564 23144 16576
rect 21577 16527 21635 16533
rect 21684 16536 23144 16564
rect 16333 16499 16391 16505
rect 16333 16465 16345 16499
rect 16379 16496 16391 16499
rect 16422 16496 16428 16508
rect 16379 16468 16428 16496
rect 16379 16465 16391 16468
rect 16333 16459 16391 16465
rect 16422 16456 16428 16468
rect 16480 16456 16486 16508
rect 21684 16496 21712 16536
rect 23138 16524 23144 16536
rect 23196 16564 23202 16576
rect 23233 16567 23291 16573
rect 23233 16564 23245 16567
rect 23196 16536 23245 16564
rect 23196 16524 23202 16536
rect 23233 16533 23245 16536
rect 23279 16533 23291 16567
rect 24812 16564 24840 16595
rect 26450 16592 26456 16604
rect 26508 16592 26514 16644
rect 26358 16564 26364 16576
rect 24812 16536 25944 16564
rect 26319 16536 26364 16564
rect 23233 16527 23291 16533
rect 19016 16468 21712 16496
rect 22405 16499 22463 16505
rect 4198 16400 4968 16428
rect 4198 16397 4210 16400
rect 4152 16391 4210 16397
rect 5474 16388 5480 16440
rect 5532 16428 5538 16440
rect 7961 16431 8019 16437
rect 7961 16428 7973 16431
rect 5532 16400 7973 16428
rect 5532 16388 5538 16400
rect 7961 16397 7973 16400
rect 8007 16428 8019 16431
rect 8513 16431 8571 16437
rect 8513 16428 8525 16431
rect 8007 16400 8525 16428
rect 8007 16397 8019 16400
rect 7961 16391 8019 16397
rect 8513 16397 8525 16400
rect 8559 16397 8571 16431
rect 11822 16428 11828 16440
rect 11783 16400 11828 16428
rect 8513 16391 8571 16397
rect 11822 16388 11828 16400
rect 11880 16388 11886 16440
rect 12653 16431 12711 16437
rect 12653 16397 12665 16431
rect 12699 16428 12711 16431
rect 13110 16428 13116 16440
rect 12699 16400 13116 16428
rect 12699 16397 12711 16400
rect 12653 16391 12711 16397
rect 13110 16388 13116 16400
rect 13168 16388 13174 16440
rect 15134 16388 15140 16440
rect 15192 16428 15198 16440
rect 16241 16431 16299 16437
rect 16241 16428 16253 16431
rect 15192 16400 16253 16428
rect 15192 16388 15198 16400
rect 16241 16397 16253 16400
rect 16287 16428 16299 16431
rect 16517 16431 16575 16437
rect 16517 16428 16529 16431
rect 16287 16400 16529 16428
rect 16287 16397 16299 16400
rect 16241 16391 16299 16397
rect 16517 16397 16529 16400
rect 16563 16428 16575 16431
rect 17158 16428 17164 16440
rect 16563 16400 17164 16428
rect 16563 16397 16575 16400
rect 16517 16391 16575 16397
rect 17158 16388 17164 16400
rect 17216 16388 17222 16440
rect 17621 16431 17679 16437
rect 17621 16397 17633 16431
rect 17667 16428 17679 16431
rect 18538 16428 18544 16440
rect 17667 16400 18544 16428
rect 17667 16397 17679 16400
rect 17621 16391 17679 16397
rect 18538 16388 18544 16400
rect 18596 16428 18602 16440
rect 18725 16431 18783 16437
rect 18725 16428 18737 16431
rect 18596 16400 18737 16428
rect 18596 16388 18602 16400
rect 18725 16397 18737 16400
rect 18771 16428 18783 16431
rect 19016 16428 19044 16468
rect 22405 16465 22417 16499
rect 22451 16496 22463 16499
rect 23322 16496 23328 16508
rect 22451 16468 23328 16496
rect 22451 16465 22463 16468
rect 22405 16459 22463 16465
rect 23322 16456 23328 16468
rect 23380 16496 23386 16508
rect 23380 16468 23644 16496
rect 23380 16456 23386 16468
rect 18771 16400 19044 16428
rect 19093 16431 19151 16437
rect 18771 16397 18783 16400
rect 18725 16391 18783 16397
rect 19093 16397 19105 16431
rect 19139 16428 19151 16431
rect 19274 16428 19280 16440
rect 19139 16400 19280 16428
rect 19139 16397 19151 16400
rect 19093 16391 19151 16397
rect 6857 16363 6915 16369
rect 6857 16360 6869 16363
rect 5768 16332 6869 16360
rect 5768 16304 5796 16332
rect 6857 16329 6869 16332
rect 6903 16329 6915 16363
rect 6857 16323 6915 16329
rect 8329 16363 8387 16369
rect 8329 16329 8341 16363
rect 8375 16329 8387 16363
rect 8329 16323 8387 16329
rect 8697 16363 8755 16369
rect 8697 16329 8709 16363
rect 8743 16360 8755 16363
rect 8970 16360 8976 16372
rect 8743 16332 8976 16360
rect 8743 16329 8755 16332
rect 8697 16323 8755 16329
rect 1242 16252 1248 16304
rect 1300 16292 1306 16304
rect 1521 16295 1579 16301
rect 1521 16292 1533 16295
rect 1300 16264 1533 16292
rect 1300 16252 1306 16264
rect 1521 16261 1533 16264
rect 1567 16261 1579 16295
rect 1521 16255 1579 16261
rect 1610 16252 1616 16304
rect 1668 16292 1674 16304
rect 1889 16295 1947 16301
rect 1889 16292 1901 16295
rect 1668 16264 1901 16292
rect 1668 16252 1674 16264
rect 1889 16261 1901 16264
rect 1935 16292 1947 16295
rect 1981 16295 2039 16301
rect 1981 16292 1993 16295
rect 1935 16264 1993 16292
rect 1935 16261 1947 16264
rect 1889 16255 1947 16261
rect 1981 16261 1993 16264
rect 2027 16261 2039 16295
rect 2990 16292 2996 16304
rect 2951 16264 2996 16292
rect 1981 16255 2039 16261
rect 2990 16252 2996 16264
rect 3048 16252 3054 16304
rect 5750 16292 5756 16304
rect 5711 16264 5756 16292
rect 5750 16252 5756 16264
rect 5808 16252 5814 16304
rect 7222 16292 7228 16304
rect 7183 16264 7228 16292
rect 7222 16252 7228 16264
rect 7280 16252 7286 16304
rect 8234 16292 8240 16304
rect 8195 16264 8240 16292
rect 8234 16252 8240 16264
rect 8292 16292 8298 16304
rect 8344 16292 8372 16323
rect 8970 16320 8976 16332
rect 9028 16360 9034 16372
rect 9338 16360 9344 16372
rect 9028 16332 9344 16360
rect 9028 16320 9034 16332
rect 9338 16320 9344 16332
rect 9396 16320 9402 16372
rect 11730 16320 11736 16372
rect 11788 16360 11794 16372
rect 11917 16363 11975 16369
rect 11917 16360 11929 16363
rect 11788 16332 11929 16360
rect 11788 16320 11794 16332
rect 11917 16329 11929 16332
rect 11963 16360 11975 16363
rect 12098 16360 12104 16372
rect 11963 16332 12104 16360
rect 11963 16329 11975 16332
rect 11917 16323 11975 16329
rect 12098 16320 12104 16332
rect 12156 16320 12162 16372
rect 15318 16320 15324 16372
rect 15376 16360 15382 16372
rect 15505 16363 15563 16369
rect 15505 16360 15517 16363
rect 15376 16332 15517 16360
rect 15376 16320 15382 16332
rect 15505 16329 15517 16332
rect 15551 16329 15563 16363
rect 15505 16323 15563 16329
rect 17437 16363 17495 16369
rect 17437 16329 17449 16363
rect 17483 16360 17495 16363
rect 19108 16360 19136 16391
rect 19274 16388 19280 16400
rect 19332 16388 19338 16440
rect 21209 16431 21267 16437
rect 21209 16397 21221 16431
rect 21255 16428 21267 16431
rect 21255 16400 21528 16428
rect 21255 16397 21267 16400
rect 21209 16391 21267 16397
rect 17483 16332 19136 16360
rect 17483 16329 17495 16332
rect 17437 16323 17495 16329
rect 21500 16304 21528 16400
rect 23230 16388 23236 16440
rect 23288 16428 23294 16440
rect 23616 16437 23644 16468
rect 23782 16456 23788 16508
rect 23840 16496 23846 16508
rect 24978 16496 24984 16508
rect 23840 16468 24984 16496
rect 23840 16456 23846 16468
rect 24978 16456 24984 16468
rect 25036 16456 25042 16508
rect 25717 16499 25775 16505
rect 25717 16465 25729 16499
rect 25763 16496 25775 16499
rect 25806 16496 25812 16508
rect 25763 16468 25812 16496
rect 25763 16465 25775 16468
rect 25717 16459 25775 16465
rect 25806 16456 25812 16468
rect 25864 16456 25870 16508
rect 25916 16505 25944 16536
rect 26358 16524 26364 16536
rect 26416 16524 26422 16576
rect 25901 16499 25959 16505
rect 25901 16465 25913 16499
rect 25947 16465 25959 16499
rect 25901 16459 25959 16465
rect 23417 16431 23475 16437
rect 23417 16428 23429 16431
rect 23288 16400 23429 16428
rect 23288 16388 23294 16400
rect 23417 16397 23429 16400
rect 23463 16397 23475 16431
rect 23417 16391 23475 16397
rect 23601 16431 23659 16437
rect 23601 16397 23613 16431
rect 23647 16397 23659 16431
rect 23601 16391 23659 16397
rect 23969 16431 24027 16437
rect 23969 16397 23981 16431
rect 24015 16397 24027 16431
rect 23969 16391 24027 16397
rect 22589 16363 22647 16369
rect 22589 16329 22601 16363
rect 22635 16360 22647 16363
rect 23690 16360 23696 16372
rect 22635 16332 23696 16360
rect 22635 16329 22647 16332
rect 22589 16323 22647 16329
rect 23690 16320 23696 16332
rect 23748 16360 23754 16372
rect 23984 16360 24012 16391
rect 24058 16388 24064 16440
rect 24116 16428 24122 16440
rect 24242 16428 24248 16440
rect 24116 16400 24248 16428
rect 24116 16388 24122 16400
rect 24242 16388 24248 16400
rect 24300 16388 24306 16440
rect 25625 16431 25683 16437
rect 25625 16397 25637 16431
rect 25671 16397 25683 16431
rect 25625 16391 25683 16397
rect 25993 16431 26051 16437
rect 25993 16397 26005 16431
rect 26039 16397 26051 16431
rect 25993 16391 26051 16397
rect 24521 16363 24579 16369
rect 23748 16332 24380 16360
rect 23748 16320 23754 16332
rect 8292 16264 8372 16292
rect 8292 16252 8298 16264
rect 8602 16252 8608 16304
rect 8660 16292 8666 16304
rect 8660 16264 8705 16292
rect 8660 16252 8666 16264
rect 10258 16252 10264 16304
rect 10316 16292 10322 16304
rect 10629 16295 10687 16301
rect 10629 16292 10641 16295
rect 10316 16264 10641 16292
rect 10316 16252 10322 16264
rect 10629 16261 10641 16264
rect 10675 16261 10687 16295
rect 10902 16292 10908 16304
rect 10863 16264 10908 16292
rect 10629 16255 10687 16261
rect 10902 16252 10908 16264
rect 10960 16252 10966 16304
rect 11178 16292 11184 16304
rect 11139 16264 11184 16292
rect 11178 16252 11184 16264
rect 11236 16252 11242 16304
rect 11454 16292 11460 16304
rect 11415 16264 11460 16292
rect 11454 16252 11460 16264
rect 11512 16252 11518 16304
rect 16698 16292 16704 16304
rect 16659 16264 16704 16292
rect 16698 16252 16704 16264
rect 16756 16252 16762 16304
rect 19366 16252 19372 16304
rect 19424 16292 19430 16304
rect 20013 16295 20071 16301
rect 20013 16292 20025 16295
rect 19424 16264 20025 16292
rect 19424 16252 19430 16264
rect 20013 16261 20025 16264
rect 20059 16292 20071 16295
rect 20286 16292 20292 16304
rect 20059 16264 20292 16292
rect 20059 16261 20071 16264
rect 20013 16255 20071 16261
rect 20286 16252 20292 16264
rect 20344 16252 20350 16304
rect 21482 16292 21488 16304
rect 21443 16264 21488 16292
rect 21482 16252 21488 16264
rect 21540 16252 21546 16304
rect 24352 16292 24380 16332
rect 24521 16329 24533 16363
rect 24567 16360 24579 16363
rect 25640 16360 25668 16391
rect 25806 16360 25812 16372
rect 24567 16332 25812 16360
rect 24567 16329 24579 16332
rect 24521 16323 24579 16329
rect 25806 16320 25812 16332
rect 25864 16320 25870 16372
rect 26008 16360 26036 16391
rect 26266 16360 26272 16372
rect 26008 16332 26272 16360
rect 26266 16320 26272 16332
rect 26324 16320 26330 16372
rect 24702 16292 24708 16304
rect 24352 16264 24708 16292
rect 24702 16252 24708 16264
rect 24760 16252 24766 16304
rect 400 16202 27264 16224
rect 400 16150 18870 16202
rect 18922 16150 18934 16202
rect 18986 16150 18998 16202
rect 19050 16150 19062 16202
rect 19114 16150 19126 16202
rect 19178 16150 27264 16202
rect 400 16128 27264 16150
rect 1702 16088 1708 16100
rect 1663 16060 1708 16088
rect 1702 16048 1708 16060
rect 1760 16048 1766 16100
rect 4097 16091 4155 16097
rect 4097 16057 4109 16091
rect 4143 16088 4155 16091
rect 4278 16088 4284 16100
rect 4143 16060 4284 16088
rect 4143 16057 4155 16060
rect 4097 16051 4155 16057
rect 4278 16048 4284 16060
rect 4336 16088 4342 16100
rect 8421 16091 8479 16097
rect 4336 16060 6624 16088
rect 4336 16048 4342 16060
rect 6596 16032 6624 16060
rect 8421 16057 8433 16091
rect 8467 16088 8479 16091
rect 9062 16088 9068 16100
rect 8467 16060 9068 16088
rect 8467 16057 8479 16060
rect 8421 16051 8479 16057
rect 9062 16048 9068 16060
rect 9120 16048 9126 16100
rect 9338 16048 9344 16100
rect 9396 16088 9402 16100
rect 9433 16091 9491 16097
rect 9433 16088 9445 16091
rect 9396 16060 9445 16088
rect 9396 16048 9402 16060
rect 9433 16057 9445 16060
rect 9479 16057 9491 16091
rect 12098 16088 12104 16100
rect 12059 16060 12104 16088
rect 9433 16051 9491 16057
rect 12098 16048 12104 16060
rect 12156 16048 12162 16100
rect 15873 16091 15931 16097
rect 15873 16057 15885 16091
rect 15919 16088 15931 16091
rect 16422 16088 16428 16100
rect 15919 16060 16428 16088
rect 15919 16057 15931 16060
rect 15873 16051 15931 16057
rect 16422 16048 16428 16060
rect 16480 16048 16486 16100
rect 17894 16048 17900 16100
rect 17952 16088 17958 16100
rect 25073 16091 25131 16097
rect 17952 16060 22724 16088
rect 17952 16048 17958 16060
rect 1794 15980 1800 16032
rect 1852 16020 1858 16032
rect 1852 15992 2116 16020
rect 1852 15980 1858 15992
rect 2088 15961 2116 15992
rect 5474 15980 5480 16032
rect 5532 16020 5538 16032
rect 6029 16023 6087 16029
rect 6029 16020 6041 16023
rect 5532 15992 6041 16020
rect 5532 15980 5538 15992
rect 6029 15989 6041 15992
rect 6075 15989 6087 16023
rect 6210 16020 6216 16032
rect 6171 15992 6216 16020
rect 6029 15983 6087 15989
rect 6210 15980 6216 15992
rect 6268 15980 6274 16032
rect 6578 16020 6584 16032
rect 6539 15992 6584 16020
rect 6578 15980 6584 15992
rect 6636 15980 6642 16032
rect 9522 16020 9528 16032
rect 8620 15992 9528 16020
rect 8620 15964 8648 15992
rect 9522 15980 9528 15992
rect 9580 15980 9586 16032
rect 11454 15980 11460 16032
rect 11512 16020 11518 16032
rect 11825 16023 11883 16029
rect 11825 16020 11837 16023
rect 11512 15992 11837 16020
rect 11512 15980 11518 15992
rect 11825 15989 11837 15992
rect 11871 16020 11883 16023
rect 12190 16020 12196 16032
rect 11871 15992 12196 16020
rect 11871 15989 11883 15992
rect 11825 15983 11883 15989
rect 12190 15980 12196 15992
rect 12248 16020 12254 16032
rect 13110 16020 13116 16032
rect 12248 15992 13116 16020
rect 12248 15980 12254 15992
rect 13110 15980 13116 15992
rect 13168 15980 13174 16032
rect 20654 15980 20660 16032
rect 20712 16020 20718 16032
rect 20712 15992 21252 16020
rect 20712 15980 20718 15992
rect 1889 15955 1947 15961
rect 1889 15921 1901 15955
rect 1935 15921 1947 15955
rect 1889 15915 1947 15921
rect 2073 15955 2131 15961
rect 2073 15921 2085 15955
rect 2119 15921 2131 15955
rect 2073 15915 2131 15921
rect 1794 15844 1800 15896
rect 1852 15884 1858 15896
rect 1904 15884 1932 15915
rect 5934 15912 5940 15964
rect 5992 15952 5998 15964
rect 6121 15955 6179 15961
rect 6121 15952 6133 15955
rect 5992 15924 6133 15952
rect 5992 15912 5998 15924
rect 6121 15921 6133 15924
rect 6167 15952 6179 15955
rect 8602 15952 8608 15964
rect 6167 15924 8608 15952
rect 6167 15921 6179 15924
rect 6121 15915 6179 15921
rect 8602 15912 8608 15924
rect 8660 15912 8666 15964
rect 9341 15955 9399 15961
rect 9341 15921 9353 15955
rect 9387 15952 9399 15955
rect 9706 15952 9712 15964
rect 9387 15924 9712 15952
rect 9387 15921 9399 15924
rect 9341 15915 9399 15921
rect 9706 15912 9712 15924
rect 9764 15912 9770 15964
rect 11362 15952 11368 15964
rect 11323 15924 11368 15952
rect 11362 15912 11368 15924
rect 11420 15912 11426 15964
rect 16606 15952 16612 15964
rect 16567 15924 16612 15952
rect 16606 15912 16612 15924
rect 16664 15912 16670 15964
rect 16974 15952 16980 15964
rect 16935 15924 16980 15952
rect 16974 15912 16980 15924
rect 17032 15912 17038 15964
rect 17066 15912 17072 15964
rect 17124 15952 17130 15964
rect 17161 15955 17219 15961
rect 17161 15952 17173 15955
rect 17124 15924 17173 15952
rect 17124 15912 17130 15924
rect 17161 15921 17173 15924
rect 17207 15952 17219 15955
rect 17802 15952 17808 15964
rect 17207 15924 17808 15952
rect 17207 15921 17219 15924
rect 17161 15915 17219 15921
rect 17802 15912 17808 15924
rect 17860 15912 17866 15964
rect 21022 15952 21028 15964
rect 20983 15924 21028 15952
rect 21022 15912 21028 15924
rect 21080 15912 21086 15964
rect 21224 15961 21252 15992
rect 22696 15964 22724 16060
rect 25073 16057 25085 16091
rect 25119 16088 25131 16091
rect 25714 16088 25720 16100
rect 25119 16060 25720 16088
rect 25119 16057 25131 16060
rect 25073 16051 25131 16057
rect 25714 16048 25720 16060
rect 25772 16048 25778 16100
rect 23414 15980 23420 16032
rect 23472 16020 23478 16032
rect 23472 15992 24564 16020
rect 23472 15980 23478 15992
rect 21209 15955 21267 15961
rect 21209 15921 21221 15955
rect 21255 15921 21267 15955
rect 21209 15915 21267 15921
rect 22678 15912 22684 15964
rect 22736 15952 22742 15964
rect 24536 15961 24564 15992
rect 23877 15955 23935 15961
rect 23877 15952 23889 15955
rect 22736 15924 23889 15952
rect 22736 15912 22742 15924
rect 23877 15921 23889 15924
rect 23923 15921 23935 15955
rect 23877 15915 23935 15921
rect 24521 15955 24579 15961
rect 24521 15921 24533 15955
rect 24567 15921 24579 15955
rect 25806 15952 25812 15964
rect 25767 15924 25812 15952
rect 24521 15915 24579 15921
rect 25806 15912 25812 15924
rect 25864 15912 25870 15964
rect 4922 15884 4928 15896
rect 1852 15856 4928 15884
rect 1852 15844 1858 15856
rect 4922 15844 4928 15856
rect 4980 15844 4986 15896
rect 5842 15884 5848 15896
rect 5803 15856 5848 15884
rect 5842 15844 5848 15856
rect 5900 15844 5906 15896
rect 6670 15844 6676 15896
rect 6728 15884 6734 15896
rect 8234 15884 8240 15896
rect 6728 15856 8240 15884
rect 6728 15844 6734 15856
rect 8234 15844 8240 15856
rect 8292 15884 8298 15896
rect 9154 15884 9160 15896
rect 8292 15856 9160 15884
rect 8292 15844 8298 15856
rect 9154 15844 9160 15856
rect 9212 15844 9218 15896
rect 9798 15844 9804 15896
rect 9856 15884 9862 15896
rect 9893 15887 9951 15893
rect 9893 15884 9905 15887
rect 9856 15856 9905 15884
rect 9856 15844 9862 15856
rect 9893 15853 9905 15856
rect 9939 15884 9951 15887
rect 9982 15884 9988 15896
rect 9939 15856 9988 15884
rect 9939 15853 9951 15856
rect 9893 15847 9951 15853
rect 9982 15844 9988 15856
rect 10040 15844 10046 15896
rect 13113 15887 13171 15893
rect 13113 15853 13125 15887
rect 13159 15884 13171 15887
rect 13386 15884 13392 15896
rect 13159 15856 13392 15884
rect 13159 15853 13171 15856
rect 13113 15847 13171 15853
rect 13386 15844 13392 15856
rect 13444 15844 13450 15896
rect 13662 15884 13668 15896
rect 13623 15856 13668 15884
rect 13662 15844 13668 15856
rect 13720 15884 13726 15896
rect 14674 15884 14680 15896
rect 13720 15856 14680 15884
rect 13720 15844 13726 15856
rect 14674 15844 14680 15856
rect 14732 15844 14738 15896
rect 15226 15844 15232 15896
rect 15284 15884 15290 15896
rect 16517 15887 16575 15893
rect 16517 15884 16529 15887
rect 15284 15856 16529 15884
rect 15284 15844 15290 15856
rect 16517 15853 16529 15856
rect 16563 15884 16575 15887
rect 16698 15884 16704 15896
rect 16563 15856 16704 15884
rect 16563 15853 16575 15856
rect 16517 15847 16575 15853
rect 16698 15844 16704 15856
rect 16756 15844 16762 15896
rect 20194 15884 20200 15896
rect 20155 15856 20200 15884
rect 20194 15844 20200 15856
rect 20252 15844 20258 15896
rect 20749 15887 20807 15893
rect 20749 15853 20761 15887
rect 20795 15853 20807 15887
rect 20749 15847 20807 15853
rect 24153 15887 24211 15893
rect 24153 15853 24165 15887
rect 24199 15884 24211 15887
rect 24242 15884 24248 15896
rect 24199 15856 24248 15884
rect 24199 15853 24211 15856
rect 24153 15847 24211 15853
rect 2070 15776 2076 15828
rect 2128 15816 2134 15828
rect 2533 15819 2591 15825
rect 2533 15816 2545 15819
rect 2128 15788 2545 15816
rect 2128 15776 2134 15788
rect 2533 15785 2545 15788
rect 2579 15816 2591 15819
rect 2990 15816 2996 15828
rect 2579 15788 2996 15816
rect 2579 15785 2591 15788
rect 2533 15779 2591 15785
rect 2990 15776 2996 15788
rect 3048 15776 3054 15828
rect 9614 15776 9620 15828
rect 9672 15816 9678 15828
rect 11822 15816 11828 15828
rect 9672 15788 11828 15816
rect 9672 15776 9678 15788
rect 11822 15776 11828 15788
rect 11880 15816 11886 15828
rect 11917 15819 11975 15825
rect 11917 15816 11929 15819
rect 11880 15788 11929 15816
rect 11880 15776 11886 15788
rect 11917 15785 11929 15788
rect 11963 15785 11975 15819
rect 13570 15816 13576 15828
rect 13531 15788 13576 15816
rect 11917 15779 11975 15785
rect 13570 15776 13576 15788
rect 13628 15776 13634 15828
rect 20286 15776 20292 15828
rect 20344 15816 20350 15828
rect 20764 15816 20792 15847
rect 24242 15844 24248 15856
rect 24300 15844 24306 15896
rect 24702 15844 24708 15896
rect 24760 15884 24766 15896
rect 24797 15887 24855 15893
rect 24797 15884 24809 15887
rect 24760 15856 24809 15884
rect 24760 15844 24766 15856
rect 24797 15853 24809 15856
rect 24843 15884 24855 15887
rect 24843 15856 26128 15884
rect 24843 15853 24855 15856
rect 24797 15847 24855 15853
rect 21482 15816 21488 15828
rect 20344 15788 21488 15816
rect 20344 15776 20350 15788
rect 21482 15776 21488 15788
rect 21540 15776 21546 15828
rect 24058 15816 24064 15828
rect 24019 15788 24064 15816
rect 24058 15776 24064 15788
rect 24116 15776 24122 15828
rect 2162 15748 2168 15760
rect 2123 15720 2168 15748
rect 2162 15708 2168 15720
rect 2220 15708 2226 15760
rect 6302 15708 6308 15760
rect 6360 15748 6366 15760
rect 6673 15751 6731 15757
rect 6673 15748 6685 15751
rect 6360 15720 6685 15748
rect 6360 15708 6366 15720
rect 6673 15717 6685 15720
rect 6719 15717 6731 15751
rect 7774 15748 7780 15760
rect 7735 15720 7780 15748
rect 6673 15711 6731 15717
rect 7774 15708 7780 15720
rect 7832 15708 7838 15760
rect 11546 15748 11552 15760
rect 11507 15720 11552 15748
rect 11546 15708 11552 15720
rect 11604 15708 11610 15760
rect 15318 15748 15324 15760
rect 15279 15720 15324 15748
rect 15318 15708 15324 15720
rect 15376 15708 15382 15760
rect 16057 15751 16115 15757
rect 16057 15717 16069 15751
rect 16103 15748 16115 15751
rect 16882 15748 16888 15760
rect 16103 15720 16888 15748
rect 16103 15717 16115 15720
rect 16057 15711 16115 15717
rect 16882 15708 16888 15720
rect 16940 15708 16946 15760
rect 23049 15751 23107 15757
rect 23049 15717 23061 15751
rect 23095 15748 23107 15751
rect 23230 15748 23236 15760
rect 23095 15720 23236 15748
rect 23095 15717 23107 15720
rect 23049 15711 23107 15717
rect 23230 15708 23236 15720
rect 23288 15708 23294 15760
rect 26100 15757 26128 15856
rect 26085 15751 26143 15757
rect 26085 15717 26097 15751
rect 26131 15748 26143 15751
rect 26266 15748 26272 15760
rect 26131 15720 26272 15748
rect 26131 15717 26143 15720
rect 26085 15711 26143 15717
rect 26266 15708 26272 15720
rect 26324 15708 26330 15760
rect 400 15658 27264 15680
rect 400 15606 3510 15658
rect 3562 15606 3574 15658
rect 3626 15606 3638 15658
rect 3690 15606 3702 15658
rect 3754 15606 3766 15658
rect 3818 15606 27264 15658
rect 400 15584 27264 15606
rect 1794 15544 1800 15556
rect 1755 15516 1800 15544
rect 1794 15504 1800 15516
rect 1852 15504 1858 15556
rect 1886 15504 1892 15556
rect 1944 15544 1950 15556
rect 2349 15547 2407 15553
rect 1944 15516 1989 15544
rect 1944 15504 1950 15516
rect 2349 15513 2361 15547
rect 2395 15544 2407 15547
rect 2438 15544 2444 15556
rect 2395 15516 2444 15544
rect 2395 15513 2407 15516
rect 2349 15507 2407 15513
rect 2438 15504 2444 15516
rect 2496 15504 2502 15556
rect 2990 15544 2996 15556
rect 2903 15516 2996 15544
rect 2990 15504 2996 15516
rect 3048 15544 3054 15556
rect 3910 15544 3916 15556
rect 3048 15516 3916 15544
rect 3048 15504 3054 15516
rect 3910 15504 3916 15516
rect 3968 15504 3974 15556
rect 4002 15504 4008 15556
rect 4060 15544 4066 15556
rect 4373 15547 4431 15553
rect 4373 15544 4385 15547
rect 4060 15516 4385 15544
rect 4060 15504 4066 15516
rect 4373 15513 4385 15516
rect 4419 15544 4431 15547
rect 4925 15547 4983 15553
rect 4925 15544 4937 15547
rect 4419 15516 4937 15544
rect 4419 15513 4431 15516
rect 4373 15507 4431 15513
rect 4925 15513 4937 15516
rect 4971 15513 4983 15547
rect 4925 15507 4983 15513
rect 7225 15547 7283 15553
rect 7225 15513 7237 15547
rect 7271 15544 7283 15547
rect 8145 15547 8203 15553
rect 8145 15544 8157 15547
rect 7271 15516 8157 15544
rect 7271 15513 7283 15516
rect 7225 15507 7283 15513
rect 8145 15513 8157 15516
rect 8191 15544 8203 15547
rect 9614 15544 9620 15556
rect 8191 15516 9620 15544
rect 8191 15513 8203 15516
rect 8145 15507 8203 15513
rect 1702 15436 1708 15488
rect 1760 15476 1766 15488
rect 2533 15479 2591 15485
rect 2533 15476 2545 15479
rect 1760 15448 2545 15476
rect 1760 15436 1766 15448
rect 2533 15445 2545 15448
rect 2579 15476 2591 15479
rect 3085 15479 3143 15485
rect 3085 15476 3097 15479
rect 2579 15448 3097 15476
rect 2579 15445 2591 15448
rect 2533 15439 2591 15445
rect 3085 15445 3097 15448
rect 3131 15445 3143 15479
rect 4940 15476 4968 15507
rect 9614 15504 9620 15516
rect 9672 15504 9678 15556
rect 9798 15544 9804 15556
rect 9759 15516 9804 15544
rect 9798 15504 9804 15516
rect 9856 15504 9862 15556
rect 11362 15544 11368 15556
rect 11323 15516 11368 15544
rect 11362 15504 11368 15516
rect 11420 15504 11426 15556
rect 11546 15544 11552 15556
rect 11507 15516 11552 15544
rect 11546 15504 11552 15516
rect 11604 15504 11610 15556
rect 15226 15544 15232 15556
rect 15187 15516 15232 15544
rect 15226 15504 15232 15516
rect 15284 15504 15290 15556
rect 15410 15504 15416 15556
rect 15468 15544 15474 15556
rect 15870 15544 15876 15556
rect 15468 15516 15876 15544
rect 15468 15504 15474 15516
rect 15870 15504 15876 15516
rect 15928 15544 15934 15556
rect 16149 15547 16207 15553
rect 16149 15544 16161 15547
rect 15928 15516 16161 15544
rect 15928 15504 15934 15516
rect 16149 15513 16161 15516
rect 16195 15513 16207 15547
rect 16882 15544 16888 15556
rect 16843 15516 16888 15544
rect 16149 15507 16207 15513
rect 16882 15504 16888 15516
rect 16940 15504 16946 15556
rect 20286 15544 20292 15556
rect 20247 15516 20292 15544
rect 20286 15504 20292 15516
rect 20344 15504 20350 15556
rect 20657 15547 20715 15553
rect 20657 15513 20669 15547
rect 20703 15544 20715 15547
rect 21022 15544 21028 15556
rect 20703 15516 21028 15544
rect 20703 15513 20715 15516
rect 20657 15507 20715 15513
rect 21022 15504 21028 15516
rect 21080 15504 21086 15556
rect 24058 15544 24064 15556
rect 24019 15516 24064 15544
rect 24058 15504 24064 15516
rect 24116 15504 24122 15556
rect 26266 15544 26272 15556
rect 26227 15516 26272 15544
rect 26266 15504 26272 15516
rect 26324 15504 26330 15556
rect 6946 15476 6952 15488
rect 4940 15448 6952 15476
rect 3085 15439 3143 15445
rect 6946 15436 6952 15448
rect 7004 15436 7010 15488
rect 7774 15436 7780 15488
rect 7832 15485 7838 15488
rect 7832 15479 7881 15485
rect 7832 15445 7835 15479
rect 7869 15445 7881 15479
rect 7832 15439 7881 15445
rect 7832 15436 7838 15439
rect 7958 15436 7964 15488
rect 8016 15476 8022 15488
rect 9249 15479 9307 15485
rect 8016 15448 8109 15476
rect 8016 15436 8022 15448
rect 9249 15445 9261 15479
rect 9295 15476 9307 15479
rect 9338 15476 9344 15488
rect 9295 15448 9344 15476
rect 9295 15445 9307 15448
rect 9249 15439 9307 15445
rect 1886 15368 1892 15420
rect 1944 15408 1950 15420
rect 2220 15411 2278 15417
rect 2220 15408 2232 15411
rect 1944 15380 2232 15408
rect 1944 15368 1950 15380
rect 2220 15377 2232 15380
rect 2266 15377 2278 15411
rect 2220 15371 2278 15377
rect 2441 15411 2499 15417
rect 2441 15377 2453 15411
rect 2487 15408 2499 15411
rect 2622 15408 2628 15420
rect 2487 15380 2628 15408
rect 2487 15377 2499 15380
rect 2441 15371 2499 15377
rect 2622 15368 2628 15380
rect 2680 15408 2686 15420
rect 3266 15408 3272 15420
rect 2680 15380 3272 15408
rect 2680 15368 2686 15380
rect 3266 15368 3272 15380
rect 3324 15368 3330 15420
rect 4557 15411 4615 15417
rect 4557 15377 4569 15411
rect 4603 15408 4615 15411
rect 5566 15408 5572 15420
rect 4603 15380 5572 15408
rect 4603 15377 4615 15380
rect 4557 15371 4615 15377
rect 874 15340 880 15352
rect 835 15312 880 15340
rect 874 15300 880 15312
rect 932 15340 938 15352
rect 1337 15343 1395 15349
rect 1337 15340 1349 15343
rect 932 15312 1349 15340
rect 932 15300 938 15312
rect 1337 15309 1349 15312
rect 1383 15309 1395 15343
rect 1337 15303 1395 15309
rect 1978 15300 1984 15352
rect 2036 15340 2042 15352
rect 4756 15349 4784 15380
rect 5566 15368 5572 15380
rect 5624 15368 5630 15420
rect 5753 15411 5811 15417
rect 5753 15377 5765 15411
rect 5799 15408 5811 15411
rect 5842 15408 5848 15420
rect 5799 15380 5848 15408
rect 5799 15377 5811 15380
rect 5753 15371 5811 15377
rect 5842 15368 5848 15380
rect 5900 15408 5906 15420
rect 5937 15411 5995 15417
rect 5937 15408 5949 15411
rect 5900 15380 5949 15408
rect 5900 15368 5906 15380
rect 5937 15377 5949 15380
rect 5983 15408 5995 15411
rect 6121 15411 6179 15417
rect 6121 15408 6133 15411
rect 5983 15380 6133 15408
rect 5983 15377 5995 15380
rect 5937 15371 5995 15377
rect 6121 15377 6133 15380
rect 6167 15408 6179 15411
rect 6670 15408 6676 15420
rect 6167 15380 6676 15408
rect 6167 15377 6179 15380
rect 6121 15371 6179 15377
rect 6670 15368 6676 15380
rect 6728 15368 6734 15420
rect 6854 15408 6860 15420
rect 6815 15380 6860 15408
rect 6854 15368 6860 15380
rect 6912 15368 6918 15420
rect 7130 15368 7136 15420
rect 7188 15408 7194 15420
rect 7501 15411 7559 15417
rect 7501 15408 7513 15411
rect 7188 15380 7513 15408
rect 7188 15368 7194 15380
rect 7501 15377 7513 15380
rect 7547 15408 7559 15411
rect 7976 15408 8004 15436
rect 7547 15380 8004 15408
rect 7547 15377 7559 15380
rect 7501 15371 7559 15377
rect 8050 15368 8056 15420
rect 8108 15408 8114 15420
rect 8513 15411 8571 15417
rect 8513 15408 8525 15411
rect 8108 15380 8525 15408
rect 8108 15368 8114 15380
rect 8513 15377 8525 15380
rect 8559 15377 8571 15411
rect 8513 15371 8571 15377
rect 2073 15343 2131 15349
rect 2073 15340 2085 15343
rect 2036 15312 2085 15340
rect 2036 15300 2042 15312
rect 2073 15309 2085 15312
rect 2119 15309 2131 15343
rect 2073 15303 2131 15309
rect 4649 15343 4707 15349
rect 4649 15309 4661 15343
rect 4695 15309 4707 15343
rect 4649 15303 4707 15309
rect 4741 15343 4799 15349
rect 4741 15309 4753 15343
rect 4787 15309 4799 15343
rect 4741 15303 4799 15309
rect 1245 15275 1303 15281
rect 1245 15241 1257 15275
rect 1291 15272 1303 15275
rect 1613 15275 1671 15281
rect 1613 15272 1625 15275
rect 1291 15244 1625 15272
rect 1291 15241 1303 15244
rect 1245 15235 1303 15241
rect 1613 15241 1625 15244
rect 1659 15272 1671 15275
rect 1702 15272 1708 15284
rect 1659 15244 1708 15272
rect 1659 15241 1671 15244
rect 1613 15235 1671 15241
rect 1702 15232 1708 15244
rect 1760 15232 1766 15284
rect 4664 15272 4692 15303
rect 5106 15300 5112 15352
rect 5164 15340 5170 15352
rect 5385 15343 5443 15349
rect 5385 15340 5397 15343
rect 5164 15312 5397 15340
rect 5164 15300 5170 15312
rect 5385 15309 5397 15312
rect 5431 15340 5443 15343
rect 6397 15343 6455 15349
rect 6397 15340 6409 15343
rect 5431 15312 6409 15340
rect 5431 15309 5443 15312
rect 5385 15303 5443 15309
rect 6397 15309 6409 15312
rect 6443 15340 6455 15343
rect 7041 15343 7099 15349
rect 7041 15340 7053 15343
rect 6443 15312 7053 15340
rect 6443 15309 6455 15312
rect 6397 15303 6455 15309
rect 7041 15309 7053 15312
rect 7087 15340 7099 15343
rect 9264 15340 9292 15439
rect 9338 15436 9344 15448
rect 9396 15436 9402 15488
rect 9522 15476 9528 15488
rect 9483 15448 9528 15476
rect 9522 15436 9528 15448
rect 9580 15436 9586 15488
rect 13570 15436 13576 15488
rect 13628 15476 13634 15488
rect 14401 15479 14459 15485
rect 14401 15476 14413 15479
rect 13628 15448 14413 15476
rect 13628 15436 13634 15448
rect 14401 15445 14413 15448
rect 14447 15445 14459 15479
rect 14401 15439 14459 15445
rect 15597 15479 15655 15485
rect 15597 15445 15609 15479
rect 15643 15476 15655 15479
rect 15778 15476 15784 15488
rect 15643 15448 15784 15476
rect 15643 15445 15655 15448
rect 15597 15439 15655 15445
rect 15778 15436 15784 15448
rect 15836 15476 15842 15488
rect 17066 15476 17072 15488
rect 15836 15448 17072 15476
rect 15836 15436 15842 15448
rect 17066 15436 17072 15448
rect 17124 15436 17130 15488
rect 20194 15436 20200 15488
rect 20252 15476 20258 15488
rect 20749 15479 20807 15485
rect 20749 15476 20761 15479
rect 20252 15448 20761 15476
rect 20252 15436 20258 15448
rect 20749 15445 20761 15448
rect 20795 15445 20807 15479
rect 20749 15439 20807 15445
rect 12469 15411 12527 15417
rect 12469 15377 12481 15411
rect 12515 15408 12527 15411
rect 14122 15408 14128 15420
rect 12515 15380 14128 15408
rect 12515 15377 12527 15380
rect 12469 15371 12527 15377
rect 7087 15312 9292 15340
rect 13113 15343 13171 15349
rect 7087 15309 7099 15312
rect 7041 15303 7099 15309
rect 13113 15309 13125 15343
rect 13159 15340 13171 15343
rect 13386 15340 13392 15352
rect 13159 15312 13392 15340
rect 13159 15309 13171 15312
rect 13113 15303 13171 15309
rect 13386 15300 13392 15312
rect 13444 15300 13450 15352
rect 14048 15349 14076 15380
rect 14122 15368 14128 15380
rect 14180 15368 14186 15420
rect 15318 15368 15324 15420
rect 15376 15408 15382 15420
rect 15413 15411 15471 15417
rect 15413 15408 15425 15411
rect 15376 15380 15425 15408
rect 15376 15368 15382 15380
rect 15413 15377 15425 15380
rect 15459 15408 15471 15411
rect 16606 15408 16612 15420
rect 15459 15380 16612 15408
rect 15459 15377 15471 15380
rect 15413 15371 15471 15377
rect 16606 15368 16612 15380
rect 16664 15368 16670 15420
rect 20473 15411 20531 15417
rect 20473 15377 20485 15411
rect 20519 15408 20531 15411
rect 20654 15408 20660 15420
rect 20519 15380 20660 15408
rect 20519 15377 20531 15380
rect 20473 15371 20531 15377
rect 20654 15368 20660 15380
rect 20712 15368 20718 15420
rect 23601 15411 23659 15417
rect 23601 15377 23613 15411
rect 23647 15408 23659 15411
rect 24076 15408 24104 15504
rect 24429 15411 24487 15417
rect 24429 15408 24441 15411
rect 23647 15380 24441 15408
rect 23647 15377 23659 15380
rect 23601 15371 23659 15377
rect 24429 15377 24441 15380
rect 24475 15377 24487 15411
rect 24429 15371 24487 15377
rect 25806 15368 25812 15420
rect 25864 15408 25870 15420
rect 26177 15411 26235 15417
rect 26177 15408 26189 15411
rect 25864 15380 26189 15408
rect 25864 15368 25870 15380
rect 26177 15377 26189 15380
rect 26223 15408 26235 15411
rect 26453 15411 26511 15417
rect 26453 15408 26465 15411
rect 26223 15380 26465 15408
rect 26223 15377 26235 15380
rect 26177 15371 26235 15377
rect 26453 15377 26465 15380
rect 26499 15377 26511 15411
rect 26453 15371 26511 15377
rect 14033 15343 14091 15349
rect 14033 15309 14045 15343
rect 14079 15309 14091 15343
rect 16057 15343 16115 15349
rect 16057 15340 16069 15343
rect 14033 15303 14091 15309
rect 14186 15312 16069 15340
rect 5124 15272 5152 15300
rect 4664 15244 5152 15272
rect 6481 15275 6539 15281
rect 6481 15241 6493 15275
rect 6527 15241 6539 15275
rect 7685 15275 7743 15281
rect 7685 15272 7697 15275
rect 6481 15235 6539 15241
rect 7332 15244 7697 15272
rect 5474 15204 5480 15216
rect 5435 15176 5480 15204
rect 5474 15164 5480 15176
rect 5532 15164 5538 15216
rect 6302 15204 6308 15216
rect 6263 15176 6308 15204
rect 6302 15164 6308 15176
rect 6360 15164 6366 15216
rect 6394 15164 6400 15216
rect 6452 15204 6458 15216
rect 6504 15204 6532 15235
rect 7332 15216 7360 15244
rect 7685 15241 7697 15244
rect 7731 15241 7743 15275
rect 7685 15235 7743 15241
rect 7866 15232 7872 15284
rect 7924 15272 7930 15284
rect 14186 15272 14214 15312
rect 16057 15309 16069 15312
rect 16103 15340 16115 15343
rect 16517 15343 16575 15349
rect 16517 15340 16529 15343
rect 16103 15312 16529 15340
rect 16103 15309 16115 15312
rect 16057 15303 16115 15309
rect 16517 15309 16529 15312
rect 16563 15340 16575 15343
rect 16701 15343 16759 15349
rect 16701 15340 16713 15343
rect 16563 15312 16713 15340
rect 16563 15309 16575 15312
rect 16517 15303 16575 15309
rect 16701 15309 16713 15312
rect 16747 15340 16759 15343
rect 16974 15340 16980 15352
rect 16747 15312 16980 15340
rect 16747 15309 16759 15312
rect 16701 15303 16759 15309
rect 16974 15300 16980 15312
rect 17032 15300 17038 15352
rect 22589 15343 22647 15349
rect 22589 15309 22601 15343
rect 22635 15340 22647 15343
rect 22770 15340 22776 15352
rect 22635 15312 22776 15340
rect 22635 15309 22647 15312
rect 22589 15303 22647 15309
rect 22770 15300 22776 15312
rect 22828 15340 22834 15352
rect 23233 15343 23291 15349
rect 23233 15340 23245 15343
rect 22828 15312 23245 15340
rect 22828 15300 22834 15312
rect 23233 15309 23245 15312
rect 23279 15340 23291 15343
rect 23782 15340 23788 15352
rect 23279 15312 23788 15340
rect 23279 15309 23291 15312
rect 23233 15303 23291 15309
rect 23782 15300 23788 15312
rect 23840 15300 23846 15352
rect 24153 15343 24211 15349
rect 24153 15309 24165 15343
rect 24199 15309 24211 15343
rect 24153 15303 24211 15309
rect 7924 15244 14214 15272
rect 7924 15232 7930 15244
rect 15778 15232 15784 15284
rect 15836 15272 15842 15284
rect 15873 15275 15931 15281
rect 15873 15272 15885 15275
rect 15836 15244 15885 15272
rect 15836 15232 15842 15244
rect 15873 15241 15885 15244
rect 15919 15241 15931 15275
rect 24168 15272 24196 15303
rect 24334 15272 24340 15284
rect 24168 15244 24340 15272
rect 15873 15235 15931 15241
rect 24334 15232 24340 15244
rect 24392 15232 24398 15284
rect 24886 15232 24892 15284
rect 24944 15232 24950 15284
rect 7314 15204 7320 15216
rect 6452 15176 6532 15204
rect 7275 15176 7320 15204
rect 6452 15164 6458 15176
rect 7314 15164 7320 15176
rect 7372 15164 7378 15216
rect 9154 15164 9160 15216
rect 9212 15204 9218 15216
rect 9341 15207 9399 15213
rect 9341 15204 9353 15207
rect 9212 15176 9353 15204
rect 9212 15164 9218 15176
rect 9341 15173 9353 15176
rect 9387 15173 9399 15207
rect 9341 15167 9399 15173
rect 9706 15164 9712 15216
rect 9764 15204 9770 15216
rect 9893 15207 9951 15213
rect 9893 15204 9905 15207
rect 9764 15176 9905 15204
rect 9764 15164 9770 15176
rect 9893 15173 9905 15176
rect 9939 15173 9951 15207
rect 12650 15204 12656 15216
rect 12611 15176 12656 15204
rect 9893 15167 9951 15173
rect 12650 15164 12656 15176
rect 12708 15164 12714 15216
rect 12837 15207 12895 15213
rect 12837 15173 12849 15207
rect 12883 15204 12895 15207
rect 13021 15207 13079 15213
rect 13021 15204 13033 15207
rect 12883 15176 13033 15204
rect 12883 15173 12895 15176
rect 12837 15167 12895 15173
rect 13021 15173 13033 15176
rect 13067 15204 13079 15207
rect 13386 15204 13392 15216
rect 13067 15176 13392 15204
rect 13067 15173 13079 15176
rect 13021 15167 13079 15173
rect 13386 15164 13392 15176
rect 13444 15164 13450 15216
rect 22678 15204 22684 15216
rect 22639 15176 22684 15204
rect 22678 15164 22684 15176
rect 22736 15164 22742 15216
rect 23230 15204 23236 15216
rect 23191 15176 23236 15204
rect 23230 15164 23236 15176
rect 23288 15164 23294 15216
rect 23785 15207 23843 15213
rect 23785 15173 23797 15207
rect 23831 15204 23843 15207
rect 24242 15204 24248 15216
rect 23831 15176 24248 15204
rect 23831 15173 23843 15176
rect 23785 15167 23843 15173
rect 24242 15164 24248 15176
rect 24300 15164 24306 15216
rect 400 15114 27264 15136
rect 400 15062 18870 15114
rect 18922 15062 18934 15114
rect 18986 15062 18998 15114
rect 19050 15062 19062 15114
rect 19114 15062 19126 15114
rect 19178 15062 27264 15114
rect 400 15040 27264 15062
rect 1978 15000 1984 15012
rect 1891 14972 1984 15000
rect 1978 14960 1984 14972
rect 2036 15000 2042 15012
rect 2162 15000 2168 15012
rect 2036 14972 2168 15000
rect 2036 14960 2042 14972
rect 2162 14960 2168 14972
rect 2220 14960 2226 15012
rect 4281 15003 4339 15009
rect 4281 14969 4293 15003
rect 4327 15000 4339 15003
rect 4554 15000 4560 15012
rect 4327 14972 4560 15000
rect 4327 14969 4339 14972
rect 4281 14963 4339 14969
rect 4554 14960 4560 14972
rect 4612 15000 4618 15012
rect 5382 15000 5388 15012
rect 4612 14972 5388 15000
rect 4612 14960 4618 14972
rect 5382 14960 5388 14972
rect 5440 14960 5446 15012
rect 5934 15000 5940 15012
rect 5895 14972 5940 15000
rect 5934 14960 5940 14972
rect 5992 14960 5998 15012
rect 6210 14960 6216 15012
rect 6268 15000 6274 15012
rect 6670 15000 6676 15012
rect 6268 14972 6676 15000
rect 6268 14960 6274 14972
rect 6670 14960 6676 14972
rect 6728 14960 6734 15012
rect 8694 14960 8700 15012
rect 8752 15000 8758 15012
rect 9614 15000 9620 15012
rect 8752 14972 9620 15000
rect 8752 14960 8758 14972
rect 9614 14960 9620 14972
rect 9672 14960 9678 15012
rect 12006 15000 12012 15012
rect 11967 14972 12012 15000
rect 12006 14960 12012 14972
rect 12064 15000 12070 15012
rect 12193 15003 12251 15009
rect 12193 15000 12205 15003
rect 12064 14972 12205 15000
rect 12064 14960 12070 14972
rect 12193 14969 12205 14972
rect 12239 14969 12251 15003
rect 12193 14963 12251 14969
rect 13205 15003 13263 15009
rect 13205 14969 13217 15003
rect 13251 15000 13263 15003
rect 13662 15000 13668 15012
rect 13251 14972 13668 15000
rect 13251 14969 13263 14972
rect 13205 14963 13263 14969
rect 13662 14960 13668 14972
rect 13720 14960 13726 15012
rect 15870 15000 15876 15012
rect 15831 14972 15876 15000
rect 15870 14960 15876 14972
rect 15928 14960 15934 15012
rect 23690 15000 23696 15012
rect 23651 14972 23696 15000
rect 23690 14960 23696 14972
rect 23748 14960 23754 15012
rect 24245 15003 24303 15009
rect 24245 14969 24257 15003
rect 24291 15000 24303 15003
rect 24886 15000 24892 15012
rect 24291 14972 24892 15000
rect 24291 14969 24303 14972
rect 24245 14963 24303 14969
rect 24886 14960 24892 14972
rect 24944 14960 24950 15012
rect 1886 14892 1892 14944
rect 1944 14932 1950 14944
rect 2441 14935 2499 14941
rect 2441 14932 2453 14935
rect 1944 14904 2453 14932
rect 1944 14892 1950 14904
rect 2441 14901 2453 14904
rect 2487 14932 2499 14935
rect 2530 14932 2536 14944
rect 2487 14904 2536 14932
rect 2487 14901 2499 14904
rect 2441 14895 2499 14901
rect 2530 14892 2536 14904
rect 2588 14892 2594 14944
rect 2714 14892 2720 14944
rect 2772 14932 2778 14944
rect 4097 14935 4155 14941
rect 4097 14932 4109 14935
rect 2772 14904 4109 14932
rect 2772 14892 2778 14904
rect 4097 14901 4109 14904
rect 4143 14932 4155 14935
rect 4370 14932 4376 14944
rect 4143 14904 4376 14932
rect 4143 14901 4155 14904
rect 4097 14895 4155 14901
rect 4370 14892 4376 14904
rect 4428 14892 4434 14944
rect 5106 14892 5112 14944
rect 5164 14932 5170 14944
rect 5477 14935 5535 14941
rect 5164 14904 5428 14932
rect 5164 14892 5170 14904
rect 2165 14867 2223 14873
rect 2165 14833 2177 14867
rect 2211 14864 2223 14867
rect 2622 14864 2628 14876
rect 2211 14836 2628 14864
rect 2211 14833 2223 14836
rect 2165 14827 2223 14833
rect 2622 14824 2628 14836
rect 2680 14864 2686 14876
rect 2806 14864 2812 14876
rect 2680 14836 2812 14864
rect 2680 14824 2686 14836
rect 2806 14824 2812 14836
rect 2864 14824 2870 14876
rect 3450 14864 3456 14876
rect 3411 14836 3456 14864
rect 3450 14824 3456 14836
rect 3508 14864 3514 14876
rect 5014 14864 5020 14876
rect 3508 14836 5020 14864
rect 3508 14824 3514 14836
rect 5014 14824 5020 14836
rect 5072 14824 5078 14876
rect 5290 14864 5296 14876
rect 5251 14836 5296 14864
rect 5290 14824 5296 14836
rect 5348 14824 5354 14876
rect 5400 14873 5428 14904
rect 5477 14901 5489 14935
rect 5523 14932 5535 14935
rect 5842 14932 5848 14944
rect 5523 14904 5848 14932
rect 5523 14901 5535 14904
rect 5477 14895 5535 14901
rect 5842 14892 5848 14904
rect 5900 14892 5906 14944
rect 6578 14932 6584 14944
rect 6539 14904 6584 14932
rect 6578 14892 6584 14904
rect 6636 14892 6642 14944
rect 12650 14892 12656 14944
rect 12708 14932 12714 14944
rect 13297 14935 13355 14941
rect 13297 14932 13309 14935
rect 12708 14904 13309 14932
rect 12708 14892 12714 14904
rect 13297 14901 13309 14904
rect 13343 14932 13355 14935
rect 13570 14932 13576 14944
rect 13343 14904 13576 14932
rect 13343 14901 13355 14904
rect 13297 14895 13355 14901
rect 13570 14892 13576 14904
rect 13628 14892 13634 14944
rect 16882 14892 16888 14944
rect 16940 14932 16946 14944
rect 16940 14904 18032 14932
rect 16940 14892 16946 14904
rect 18004 14876 18032 14904
rect 23414 14892 23420 14944
rect 23472 14932 23478 14944
rect 23785 14935 23843 14941
rect 23785 14932 23797 14935
rect 23472 14904 23797 14932
rect 23472 14892 23478 14904
rect 23785 14901 23797 14904
rect 23831 14932 23843 14935
rect 24058 14932 24064 14944
rect 23831 14904 24064 14932
rect 23831 14901 23843 14904
rect 23785 14895 23843 14901
rect 24058 14892 24064 14904
rect 24116 14892 24122 14944
rect 24334 14932 24340 14944
rect 24295 14904 24340 14932
rect 24334 14892 24340 14904
rect 24392 14892 24398 14944
rect 24613 14935 24671 14941
rect 24613 14901 24625 14935
rect 24659 14932 24671 14935
rect 25806 14932 25812 14944
rect 24659 14904 25812 14932
rect 24659 14901 24671 14904
rect 24613 14895 24671 14901
rect 25806 14892 25812 14904
rect 25864 14892 25870 14944
rect 5385 14867 5443 14873
rect 5385 14833 5397 14867
rect 5431 14833 5443 14867
rect 6118 14864 6124 14876
rect 5385 14827 5443 14833
rect 5492 14836 6124 14864
rect 3266 14756 3272 14808
rect 3324 14796 3330 14808
rect 3361 14799 3419 14805
rect 3361 14796 3373 14799
rect 3324 14768 3373 14796
rect 3324 14756 3330 14768
rect 3361 14765 3373 14768
rect 3407 14765 3419 14799
rect 3361 14759 3419 14765
rect 5109 14799 5167 14805
rect 5109 14765 5121 14799
rect 5155 14796 5167 14799
rect 5492 14796 5520 14836
rect 6118 14824 6124 14836
rect 6176 14824 6182 14876
rect 6397 14867 6455 14873
rect 6397 14833 6409 14867
rect 6443 14864 6455 14867
rect 6854 14864 6860 14876
rect 6443 14836 6860 14864
rect 6443 14833 6455 14836
rect 6397 14827 6455 14833
rect 6854 14824 6860 14836
rect 6912 14824 6918 14876
rect 7317 14867 7375 14873
rect 7317 14833 7329 14867
rect 7363 14864 7375 14867
rect 8418 14864 8424 14876
rect 7363 14836 8424 14864
rect 7363 14833 7375 14836
rect 7317 14827 7375 14833
rect 8418 14824 8424 14836
rect 8476 14824 8482 14876
rect 8970 14864 8976 14876
rect 8931 14836 8976 14864
rect 8970 14824 8976 14836
rect 9028 14824 9034 14876
rect 9062 14824 9068 14876
rect 9120 14864 9126 14876
rect 9157 14867 9215 14873
rect 9157 14864 9169 14867
rect 9120 14836 9169 14864
rect 9120 14824 9126 14836
rect 9157 14833 9169 14836
rect 9203 14833 9215 14867
rect 9157 14827 9215 14833
rect 11365 14867 11423 14873
rect 11365 14833 11377 14867
rect 11411 14864 11423 14867
rect 11638 14864 11644 14876
rect 11411 14836 11644 14864
rect 11411 14833 11423 14836
rect 11365 14827 11423 14833
rect 11638 14824 11644 14836
rect 11696 14824 11702 14876
rect 16422 14824 16428 14876
rect 16480 14864 16486 14876
rect 16977 14867 17035 14873
rect 16977 14864 16989 14867
rect 16480 14836 16989 14864
rect 16480 14824 16486 14836
rect 16977 14833 16989 14836
rect 17023 14833 17035 14867
rect 17158 14864 17164 14876
rect 17119 14836 17164 14864
rect 16977 14827 17035 14833
rect 17158 14824 17164 14836
rect 17216 14824 17222 14876
rect 17986 14864 17992 14876
rect 17899 14836 17992 14864
rect 17986 14824 17992 14836
rect 18044 14824 18050 14876
rect 22770 14864 22776 14876
rect 22731 14836 22776 14864
rect 22770 14824 22776 14836
rect 22828 14824 22834 14876
rect 22957 14867 23015 14873
rect 22957 14833 22969 14867
rect 23003 14864 23015 14867
rect 23046 14864 23052 14876
rect 23003 14836 23052 14864
rect 23003 14833 23015 14836
rect 22957 14827 23015 14833
rect 23046 14824 23052 14836
rect 23104 14824 23110 14876
rect 23322 14864 23328 14876
rect 23283 14836 23328 14864
rect 23322 14824 23328 14836
rect 23380 14824 23386 14876
rect 23690 14824 23696 14876
rect 23748 14864 23754 14876
rect 24352 14864 24380 14892
rect 23748 14836 24380 14864
rect 23748 14824 23754 14836
rect 5155 14768 5520 14796
rect 5155 14765 5167 14768
rect 5109 14759 5167 14765
rect 5750 14756 5756 14808
rect 5808 14796 5814 14808
rect 5845 14799 5903 14805
rect 5845 14796 5857 14799
rect 5808 14768 5857 14796
rect 5808 14756 5814 14768
rect 5845 14765 5857 14768
rect 5891 14765 5903 14799
rect 5845 14759 5903 14765
rect 6946 14756 6952 14808
rect 7004 14796 7010 14808
rect 7406 14796 7412 14808
rect 7004 14768 7412 14796
rect 7004 14756 7010 14768
rect 7406 14756 7412 14768
rect 7464 14796 7470 14808
rect 7685 14799 7743 14805
rect 7685 14796 7697 14799
rect 7464 14768 7697 14796
rect 7464 14756 7470 14768
rect 7685 14765 7697 14768
rect 7731 14796 7743 14799
rect 8510 14796 8516 14808
rect 7731 14768 8516 14796
rect 7731 14765 7743 14768
rect 7685 14759 7743 14765
rect 8510 14756 8516 14768
rect 8568 14756 8574 14808
rect 9338 14756 9344 14808
rect 9396 14796 9402 14808
rect 10718 14796 10724 14808
rect 9396 14768 10724 14796
rect 9396 14756 9402 14768
rect 10718 14756 10724 14768
rect 10776 14756 10782 14808
rect 11733 14799 11791 14805
rect 11733 14765 11745 14799
rect 11779 14796 11791 14799
rect 12190 14796 12196 14808
rect 11779 14768 12196 14796
rect 11779 14765 11791 14768
rect 11733 14759 11791 14765
rect 12190 14756 12196 14768
rect 12248 14756 12254 14808
rect 16146 14796 16152 14808
rect 16107 14768 16152 14796
rect 16146 14756 16152 14768
rect 16204 14756 16210 14808
rect 16606 14756 16612 14808
rect 16664 14796 16670 14808
rect 16701 14799 16759 14805
rect 16701 14796 16713 14799
rect 16664 14768 16713 14796
rect 16664 14756 16670 14768
rect 16701 14765 16713 14768
rect 16747 14765 16759 14799
rect 22310 14796 22316 14808
rect 22271 14768 22316 14796
rect 16701 14759 16759 14765
rect 22310 14756 22316 14768
rect 22368 14756 22374 14808
rect 23230 14796 23236 14808
rect 23191 14768 23236 14796
rect 23230 14756 23236 14768
rect 23288 14756 23294 14808
rect 4094 14688 4100 14740
rect 4152 14728 4158 14740
rect 5198 14728 5204 14740
rect 4152 14700 5204 14728
rect 4152 14688 4158 14700
rect 5198 14688 5204 14700
rect 5256 14688 5262 14740
rect 6486 14688 6492 14740
rect 6544 14728 6550 14740
rect 6762 14728 6768 14740
rect 6544 14700 6768 14728
rect 6544 14688 6550 14700
rect 6762 14688 6768 14700
rect 6820 14728 6826 14740
rect 11546 14737 11552 14740
rect 7593 14731 7651 14737
rect 7593 14728 7605 14731
rect 6820 14700 7605 14728
rect 6820 14688 6826 14700
rect 7593 14697 7605 14700
rect 7639 14697 7651 14731
rect 11530 14731 11552 14737
rect 11530 14728 11542 14731
rect 11459 14700 11542 14728
rect 7593 14691 7651 14697
rect 11530 14697 11542 14700
rect 11604 14728 11610 14740
rect 12377 14731 12435 14737
rect 12377 14728 12389 14731
rect 11604 14700 12389 14728
rect 11530 14691 11552 14697
rect 11546 14688 11552 14691
rect 11604 14688 11610 14700
rect 12377 14697 12389 14700
rect 12423 14728 12435 14731
rect 12926 14728 12932 14740
rect 12423 14700 12932 14728
rect 12423 14697 12435 14700
rect 12377 14691 12435 14697
rect 12926 14688 12932 14700
rect 12984 14688 12990 14740
rect 2349 14663 2407 14669
rect 2349 14629 2361 14663
rect 2395 14660 2407 14663
rect 2438 14660 2444 14672
rect 2395 14632 2444 14660
rect 2395 14629 2407 14632
rect 2349 14623 2407 14629
rect 2438 14620 2444 14632
rect 2496 14660 2502 14672
rect 3082 14660 3088 14672
rect 2496 14632 3088 14660
rect 2496 14620 2502 14632
rect 3082 14620 3088 14632
rect 3140 14660 3146 14672
rect 3637 14663 3695 14669
rect 3637 14660 3649 14663
rect 3140 14632 3649 14660
rect 3140 14620 3146 14632
rect 3637 14629 3649 14632
rect 3683 14629 3695 14663
rect 3637 14623 3695 14629
rect 5842 14620 5848 14672
rect 5900 14660 5906 14672
rect 6121 14663 6179 14669
rect 6121 14660 6133 14663
rect 5900 14632 6133 14660
rect 5900 14620 5906 14632
rect 6121 14629 6133 14632
rect 6167 14660 6179 14663
rect 6394 14660 6400 14672
rect 6167 14632 6400 14660
rect 6167 14629 6179 14632
rect 6121 14623 6179 14629
rect 6394 14620 6400 14632
rect 6452 14620 6458 14672
rect 6854 14620 6860 14672
rect 6912 14660 6918 14672
rect 7222 14660 7228 14672
rect 6912 14632 7228 14660
rect 6912 14620 6918 14632
rect 7222 14620 7228 14632
rect 7280 14660 7286 14672
rect 7455 14663 7513 14669
rect 7455 14660 7467 14663
rect 7280 14632 7467 14660
rect 7280 14620 7286 14632
rect 7455 14629 7467 14632
rect 7501 14629 7513 14663
rect 7455 14623 7513 14629
rect 7774 14620 7780 14672
rect 7832 14660 7838 14672
rect 7961 14663 8019 14669
rect 7961 14660 7973 14663
rect 7832 14632 7973 14660
rect 7832 14620 7838 14632
rect 7961 14629 7973 14632
rect 8007 14660 8019 14663
rect 8602 14660 8608 14672
rect 8007 14632 8608 14660
rect 8007 14629 8019 14632
rect 7961 14623 8019 14629
rect 8602 14620 8608 14632
rect 8660 14620 8666 14672
rect 8786 14620 8792 14672
rect 8844 14660 8850 14672
rect 9249 14663 9307 14669
rect 9249 14660 9261 14663
rect 8844 14632 9261 14660
rect 8844 14620 8850 14632
rect 9249 14629 9261 14632
rect 9295 14660 9307 14663
rect 9338 14660 9344 14672
rect 9295 14632 9344 14660
rect 9295 14629 9307 14632
rect 9249 14623 9307 14629
rect 9338 14620 9344 14632
rect 9396 14620 9402 14672
rect 9430 14620 9436 14672
rect 9488 14660 9494 14672
rect 9798 14660 9804 14672
rect 9488 14632 9804 14660
rect 9488 14620 9494 14632
rect 9798 14620 9804 14632
rect 9856 14660 9862 14672
rect 9893 14663 9951 14669
rect 9893 14660 9905 14663
rect 9856 14632 9905 14660
rect 9856 14620 9862 14632
rect 9893 14629 9905 14632
rect 9939 14629 9951 14663
rect 9893 14623 9951 14629
rect 10169 14663 10227 14669
rect 10169 14629 10181 14663
rect 10215 14660 10227 14663
rect 10626 14660 10632 14672
rect 10215 14632 10632 14660
rect 10215 14629 10227 14632
rect 10169 14623 10227 14629
rect 10626 14620 10632 14632
rect 10684 14620 10690 14672
rect 11641 14663 11699 14669
rect 11641 14629 11653 14663
rect 11687 14660 11699 14663
rect 11730 14660 11736 14672
rect 11687 14632 11736 14660
rect 11687 14629 11699 14632
rect 11641 14623 11699 14629
rect 11730 14620 11736 14632
rect 11788 14620 11794 14672
rect 17434 14620 17440 14672
rect 17492 14660 17498 14672
rect 17805 14663 17863 14669
rect 17805 14660 17817 14663
rect 17492 14632 17817 14660
rect 17492 14620 17498 14632
rect 17805 14629 17817 14632
rect 17851 14660 17863 14663
rect 18265 14663 18323 14669
rect 18265 14660 18277 14663
rect 17851 14632 18277 14660
rect 17851 14629 17863 14632
rect 17805 14623 17863 14629
rect 18265 14629 18277 14632
rect 18311 14660 18323 14663
rect 18722 14660 18728 14672
rect 18311 14632 18728 14660
rect 18311 14629 18323 14632
rect 18265 14623 18323 14629
rect 18722 14620 18728 14632
rect 18780 14620 18786 14672
rect 19829 14663 19887 14669
rect 19829 14629 19841 14663
rect 19875 14660 19887 14663
rect 20470 14660 20476 14672
rect 19875 14632 20476 14660
rect 19875 14629 19887 14632
rect 19829 14623 19887 14629
rect 20470 14620 20476 14632
rect 20528 14620 20534 14672
rect 400 14570 27264 14592
rect 400 14518 3510 14570
rect 3562 14518 3574 14570
rect 3626 14518 3638 14570
rect 3690 14518 3702 14570
rect 3754 14518 3766 14570
rect 3818 14518 27264 14570
rect 400 14496 27264 14518
rect 1521 14459 1579 14465
rect 1521 14425 1533 14459
rect 1567 14456 1579 14459
rect 2257 14459 2315 14465
rect 2257 14456 2269 14459
rect 1567 14428 2269 14456
rect 1567 14425 1579 14428
rect 1521 14419 1579 14425
rect 2257 14425 2269 14428
rect 2303 14456 2315 14459
rect 3082 14456 3088 14468
rect 2303 14428 3088 14456
rect 2303 14425 2315 14428
rect 2257 14419 2315 14425
rect 3082 14416 3088 14428
rect 3140 14416 3146 14468
rect 3358 14416 3364 14468
rect 3416 14456 3422 14468
rect 3545 14459 3603 14465
rect 3545 14456 3557 14459
rect 3416 14428 3557 14456
rect 3416 14416 3422 14428
rect 3545 14425 3557 14428
rect 3591 14425 3603 14459
rect 3545 14419 3603 14425
rect 3821 14459 3879 14465
rect 3821 14425 3833 14459
rect 3867 14456 3879 14459
rect 4078 14459 4136 14465
rect 4078 14456 4090 14459
rect 3867 14428 4090 14456
rect 3867 14425 3879 14428
rect 3821 14419 3879 14425
rect 4078 14425 4090 14428
rect 4124 14456 4136 14459
rect 4124 14428 4324 14456
rect 4124 14425 4136 14428
rect 4078 14419 4136 14425
rect 1150 14348 1156 14400
rect 1208 14388 1214 14400
rect 1337 14391 1395 14397
rect 1337 14388 1349 14391
rect 1208 14360 1349 14388
rect 1208 14348 1214 14360
rect 1337 14357 1349 14360
rect 1383 14388 1395 14391
rect 1794 14388 1800 14400
rect 1383 14360 1800 14388
rect 1383 14357 1395 14360
rect 1337 14351 1395 14357
rect 1794 14348 1800 14360
rect 1852 14348 1858 14400
rect 1889 14391 1947 14397
rect 1889 14357 1901 14391
rect 1935 14388 1947 14391
rect 4186 14388 4192 14400
rect 1935 14360 2392 14388
rect 4147 14360 4192 14388
rect 1935 14357 1947 14360
rect 1889 14351 1947 14357
rect 2364 14329 2392 14360
rect 4186 14348 4192 14360
rect 4244 14348 4250 14400
rect 4296 14388 4324 14428
rect 4554 14416 4560 14468
rect 4612 14456 4618 14468
rect 4612 14428 4657 14456
rect 4612 14416 4618 14428
rect 5014 14416 5020 14468
rect 5072 14456 5078 14468
rect 6486 14456 6492 14468
rect 5072 14428 6492 14456
rect 5072 14416 5078 14428
rect 6486 14416 6492 14428
rect 6544 14416 6550 14468
rect 6765 14459 6823 14465
rect 6765 14425 6777 14459
rect 6811 14456 6823 14459
rect 6854 14456 6860 14468
rect 6811 14428 6860 14456
rect 6811 14425 6823 14428
rect 6765 14419 6823 14425
rect 6854 14416 6860 14428
rect 6912 14416 6918 14468
rect 6946 14416 6952 14468
rect 7004 14456 7010 14468
rect 8418 14456 8424 14468
rect 7004 14428 7049 14456
rect 8379 14428 8424 14456
rect 7004 14416 7010 14428
rect 8418 14416 8424 14428
rect 8476 14416 8482 14468
rect 8602 14456 8608 14468
rect 8563 14428 8608 14456
rect 8602 14416 8608 14428
rect 8660 14416 8666 14468
rect 8970 14416 8976 14468
rect 9028 14456 9034 14468
rect 9157 14459 9215 14465
rect 9157 14456 9169 14459
rect 9028 14428 9169 14456
rect 9028 14416 9034 14428
rect 9157 14425 9169 14428
rect 9203 14425 9215 14459
rect 9338 14456 9344 14468
rect 9299 14428 9344 14456
rect 9157 14419 9215 14425
rect 9338 14416 9344 14428
rect 9396 14416 9402 14468
rect 9522 14456 9528 14468
rect 9483 14428 9528 14456
rect 9522 14416 9528 14428
rect 9580 14456 9586 14468
rect 9982 14456 9988 14468
rect 9580 14428 9988 14456
rect 9580 14416 9586 14428
rect 9982 14416 9988 14428
rect 10040 14416 10046 14468
rect 10718 14456 10724 14468
rect 10679 14428 10724 14456
rect 10718 14416 10724 14428
rect 10776 14416 10782 14468
rect 11362 14416 11368 14468
rect 11420 14456 11426 14468
rect 12098 14456 12104 14468
rect 11420 14428 12104 14456
rect 11420 14416 11426 14428
rect 12098 14416 12104 14428
rect 12156 14456 12162 14468
rect 12193 14459 12251 14465
rect 12193 14456 12205 14459
rect 12156 14428 12205 14456
rect 12156 14416 12162 14428
rect 12193 14425 12205 14428
rect 12239 14425 12251 14459
rect 12926 14456 12932 14468
rect 12887 14428 12932 14456
rect 12193 14419 12251 14425
rect 12926 14416 12932 14428
rect 12984 14416 12990 14468
rect 13570 14416 13576 14468
rect 13628 14456 13634 14468
rect 13849 14459 13907 14465
rect 13849 14456 13861 14459
rect 13628 14428 13861 14456
rect 13628 14416 13634 14428
rect 13849 14425 13861 14428
rect 13895 14425 13907 14459
rect 13849 14419 13907 14425
rect 16146 14416 16152 14468
rect 16204 14456 16210 14468
rect 16701 14459 16759 14465
rect 16701 14456 16713 14459
rect 16204 14428 16713 14456
rect 16204 14416 16210 14428
rect 16701 14425 16713 14428
rect 16747 14456 16759 14459
rect 17069 14459 17127 14465
rect 17069 14456 17081 14459
rect 16747 14428 17081 14456
rect 16747 14425 16759 14428
rect 16701 14419 16759 14425
rect 17069 14425 17081 14428
rect 17115 14425 17127 14459
rect 17434 14456 17440 14468
rect 17395 14428 17440 14456
rect 17069 14419 17127 14425
rect 6578 14388 6584 14400
rect 4296 14360 6584 14388
rect 6578 14348 6584 14360
rect 6636 14348 6642 14400
rect 7498 14388 7504 14400
rect 7411 14360 7504 14388
rect 7498 14348 7504 14360
rect 7556 14388 7562 14400
rect 8237 14391 8295 14397
rect 8237 14388 8249 14391
rect 7556 14360 8249 14388
rect 7556 14348 7562 14360
rect 8237 14357 8249 14360
rect 8283 14357 8295 14391
rect 8237 14351 8295 14357
rect 2128 14323 2186 14329
rect 2128 14320 2140 14323
rect 1720 14292 2140 14320
rect 1720 14252 1748 14292
rect 2128 14289 2140 14292
rect 2174 14289 2186 14323
rect 2128 14283 2186 14289
rect 2349 14323 2407 14329
rect 2349 14289 2361 14323
rect 2395 14320 2407 14323
rect 2714 14320 2720 14332
rect 2395 14292 2720 14320
rect 2395 14289 2407 14292
rect 2349 14283 2407 14289
rect 2714 14280 2720 14292
rect 2772 14280 2778 14332
rect 4281 14323 4339 14329
rect 4281 14289 4293 14323
rect 4327 14320 4339 14323
rect 4370 14320 4376 14332
rect 4327 14292 4376 14320
rect 4327 14289 4339 14292
rect 4281 14283 4339 14289
rect 4370 14280 4376 14292
rect 4428 14280 4434 14332
rect 5106 14320 5112 14332
rect 5067 14292 5112 14320
rect 5106 14280 5112 14292
rect 5164 14280 5170 14332
rect 7372 14323 7430 14329
rect 7372 14320 7384 14323
rect 6320 14292 7384 14320
rect 1628 14224 1748 14252
rect 1334 14076 1340 14128
rect 1392 14116 1398 14128
rect 1628 14125 1656 14224
rect 1794 14212 1800 14264
rect 1852 14252 1858 14264
rect 3082 14252 3088 14264
rect 1852 14224 3088 14252
rect 1852 14212 1858 14224
rect 1978 14184 1984 14196
rect 1891 14156 1984 14184
rect 1978 14144 1984 14156
rect 2036 14144 2042 14196
rect 2732 14193 2760 14224
rect 3082 14212 3088 14224
rect 3140 14212 3146 14264
rect 5750 14252 5756 14264
rect 5711 14224 5756 14252
rect 5750 14212 5756 14224
rect 5808 14212 5814 14264
rect 2717 14187 2775 14193
rect 2717 14153 2729 14187
rect 2763 14153 2775 14187
rect 3913 14187 3971 14193
rect 3913 14184 3925 14187
rect 2717 14147 2775 14153
rect 3008 14156 3925 14184
rect 1613 14119 1671 14125
rect 1613 14116 1625 14119
rect 1392 14088 1625 14116
rect 1392 14076 1398 14088
rect 1613 14085 1625 14088
rect 1659 14085 1671 14119
rect 1996 14116 2024 14144
rect 3008 14128 3036 14156
rect 3913 14153 3925 14156
rect 3959 14184 3971 14187
rect 4741 14187 4799 14193
rect 4741 14184 4753 14187
rect 3959 14156 4753 14184
rect 3959 14153 3971 14156
rect 3913 14147 3971 14153
rect 4741 14153 4753 14156
rect 4787 14153 4799 14187
rect 4741 14147 4799 14153
rect 2809 14119 2867 14125
rect 2809 14116 2821 14119
rect 1996 14088 2821 14116
rect 1613 14079 1671 14085
rect 2809 14085 2821 14088
rect 2855 14116 2867 14119
rect 2990 14116 2996 14128
rect 2855 14088 2996 14116
rect 2855 14085 2867 14088
rect 2809 14079 2867 14085
rect 2990 14076 2996 14088
rect 3048 14076 3054 14128
rect 3266 14116 3272 14128
rect 3227 14088 3272 14116
rect 3266 14076 3272 14088
rect 3324 14076 3330 14128
rect 3358 14076 3364 14128
rect 3416 14116 3422 14128
rect 5382 14116 5388 14128
rect 3416 14088 3461 14116
rect 5343 14088 5388 14116
rect 3416 14076 3422 14088
rect 5382 14076 5388 14088
rect 5440 14076 5446 14128
rect 5569 14119 5627 14125
rect 5569 14085 5581 14119
rect 5615 14116 5627 14119
rect 5750 14116 5756 14128
rect 5615 14088 5756 14116
rect 5615 14085 5627 14088
rect 5569 14079 5627 14085
rect 5750 14076 5756 14088
rect 5808 14076 5814 14128
rect 5937 14119 5995 14125
rect 5937 14085 5949 14119
rect 5983 14116 5995 14119
rect 6118 14116 6124 14128
rect 5983 14088 6124 14116
rect 5983 14085 5995 14088
rect 5937 14079 5995 14085
rect 6118 14076 6124 14088
rect 6176 14076 6182 14128
rect 6210 14076 6216 14128
rect 6268 14116 6274 14128
rect 6320 14125 6348 14292
rect 7372 14289 7384 14292
rect 7418 14289 7430 14323
rect 7372 14283 7430 14289
rect 7593 14323 7651 14329
rect 7593 14289 7605 14323
rect 7639 14320 7651 14323
rect 8050 14320 8056 14332
rect 7639 14292 8056 14320
rect 7639 14289 7651 14292
rect 7593 14283 7651 14289
rect 8050 14280 8056 14292
rect 8108 14320 8114 14332
rect 8988 14320 9016 14416
rect 9062 14348 9068 14400
rect 9120 14388 9126 14400
rect 10074 14388 10080 14400
rect 9120 14360 10080 14388
rect 9120 14348 9126 14360
rect 10074 14348 10080 14360
rect 10132 14348 10138 14400
rect 10166 14348 10172 14400
rect 10224 14388 10230 14400
rect 11546 14388 11552 14400
rect 10224 14360 11552 14388
rect 10224 14348 10230 14360
rect 11546 14348 11552 14360
rect 11604 14388 11610 14400
rect 11871 14391 11929 14397
rect 11871 14388 11883 14391
rect 11604 14360 11883 14388
rect 11604 14348 11610 14360
rect 11871 14357 11883 14360
rect 11917 14357 11929 14391
rect 12006 14388 12012 14400
rect 11967 14360 12012 14388
rect 11871 14351 11929 14357
rect 12006 14348 12012 14360
rect 12064 14348 12070 14400
rect 16422 14388 16428 14400
rect 16383 14360 16428 14388
rect 16422 14348 16428 14360
rect 16480 14348 16486 14400
rect 16606 14388 16612 14400
rect 16567 14360 16612 14388
rect 16606 14348 16612 14360
rect 16664 14348 16670 14400
rect 8108 14292 9016 14320
rect 10629 14323 10687 14329
rect 8108 14280 8114 14292
rect 10629 14289 10641 14323
rect 10675 14320 10687 14323
rect 11270 14320 11276 14332
rect 10675 14292 11276 14320
rect 10675 14289 10687 14292
rect 10629 14283 10687 14289
rect 11270 14280 11276 14292
rect 11328 14280 11334 14332
rect 11454 14280 11460 14332
rect 11512 14320 11518 14332
rect 12101 14323 12159 14329
rect 12101 14320 12113 14323
rect 11512 14292 12113 14320
rect 11512 14280 11518 14292
rect 12101 14289 12113 14292
rect 12147 14320 12159 14323
rect 12561 14323 12619 14329
rect 12561 14320 12573 14323
rect 12147 14292 12573 14320
rect 12147 14289 12159 14292
rect 12101 14283 12159 14289
rect 12561 14289 12573 14292
rect 12607 14289 12619 14323
rect 12561 14283 12619 14289
rect 7130 14252 7136 14264
rect 7043 14224 7136 14252
rect 7130 14212 7136 14224
rect 7188 14252 7194 14264
rect 7225 14255 7283 14261
rect 7225 14252 7237 14255
rect 7188 14224 7237 14252
rect 7188 14212 7194 14224
rect 7225 14221 7237 14224
rect 7271 14221 7283 14255
rect 7225 14215 7283 14221
rect 9522 14212 9528 14264
rect 9580 14252 9586 14264
rect 9893 14255 9951 14261
rect 9893 14252 9905 14255
rect 9580 14224 9905 14252
rect 9580 14212 9586 14224
rect 9893 14221 9905 14224
rect 9939 14221 9951 14255
rect 9893 14215 9951 14221
rect 9982 14212 9988 14264
rect 10040 14212 10046 14264
rect 10169 14255 10227 14261
rect 10169 14221 10181 14255
rect 10215 14252 10227 14255
rect 10442 14252 10448 14264
rect 10215 14224 10448 14252
rect 10215 14221 10227 14224
rect 10169 14215 10227 14221
rect 10442 14212 10448 14224
rect 10500 14252 10506 14264
rect 10718 14252 10724 14264
rect 10500 14224 10724 14252
rect 10500 14212 10506 14224
rect 10718 14212 10724 14224
rect 10776 14212 10782 14264
rect 10902 14212 10908 14264
rect 10960 14252 10966 14264
rect 11546 14252 11552 14264
rect 10960 14224 11552 14252
rect 10960 14212 10966 14224
rect 11546 14212 11552 14224
rect 11604 14212 11610 14264
rect 13570 14252 13576 14264
rect 13531 14224 13576 14252
rect 13570 14212 13576 14224
rect 13628 14212 13634 14264
rect 17084 14252 17112 14419
rect 17434 14416 17440 14428
rect 17492 14416 17498 14468
rect 22589 14459 22647 14465
rect 22589 14425 22601 14459
rect 22635 14456 22647 14459
rect 23230 14456 23236 14468
rect 22635 14428 23236 14456
rect 22635 14425 22647 14428
rect 22589 14419 22647 14425
rect 23230 14416 23236 14428
rect 23288 14416 23294 14468
rect 20194 14388 20200 14400
rect 18464 14360 20200 14388
rect 18464 14332 18492 14360
rect 20194 14348 20200 14360
rect 20252 14348 20258 14400
rect 20562 14388 20568 14400
rect 20523 14360 20568 14388
rect 20562 14348 20568 14360
rect 20620 14348 20626 14400
rect 22221 14391 22279 14397
rect 22221 14357 22233 14391
rect 22267 14388 22279 14391
rect 22773 14391 22831 14397
rect 22773 14388 22785 14391
rect 22267 14360 22785 14388
rect 22267 14357 22279 14360
rect 22221 14351 22279 14357
rect 22773 14357 22785 14360
rect 22819 14388 22831 14391
rect 23322 14388 23328 14400
rect 22819 14360 23328 14388
rect 22819 14357 22831 14360
rect 22773 14351 22831 14357
rect 23322 14348 23328 14360
rect 23380 14388 23386 14400
rect 23380 14360 23552 14388
rect 23380 14348 23386 14360
rect 18446 14320 18452 14332
rect 18359 14292 18452 14320
rect 18446 14280 18452 14292
rect 18504 14280 18510 14332
rect 19645 14323 19703 14329
rect 19645 14289 19657 14323
rect 19691 14320 19703 14323
rect 19918 14320 19924 14332
rect 19691 14292 19924 14320
rect 19691 14289 19703 14292
rect 19645 14283 19703 14289
rect 19918 14280 19924 14292
rect 19976 14280 19982 14332
rect 21666 14320 21672 14332
rect 20120 14292 21672 14320
rect 18357 14255 18415 14261
rect 18357 14252 18369 14255
rect 17084 14224 18369 14252
rect 18357 14221 18369 14224
rect 18403 14221 18415 14255
rect 18722 14252 18728 14264
rect 18683 14224 18728 14252
rect 18357 14215 18415 14221
rect 18722 14212 18728 14224
rect 18780 14212 18786 14264
rect 18909 14255 18967 14261
rect 18909 14221 18921 14255
rect 18955 14252 18967 14255
rect 19274 14252 19280 14264
rect 18955 14224 19280 14252
rect 18955 14221 18967 14224
rect 18909 14215 18967 14221
rect 19274 14212 19280 14224
rect 19332 14212 19338 14264
rect 20120 14261 20148 14292
rect 21666 14280 21672 14292
rect 21724 14320 21730 14332
rect 22957 14323 23015 14329
rect 22957 14320 22969 14323
rect 21724 14292 22969 14320
rect 21724 14280 21730 14292
rect 22957 14289 22969 14292
rect 23003 14320 23015 14323
rect 23414 14320 23420 14332
rect 23003 14292 23420 14320
rect 23003 14289 23015 14292
rect 22957 14283 23015 14289
rect 23414 14280 23420 14292
rect 23472 14280 23478 14332
rect 23524 14329 23552 14360
rect 23509 14323 23567 14329
rect 23509 14289 23521 14323
rect 23555 14289 23567 14323
rect 23509 14283 23567 14289
rect 23598 14280 23604 14332
rect 23656 14320 23662 14332
rect 23656 14292 24012 14320
rect 23656 14280 23662 14292
rect 19461 14255 19519 14261
rect 19461 14221 19473 14255
rect 19507 14252 19519 14255
rect 20105 14255 20163 14261
rect 20105 14252 20117 14255
rect 19507 14224 20117 14252
rect 19507 14221 19519 14224
rect 19461 14215 19519 14221
rect 20105 14221 20117 14224
rect 20151 14221 20163 14255
rect 20105 14215 20163 14221
rect 20470 14212 20476 14264
rect 20528 14252 20534 14264
rect 20565 14255 20623 14261
rect 20565 14252 20577 14255
rect 20528 14224 20577 14252
rect 20528 14212 20534 14224
rect 20565 14221 20577 14224
rect 20611 14221 20623 14255
rect 20565 14215 20623 14221
rect 22405 14255 22463 14261
rect 22405 14221 22417 14255
rect 22451 14252 22463 14255
rect 22770 14252 22776 14264
rect 22451 14224 22776 14252
rect 22451 14221 22463 14224
rect 22405 14215 22463 14221
rect 22770 14212 22776 14224
rect 22828 14212 22834 14264
rect 23782 14252 23788 14264
rect 23743 14224 23788 14252
rect 23782 14212 23788 14224
rect 23840 14212 23846 14264
rect 23984 14261 24012 14292
rect 24886 14280 24892 14332
rect 24944 14320 24950 14332
rect 25625 14323 25683 14329
rect 25625 14320 25637 14323
rect 24944 14292 25637 14320
rect 24944 14280 24950 14292
rect 25625 14289 25637 14292
rect 25671 14320 25683 14323
rect 26177 14323 26235 14329
rect 26177 14320 26189 14323
rect 25671 14292 26189 14320
rect 25671 14289 25683 14292
rect 25625 14283 25683 14289
rect 26177 14289 26189 14292
rect 26223 14289 26235 14323
rect 26177 14283 26235 14289
rect 23969 14255 24027 14261
rect 23969 14221 23981 14255
rect 24015 14252 24027 14255
rect 24061 14255 24119 14261
rect 24061 14252 24073 14255
rect 24015 14224 24073 14252
rect 24015 14221 24027 14224
rect 23969 14215 24027 14221
rect 24061 14221 24073 14224
rect 24107 14221 24119 14255
rect 24061 14215 24119 14221
rect 24426 14212 24432 14264
rect 24484 14252 24490 14264
rect 25441 14255 25499 14261
rect 25441 14252 25453 14255
rect 24484 14224 25453 14252
rect 24484 14212 24490 14224
rect 25441 14221 25453 14224
rect 25487 14252 25499 14255
rect 25990 14252 25996 14264
rect 25487 14224 25996 14252
rect 25487 14221 25499 14224
rect 25441 14215 25499 14221
rect 25990 14212 25996 14224
rect 26048 14212 26054 14264
rect 7682 14144 7688 14196
rect 7740 14184 7746 14196
rect 7961 14187 8019 14193
rect 7961 14184 7973 14187
rect 7740 14156 7973 14184
rect 7740 14144 7746 14156
rect 7961 14153 7973 14156
rect 8007 14184 8019 14187
rect 8789 14187 8847 14193
rect 8789 14184 8801 14187
rect 8007 14156 8801 14184
rect 8007 14153 8019 14156
rect 7961 14147 8019 14153
rect 8789 14153 8801 14156
rect 8835 14153 8847 14187
rect 10000 14184 10028 14212
rect 10261 14187 10319 14193
rect 10261 14184 10273 14187
rect 10000 14156 10273 14184
rect 8789 14147 8847 14153
rect 10261 14153 10273 14156
rect 10307 14184 10319 14187
rect 10350 14184 10356 14196
rect 10307 14156 10356 14184
rect 10307 14153 10319 14156
rect 10261 14147 10319 14153
rect 10350 14144 10356 14156
rect 10408 14144 10414 14196
rect 11089 14187 11147 14193
rect 11089 14153 11101 14187
rect 11135 14184 11147 14187
rect 11273 14187 11331 14193
rect 11273 14184 11285 14187
rect 11135 14156 11285 14184
rect 11135 14153 11147 14156
rect 11089 14147 11147 14153
rect 11273 14153 11285 14156
rect 11319 14184 11331 14187
rect 11730 14184 11736 14196
rect 11319 14156 11736 14184
rect 11319 14153 11331 14156
rect 11273 14147 11331 14153
rect 11730 14144 11736 14156
rect 11788 14144 11794 14196
rect 12834 14184 12840 14196
rect 12795 14156 12840 14184
rect 12834 14144 12840 14156
rect 12892 14144 12898 14196
rect 16241 14187 16299 14193
rect 16241 14153 16253 14187
rect 16287 14184 16299 14187
rect 17158 14184 17164 14196
rect 16287 14156 17164 14184
rect 16287 14153 16299 14156
rect 16241 14147 16299 14153
rect 17158 14144 17164 14156
rect 17216 14144 17222 14196
rect 17713 14187 17771 14193
rect 17713 14184 17725 14187
rect 17452 14156 17725 14184
rect 6305 14119 6363 14125
rect 6305 14116 6317 14119
rect 6268 14088 6317 14116
rect 6268 14076 6274 14088
rect 6305 14085 6317 14088
rect 6351 14085 6363 14119
rect 8050 14116 8056 14128
rect 8011 14088 8056 14116
rect 6305 14079 6363 14085
rect 8050 14076 8056 14088
rect 8108 14076 8114 14128
rect 9338 14076 9344 14128
rect 9396 14116 9402 14128
rect 9709 14119 9767 14125
rect 9709 14116 9721 14119
rect 9396 14088 9721 14116
rect 9396 14076 9402 14088
rect 9709 14085 9721 14088
rect 9755 14116 9767 14119
rect 10077 14119 10135 14125
rect 10077 14116 10089 14119
rect 9755 14088 10089 14116
rect 9755 14085 9767 14088
rect 9709 14079 9767 14085
rect 10077 14085 10089 14088
rect 10123 14116 10135 14119
rect 11457 14119 11515 14125
rect 11457 14116 11469 14119
rect 10123 14088 11469 14116
rect 10123 14085 10135 14088
rect 10077 14079 10135 14085
rect 11457 14085 11469 14088
rect 11503 14116 11515 14119
rect 11822 14116 11828 14128
rect 11503 14088 11828 14116
rect 11503 14085 11515 14088
rect 11457 14079 11515 14085
rect 11822 14076 11828 14088
rect 11880 14076 11886 14128
rect 13665 14119 13723 14125
rect 13665 14085 13677 14119
rect 13711 14116 13723 14119
rect 14030 14116 14036 14128
rect 13711 14088 14036 14116
rect 13711 14085 13723 14088
rect 13665 14079 13723 14085
rect 14030 14076 14036 14088
rect 14088 14076 14094 14128
rect 16977 14119 17035 14125
rect 16977 14085 16989 14119
rect 17023 14116 17035 14119
rect 17452 14116 17480 14156
rect 17713 14153 17725 14156
rect 17759 14184 17771 14187
rect 17802 14184 17808 14196
rect 17759 14156 17808 14184
rect 17759 14153 17771 14156
rect 17713 14147 17771 14153
rect 17802 14144 17808 14156
rect 17860 14144 17866 14196
rect 17023 14088 17480 14116
rect 17621 14119 17679 14125
rect 17023 14085 17035 14088
rect 16977 14079 17035 14085
rect 17621 14085 17633 14119
rect 17667 14116 17679 14119
rect 18446 14116 18452 14128
rect 17667 14088 18452 14116
rect 17667 14085 17679 14088
rect 17621 14079 17679 14085
rect 18446 14076 18452 14088
rect 18504 14076 18510 14128
rect 22037 14119 22095 14125
rect 22037 14085 22049 14119
rect 22083 14116 22095 14119
rect 23046 14116 23052 14128
rect 22083 14088 23052 14116
rect 22083 14085 22095 14088
rect 22037 14079 22095 14085
rect 23046 14076 23052 14088
rect 23104 14076 23110 14128
rect 400 14026 27264 14048
rect 400 13974 18870 14026
rect 18922 13974 18934 14026
rect 18986 13974 18998 14026
rect 19050 13974 19062 14026
rect 19114 13974 19126 14026
rect 19178 13974 27264 14026
rect 400 13952 27264 13974
rect 4278 13912 4284 13924
rect 4239 13884 4284 13912
rect 4278 13872 4284 13884
rect 4336 13872 4342 13924
rect 4370 13872 4376 13924
rect 4428 13912 4434 13924
rect 4741 13915 4799 13921
rect 4741 13912 4753 13915
rect 4428 13884 4753 13912
rect 4428 13872 4434 13884
rect 4741 13881 4753 13884
rect 4787 13912 4799 13915
rect 6302 13912 6308 13924
rect 4787 13884 6308 13912
rect 4787 13881 4799 13884
rect 4741 13875 4799 13881
rect 6302 13872 6308 13884
rect 6360 13912 6366 13924
rect 9706 13912 9712 13924
rect 6360 13884 9712 13912
rect 6360 13872 6366 13884
rect 9706 13872 9712 13884
rect 9764 13912 9770 13924
rect 9764 13884 10028 13912
rect 9764 13872 9770 13884
rect 10000 13856 10028 13884
rect 10074 13872 10080 13924
rect 10132 13912 10138 13924
rect 12098 13912 12104 13924
rect 10132 13884 10580 13912
rect 12059 13884 12104 13912
rect 10132 13872 10138 13884
rect 10552 13856 10580 13884
rect 12098 13872 12104 13884
rect 12156 13872 12162 13924
rect 17986 13912 17992 13924
rect 17947 13884 17992 13912
rect 17986 13872 17992 13884
rect 18044 13872 18050 13924
rect 18538 13872 18544 13924
rect 18596 13912 18602 13924
rect 19366 13912 19372 13924
rect 18596 13884 19372 13912
rect 18596 13872 18602 13884
rect 19366 13872 19372 13884
rect 19424 13872 19430 13924
rect 19829 13915 19887 13921
rect 19829 13881 19841 13915
rect 19875 13912 19887 13915
rect 20562 13912 20568 13924
rect 19875 13884 20568 13912
rect 19875 13881 19887 13884
rect 19829 13875 19887 13881
rect 4002 13844 4008 13856
rect 3915 13816 4008 13844
rect 4002 13804 4008 13816
rect 4060 13844 4066 13856
rect 5658 13844 5664 13856
rect 4060 13816 5664 13844
rect 4060 13804 4066 13816
rect 5658 13804 5664 13816
rect 5716 13804 5722 13856
rect 7406 13804 7412 13856
rect 7464 13844 7470 13856
rect 7593 13847 7651 13853
rect 7593 13844 7605 13847
rect 7464 13816 7605 13844
rect 7464 13804 7470 13816
rect 7593 13813 7605 13816
rect 7639 13813 7651 13847
rect 7593 13807 7651 13813
rect 7685 13847 7743 13853
rect 7685 13813 7697 13847
rect 7731 13844 7743 13847
rect 8050 13844 8056 13856
rect 7731 13816 8056 13844
rect 7731 13813 7743 13816
rect 7685 13807 7743 13813
rect 8050 13804 8056 13816
rect 8108 13804 8114 13856
rect 9982 13844 9988 13856
rect 9943 13816 9988 13844
rect 9982 13804 9988 13816
rect 10040 13804 10046 13856
rect 10169 13847 10227 13853
rect 10169 13813 10181 13847
rect 10215 13844 10227 13847
rect 10350 13844 10356 13856
rect 10215 13816 10356 13844
rect 10215 13813 10227 13816
rect 10169 13807 10227 13813
rect 10350 13804 10356 13816
rect 10408 13804 10414 13856
rect 10534 13844 10540 13856
rect 10447 13816 10540 13844
rect 10534 13804 10540 13816
rect 10592 13844 10598 13856
rect 18004 13844 18032 13872
rect 10592 13816 11592 13844
rect 18004 13816 18731 13844
rect 10592 13804 10598 13816
rect 1702 13736 1708 13788
rect 1760 13776 1766 13788
rect 1797 13779 1855 13785
rect 1797 13776 1809 13779
rect 1760 13748 1809 13776
rect 1760 13736 1766 13748
rect 1797 13745 1809 13748
rect 1843 13745 1855 13779
rect 1797 13739 1855 13745
rect 1981 13779 2039 13785
rect 1981 13745 1993 13779
rect 2027 13776 2039 13779
rect 2254 13776 2260 13788
rect 2027 13748 2260 13776
rect 2027 13745 2039 13748
rect 1981 13739 2039 13745
rect 2254 13736 2260 13748
rect 2312 13776 2318 13788
rect 4094 13776 4100 13788
rect 2312 13748 4100 13776
rect 2312 13736 2318 13748
rect 4094 13736 4100 13748
rect 4152 13776 4158 13788
rect 4189 13779 4247 13785
rect 4189 13776 4201 13779
rect 4152 13748 4201 13776
rect 4152 13736 4158 13748
rect 4189 13745 4201 13748
rect 4235 13745 4247 13779
rect 4189 13739 4247 13745
rect 6854 13736 6860 13788
rect 6912 13776 6918 13788
rect 7501 13779 7559 13785
rect 7501 13776 7513 13779
rect 6912 13748 7513 13776
rect 6912 13736 6918 13748
rect 7501 13745 7513 13748
rect 7547 13745 7559 13779
rect 7501 13739 7559 13745
rect 10074 13736 10080 13788
rect 10132 13776 10138 13788
rect 10442 13776 10448 13788
rect 10132 13748 10448 13776
rect 10132 13736 10138 13748
rect 10442 13736 10448 13748
rect 10500 13736 10506 13788
rect 11270 13736 11276 13788
rect 11328 13776 11334 13788
rect 11564 13785 11592 13816
rect 11365 13779 11423 13785
rect 11365 13776 11377 13779
rect 11328 13748 11377 13776
rect 11328 13736 11334 13748
rect 11365 13745 11377 13748
rect 11411 13745 11423 13779
rect 11365 13739 11423 13745
rect 11549 13779 11607 13785
rect 11549 13745 11561 13779
rect 11595 13745 11607 13779
rect 11549 13739 11607 13745
rect 15781 13779 15839 13785
rect 15781 13745 15793 13779
rect 15827 13745 15839 13779
rect 18538 13776 18544 13788
rect 18499 13748 18544 13776
rect 15781 13739 15839 13745
rect 3082 13668 3088 13720
rect 3140 13708 3146 13720
rect 5842 13708 5848 13720
rect 3140 13680 5848 13708
rect 3140 13668 3146 13680
rect 5842 13668 5848 13680
rect 5900 13668 5906 13720
rect 7317 13711 7375 13717
rect 7317 13677 7329 13711
rect 7363 13677 7375 13711
rect 7317 13671 7375 13677
rect 4186 13600 4192 13652
rect 4244 13640 4250 13652
rect 7332 13640 7360 13671
rect 7958 13668 7964 13720
rect 8016 13708 8022 13720
rect 8053 13711 8111 13717
rect 8053 13708 8065 13711
rect 8016 13680 8065 13708
rect 8016 13668 8022 13680
rect 8053 13677 8065 13680
rect 8099 13677 8111 13711
rect 8053 13671 8111 13677
rect 9522 13668 9528 13720
rect 9580 13708 9586 13720
rect 9801 13711 9859 13717
rect 9801 13708 9813 13711
rect 9580 13680 9813 13708
rect 9580 13668 9586 13680
rect 9801 13677 9813 13680
rect 9847 13677 9859 13711
rect 9801 13671 9859 13677
rect 9982 13668 9988 13720
rect 10040 13708 10046 13720
rect 12006 13708 12012 13720
rect 10040 13680 12012 13708
rect 10040 13668 10046 13680
rect 12006 13668 12012 13680
rect 12064 13708 12070 13720
rect 12193 13711 12251 13717
rect 12193 13708 12205 13711
rect 12064 13680 12205 13708
rect 12064 13668 12070 13680
rect 12193 13677 12205 13680
rect 12239 13708 12251 13711
rect 13938 13708 13944 13720
rect 12239 13680 13944 13708
rect 12239 13677 12251 13680
rect 12193 13671 12251 13677
rect 13938 13668 13944 13680
rect 13996 13708 14002 13720
rect 15796 13708 15824 13739
rect 18538 13736 18544 13748
rect 18596 13736 18602 13788
rect 18703 13785 18731 13816
rect 18688 13779 18746 13785
rect 18688 13745 18700 13779
rect 18734 13776 18746 13779
rect 18814 13776 18820 13788
rect 18734 13748 18820 13776
rect 18734 13745 18746 13748
rect 18688 13739 18746 13745
rect 18814 13736 18820 13748
rect 18872 13736 18878 13788
rect 15962 13708 15968 13720
rect 13996 13680 15968 13708
rect 13996 13668 14002 13680
rect 15962 13668 15968 13680
rect 16020 13668 16026 13720
rect 18446 13668 18452 13720
rect 18504 13708 18510 13720
rect 18909 13711 18967 13717
rect 18909 13708 18921 13711
rect 18504 13680 18921 13708
rect 18504 13668 18510 13680
rect 18909 13677 18921 13680
rect 18955 13677 18967 13711
rect 18909 13671 18967 13677
rect 8602 13640 8608 13652
rect 4244 13612 8608 13640
rect 4244 13600 4250 13612
rect 8602 13600 8608 13612
rect 8660 13640 8666 13652
rect 9154 13640 9160 13652
rect 8660 13612 9160 13640
rect 8660 13600 8666 13612
rect 9154 13600 9160 13612
rect 9212 13640 9218 13652
rect 11454 13640 11460 13652
rect 9212 13612 9936 13640
rect 9212 13600 9218 13612
rect 1334 13532 1340 13584
rect 1392 13572 1398 13584
rect 2073 13575 2131 13581
rect 2073 13572 2085 13575
rect 1392 13544 2085 13572
rect 1392 13532 1398 13544
rect 2073 13541 2085 13544
rect 2119 13541 2131 13575
rect 6118 13572 6124 13584
rect 6079 13544 6124 13572
rect 2073 13535 2131 13541
rect 6118 13532 6124 13544
rect 6176 13572 6182 13584
rect 7130 13572 7136 13584
rect 6176 13544 7136 13572
rect 6176 13532 6182 13544
rect 7130 13532 7136 13544
rect 7188 13532 7194 13584
rect 8142 13572 8148 13584
rect 8103 13544 8148 13572
rect 8142 13532 8148 13544
rect 8200 13532 8206 13584
rect 9246 13572 9252 13584
rect 9207 13544 9252 13572
rect 9246 13532 9252 13544
rect 9304 13532 9310 13584
rect 9908 13572 9936 13612
rect 10046 13612 11460 13640
rect 10046 13572 10074 13612
rect 11454 13600 11460 13612
rect 11512 13600 11518 13652
rect 11822 13600 11828 13652
rect 11880 13640 11886 13652
rect 15778 13640 15784 13652
rect 11880 13612 15784 13640
rect 11880 13600 11886 13612
rect 15778 13600 15784 13612
rect 15836 13640 15842 13652
rect 15873 13643 15931 13649
rect 15873 13640 15885 13643
rect 15836 13612 15885 13640
rect 15836 13600 15842 13612
rect 15873 13609 15885 13612
rect 15919 13609 15931 13643
rect 15873 13603 15931 13609
rect 18722 13600 18728 13652
rect 18780 13640 18786 13652
rect 18817 13643 18875 13649
rect 18817 13640 18829 13643
rect 18780 13612 18829 13640
rect 18780 13600 18786 13612
rect 18817 13609 18829 13612
rect 18863 13640 18875 13643
rect 19844 13640 19872 13875
rect 20562 13872 20568 13884
rect 20620 13872 20626 13924
rect 22310 13912 22316 13924
rect 22271 13884 22316 13912
rect 22310 13872 22316 13884
rect 22368 13872 22374 13924
rect 23046 13912 23052 13924
rect 23007 13884 23052 13912
rect 23046 13872 23052 13884
rect 23104 13872 23110 13924
rect 23414 13912 23420 13924
rect 23375 13884 23420 13912
rect 23414 13872 23420 13884
rect 23472 13872 23478 13924
rect 23693 13915 23751 13921
rect 23693 13881 23705 13915
rect 23739 13912 23751 13915
rect 23782 13912 23788 13924
rect 23739 13884 23788 13912
rect 23739 13881 23751 13884
rect 23693 13875 23751 13881
rect 23782 13872 23788 13884
rect 23840 13872 23846 13924
rect 20197 13847 20255 13853
rect 20197 13813 20209 13847
rect 20243 13844 20255 13847
rect 20470 13844 20476 13856
rect 20243 13816 20476 13844
rect 20243 13813 20255 13816
rect 20197 13807 20255 13813
rect 20470 13804 20476 13816
rect 20528 13804 20534 13856
rect 20378 13776 20384 13788
rect 20339 13748 20384 13776
rect 20378 13736 20384 13748
rect 20436 13736 20442 13788
rect 21666 13776 21672 13788
rect 21579 13748 21672 13776
rect 21666 13736 21672 13748
rect 21724 13776 21730 13788
rect 22126 13776 22132 13788
rect 21724 13748 22132 13776
rect 21724 13736 21730 13748
rect 22126 13736 22132 13748
rect 22184 13736 22190 13788
rect 23233 13779 23291 13785
rect 23233 13745 23245 13779
rect 23279 13776 23291 13779
rect 23322 13776 23328 13788
rect 23279 13748 23328 13776
rect 23279 13745 23291 13748
rect 23233 13739 23291 13745
rect 23322 13736 23328 13748
rect 23380 13736 23386 13788
rect 19918 13668 19924 13720
rect 19976 13708 19982 13720
rect 21577 13711 21635 13717
rect 21577 13708 21589 13711
rect 19976 13680 21589 13708
rect 19976 13668 19982 13680
rect 21577 13677 21589 13680
rect 21623 13708 21635 13711
rect 21942 13708 21948 13720
rect 21623 13680 21948 13708
rect 21623 13677 21635 13680
rect 21577 13671 21635 13677
rect 21942 13668 21948 13680
rect 22000 13668 22006 13720
rect 18863 13612 19872 13640
rect 18863 13609 18875 13612
rect 18817 13603 18875 13609
rect 11638 13572 11644 13584
rect 9908 13544 10074 13572
rect 11599 13544 11644 13572
rect 11638 13532 11644 13544
rect 11696 13532 11702 13584
rect 13294 13572 13300 13584
rect 13255 13544 13300 13572
rect 13294 13532 13300 13544
rect 13352 13532 13358 13584
rect 17805 13575 17863 13581
rect 17805 13541 17817 13575
rect 17851 13572 17863 13575
rect 18630 13572 18636 13584
rect 17851 13544 18636 13572
rect 17851 13541 17863 13544
rect 17805 13535 17863 13541
rect 18630 13532 18636 13544
rect 18688 13532 18694 13584
rect 19182 13572 19188 13584
rect 19143 13544 19188 13572
rect 19182 13532 19188 13544
rect 19240 13532 19246 13584
rect 19274 13532 19280 13584
rect 19332 13572 19338 13584
rect 20473 13575 20531 13581
rect 20473 13572 20485 13575
rect 19332 13544 20485 13572
rect 19332 13532 19338 13544
rect 20473 13541 20485 13544
rect 20519 13541 20531 13575
rect 20473 13535 20531 13541
rect 20933 13575 20991 13581
rect 20933 13541 20945 13575
rect 20979 13572 20991 13575
rect 21206 13572 21212 13584
rect 20979 13544 21212 13572
rect 20979 13541 20991 13544
rect 20933 13535 20991 13541
rect 21206 13532 21212 13544
rect 21264 13572 21270 13584
rect 21853 13575 21911 13581
rect 21853 13572 21865 13575
rect 21264 13544 21865 13572
rect 21264 13532 21270 13544
rect 21853 13541 21865 13544
rect 21899 13541 21911 13575
rect 21853 13535 21911 13541
rect 400 13482 27264 13504
rect 400 13430 3510 13482
rect 3562 13430 3574 13482
rect 3626 13430 3638 13482
rect 3690 13430 3702 13482
rect 3754 13430 3766 13482
rect 3818 13430 27264 13482
rect 400 13408 27264 13430
rect 1705 13371 1763 13377
rect 1705 13337 1717 13371
rect 1751 13368 1763 13371
rect 1889 13371 1947 13377
rect 1889 13368 1901 13371
rect 1751 13340 1901 13368
rect 1751 13337 1763 13340
rect 1705 13331 1763 13337
rect 1889 13337 1901 13340
rect 1935 13368 1947 13371
rect 2254 13368 2260 13380
rect 1935 13340 2260 13368
rect 1935 13337 1947 13340
rect 1889 13331 1947 13337
rect 2254 13328 2260 13340
rect 2312 13328 2318 13380
rect 2806 13368 2812 13380
rect 2767 13340 2812 13368
rect 2806 13328 2812 13340
rect 2864 13328 2870 13380
rect 3266 13368 3272 13380
rect 3227 13340 3272 13368
rect 3266 13328 3272 13340
rect 3324 13328 3330 13380
rect 3545 13371 3603 13377
rect 3545 13337 3557 13371
rect 3591 13368 3603 13371
rect 4002 13368 4008 13380
rect 3591 13340 4008 13368
rect 3591 13337 3603 13340
rect 3545 13331 3603 13337
rect 4002 13328 4008 13340
rect 4060 13328 4066 13380
rect 5106 13368 5112 13380
rect 5067 13340 5112 13368
rect 5106 13328 5112 13340
rect 5164 13328 5170 13380
rect 5569 13371 5627 13377
rect 5569 13337 5581 13371
rect 5615 13368 5627 13371
rect 6670 13368 6676 13380
rect 5615 13340 6676 13368
rect 5615 13337 5627 13340
rect 5569 13331 5627 13337
rect 6670 13328 6676 13340
rect 6728 13328 6734 13380
rect 6854 13328 6860 13380
rect 6912 13328 6918 13380
rect 7406 13368 7412 13380
rect 7367 13340 7412 13368
rect 7406 13328 7412 13340
rect 7464 13368 7470 13380
rect 7464 13340 7728 13368
rect 7464 13328 7470 13340
rect 2824 13300 2852 13328
rect 3637 13303 3695 13309
rect 3637 13300 3649 13303
rect 2824 13272 3649 13300
rect 2824 13232 2852 13272
rect 3637 13269 3649 13272
rect 3683 13300 3695 13303
rect 3683 13272 4416 13300
rect 3683 13269 3695 13272
rect 3637 13263 3695 13269
rect 1996 13204 2852 13232
rect 1996 13173 2024 13204
rect 3358 13192 3364 13244
rect 3416 13232 3422 13244
rect 4097 13235 4155 13241
rect 4097 13232 4109 13235
rect 3416 13204 4109 13232
rect 3416 13192 3422 13204
rect 4097 13201 4109 13204
rect 4143 13232 4155 13235
rect 4186 13232 4192 13244
rect 4143 13204 4192 13232
rect 4143 13201 4155 13204
rect 4097 13195 4155 13201
rect 4186 13192 4192 13204
rect 4244 13192 4250 13244
rect 4388 13232 4416 13272
rect 6302 13260 6308 13312
rect 6360 13300 6366 13312
rect 6872 13300 6900 13328
rect 6949 13303 7007 13309
rect 6949 13300 6961 13303
rect 6360 13272 6961 13300
rect 6360 13260 6366 13272
rect 6949 13269 6961 13272
rect 6995 13300 7007 13303
rect 7133 13303 7191 13309
rect 7133 13300 7145 13303
rect 6995 13272 7145 13300
rect 6995 13269 7007 13272
rect 6949 13263 7007 13269
rect 7133 13269 7145 13272
rect 7179 13269 7191 13303
rect 7700 13300 7728 13340
rect 7774 13328 7780 13380
rect 7832 13368 7838 13380
rect 7961 13371 8019 13377
rect 7961 13368 7973 13371
rect 7832 13340 7973 13368
rect 7832 13328 7838 13340
rect 7961 13337 7973 13340
rect 8007 13337 8019 13371
rect 7961 13331 8019 13337
rect 8142 13328 8148 13380
rect 8200 13368 8206 13380
rect 10074 13368 10080 13380
rect 8200 13340 8245 13368
rect 8344 13340 10080 13368
rect 8200 13328 8206 13340
rect 8344 13312 8372 13340
rect 10074 13328 10080 13340
rect 10132 13328 10138 13380
rect 10534 13368 10540 13380
rect 10495 13340 10540 13368
rect 10534 13328 10540 13340
rect 10592 13368 10598 13380
rect 11365 13371 11423 13377
rect 11365 13368 11377 13371
rect 10592 13340 11377 13368
rect 10592 13328 10598 13340
rect 11365 13337 11377 13340
rect 11411 13337 11423 13371
rect 15778 13368 15784 13380
rect 15739 13340 15784 13368
rect 11365 13331 11423 13337
rect 15778 13328 15784 13340
rect 15836 13328 15842 13380
rect 15962 13368 15968 13380
rect 15923 13340 15968 13368
rect 15962 13328 15968 13340
rect 16020 13328 16026 13380
rect 17802 13368 17808 13380
rect 17763 13340 17808 13368
rect 17802 13328 17808 13340
rect 17860 13328 17866 13380
rect 18446 13328 18452 13380
rect 18504 13368 18510 13380
rect 18541 13371 18599 13377
rect 18541 13368 18553 13371
rect 18504 13340 18553 13368
rect 18504 13328 18510 13340
rect 18541 13337 18553 13340
rect 18587 13337 18599 13371
rect 18722 13368 18728 13380
rect 18683 13340 18728 13368
rect 18541 13331 18599 13337
rect 18722 13328 18728 13340
rect 18780 13328 18786 13380
rect 18814 13328 18820 13380
rect 18872 13368 18878 13380
rect 18909 13371 18967 13377
rect 18909 13368 18921 13371
rect 18872 13340 18921 13368
rect 18872 13328 18878 13340
rect 18909 13337 18921 13340
rect 18955 13337 18967 13371
rect 18909 13331 18967 13337
rect 19185 13371 19243 13377
rect 19185 13337 19197 13371
rect 19231 13368 19243 13371
rect 19366 13368 19372 13380
rect 19231 13340 19372 13368
rect 19231 13337 19243 13340
rect 19185 13331 19243 13337
rect 19366 13328 19372 13340
rect 19424 13328 19430 13380
rect 20013 13371 20071 13377
rect 20013 13337 20025 13371
rect 20059 13368 20071 13371
rect 20470 13368 20476 13380
rect 20059 13340 20476 13368
rect 20059 13337 20071 13340
rect 20013 13331 20071 13337
rect 20470 13328 20476 13340
rect 20528 13328 20534 13380
rect 21942 13368 21948 13380
rect 21903 13340 21948 13368
rect 21942 13328 21948 13340
rect 22000 13328 22006 13380
rect 22126 13368 22132 13380
rect 22087 13340 22132 13368
rect 22126 13328 22132 13340
rect 22184 13328 22190 13380
rect 23046 13328 23052 13380
rect 23104 13368 23110 13380
rect 23141 13371 23199 13377
rect 23141 13368 23153 13371
rect 23104 13340 23153 13368
rect 23104 13328 23110 13340
rect 23141 13337 23153 13340
rect 23187 13337 23199 13371
rect 24061 13371 24119 13377
rect 24061 13368 24073 13371
rect 23141 13331 23199 13337
rect 23846 13340 24073 13368
rect 8326 13300 8332 13312
rect 7700 13272 8332 13300
rect 7133 13263 7191 13269
rect 8326 13260 8332 13272
rect 8384 13260 8390 13312
rect 8878 13260 8884 13312
rect 8936 13300 8942 13312
rect 9341 13303 9399 13309
rect 9341 13300 9353 13303
rect 8936 13272 9353 13300
rect 8936 13260 8942 13272
rect 9341 13269 9353 13272
rect 9387 13269 9399 13303
rect 9341 13263 9399 13269
rect 9798 13260 9804 13312
rect 9856 13300 9862 13312
rect 11181 13303 11239 13309
rect 11181 13300 11193 13303
rect 9856 13272 11193 13300
rect 9856 13260 9862 13272
rect 11181 13269 11193 13272
rect 11227 13300 11239 13303
rect 11270 13300 11276 13312
rect 11227 13272 11276 13300
rect 11227 13269 11239 13272
rect 11181 13263 11239 13269
rect 11270 13260 11276 13272
rect 11328 13260 11334 13312
rect 12929 13303 12987 13309
rect 12929 13269 12941 13303
rect 12975 13300 12987 13303
rect 17250 13300 17256 13312
rect 12975 13272 17256 13300
rect 12975 13269 12987 13272
rect 12929 13263 12987 13269
rect 4925 13235 4983 13241
rect 4925 13232 4937 13235
rect 4388 13204 4937 13232
rect 4925 13201 4937 13204
rect 4971 13201 4983 13235
rect 4925 13195 4983 13201
rect 7593 13235 7651 13241
rect 7593 13201 7605 13235
rect 7639 13232 7651 13235
rect 8053 13235 8111 13241
rect 7639 13204 8004 13232
rect 7639 13201 7651 13204
rect 7593 13195 7651 13201
rect 1981 13167 2039 13173
rect 1981 13133 1993 13167
rect 2027 13133 2039 13167
rect 1981 13127 2039 13133
rect 2165 13167 2223 13173
rect 2165 13133 2177 13167
rect 2211 13133 2223 13167
rect 2165 13127 2223 13133
rect 4465 13167 4523 13173
rect 4465 13133 4477 13167
rect 4511 13164 4523 13167
rect 4646 13164 4652 13176
rect 4511 13136 4652 13164
rect 4511 13133 4523 13136
rect 4465 13127 4523 13133
rect 1886 13056 1892 13108
rect 1944 13096 1950 13108
rect 2180 13096 2208 13127
rect 4646 13124 4652 13136
rect 4704 13164 4710 13176
rect 5106 13164 5112 13176
rect 4704 13136 5112 13164
rect 4704 13124 4710 13136
rect 5106 13124 5112 13136
rect 5164 13124 5170 13176
rect 5658 13164 5664 13176
rect 5619 13136 5664 13164
rect 5658 13124 5664 13136
rect 5716 13124 5722 13176
rect 5750 13124 5756 13176
rect 5808 13164 5814 13176
rect 5937 13167 5995 13173
rect 5937 13164 5949 13167
rect 5808 13136 5949 13164
rect 5808 13124 5814 13136
rect 5937 13133 5949 13136
rect 5983 13164 5995 13167
rect 7222 13164 7228 13176
rect 5983 13136 7228 13164
rect 5983 13133 5995 13136
rect 5937 13127 5995 13133
rect 2625 13099 2683 13105
rect 2625 13096 2637 13099
rect 1944 13068 2637 13096
rect 1944 13056 1950 13068
rect 2625 13065 2637 13068
rect 2671 13065 2683 13099
rect 2625 13059 2683 13065
rect 4370 13056 4376 13108
rect 4428 13096 4434 13108
rect 4554 13096 4560 13108
rect 4428 13068 4473 13096
rect 4515 13068 4560 13096
rect 4428 13056 4434 13068
rect 4554 13056 4560 13068
rect 4612 13056 4618 13108
rect 5290 13056 5296 13108
rect 5348 13096 5354 13108
rect 6118 13096 6124 13108
rect 5348 13068 6124 13096
rect 5348 13056 5354 13068
rect 6118 13056 6124 13068
rect 6176 13056 6182 13108
rect 6504 13105 6532 13136
rect 7222 13124 7228 13136
rect 7280 13124 7286 13176
rect 7682 13164 7688 13176
rect 7643 13136 7688 13164
rect 7682 13124 7688 13136
rect 7740 13124 7746 13176
rect 7832 13167 7890 13173
rect 7832 13133 7844 13167
rect 7878 13133 7890 13167
rect 7976 13164 8004 13204
rect 8053 13201 8065 13235
rect 8099 13232 8111 13235
rect 8513 13235 8571 13241
rect 8513 13232 8525 13235
rect 8099 13204 8525 13232
rect 8099 13201 8111 13204
rect 8053 13195 8111 13201
rect 8513 13201 8525 13204
rect 8559 13232 8571 13235
rect 10997 13235 11055 13241
rect 10997 13232 11009 13235
rect 8559 13204 11009 13232
rect 8559 13201 8571 13204
rect 8513 13195 8571 13201
rect 10997 13201 11009 13204
rect 11043 13201 11055 13235
rect 13386 13232 13392 13244
rect 13347 13204 13392 13232
rect 10997 13195 11055 13201
rect 8602 13164 8608 13176
rect 7976 13136 8608 13164
rect 7832 13127 7890 13133
rect 6489 13099 6547 13105
rect 6489 13065 6501 13099
rect 6535 13065 6547 13099
rect 6854 13096 6860 13108
rect 6767 13068 6860 13096
rect 6489 13059 6547 13065
rect 6854 13056 6860 13068
rect 6912 13096 6918 13108
rect 7498 13096 7504 13108
rect 6912 13068 7504 13096
rect 6912 13056 6918 13068
rect 7498 13056 7504 13068
rect 7556 13056 7562 13108
rect 7847 13040 7875 13127
rect 8602 13124 8608 13136
rect 8660 13124 8666 13176
rect 8786 13124 8792 13176
rect 8844 13164 8850 13176
rect 9246 13164 9252 13176
rect 8844 13136 9252 13164
rect 8844 13124 8850 13136
rect 9246 13124 9252 13136
rect 9304 13124 9310 13176
rect 9525 13167 9583 13173
rect 9525 13133 9537 13167
rect 9571 13164 9583 13167
rect 9798 13164 9804 13176
rect 9571 13136 9804 13164
rect 9571 13133 9583 13136
rect 9525 13127 9583 13133
rect 9157 13099 9215 13105
rect 9157 13065 9169 13099
rect 9203 13096 9215 13099
rect 9540 13096 9568 13127
rect 9798 13124 9804 13136
rect 9856 13124 9862 13176
rect 9982 13124 9988 13176
rect 10040 13164 10046 13176
rect 10629 13167 10687 13173
rect 10629 13164 10641 13167
rect 10040 13136 10641 13164
rect 10040 13124 10046 13136
rect 10629 13133 10641 13136
rect 10675 13133 10687 13167
rect 10629 13127 10687 13133
rect 9203 13068 9568 13096
rect 11012 13096 11040 13195
rect 13386 13192 13392 13204
rect 13444 13192 13450 13244
rect 14232 13241 14260 13272
rect 17250 13260 17256 13272
rect 17308 13260 17314 13312
rect 18630 13260 18636 13312
rect 18688 13300 18694 13312
rect 19274 13300 19280 13312
rect 18688 13272 19280 13300
rect 18688 13260 18694 13272
rect 19274 13260 19280 13272
rect 19332 13300 19338 13312
rect 19737 13303 19795 13309
rect 19737 13300 19749 13303
rect 19332 13272 19749 13300
rect 19332 13260 19338 13272
rect 19737 13269 19749 13272
rect 19783 13269 19795 13303
rect 19737 13263 19795 13269
rect 20381 13303 20439 13309
rect 20381 13269 20393 13303
rect 20427 13300 20439 13303
rect 21850 13300 21856 13312
rect 20427 13272 21856 13300
rect 20427 13269 20439 13272
rect 20381 13263 20439 13269
rect 21850 13260 21856 13272
rect 21908 13260 21914 13312
rect 23846 13300 23874 13340
rect 24061 13337 24073 13340
rect 24107 13337 24119 13371
rect 24061 13331 24119 13337
rect 24150 13328 24156 13380
rect 24208 13368 24214 13380
rect 24429 13371 24487 13377
rect 24429 13368 24441 13371
rect 24208 13340 24441 13368
rect 24208 13328 24214 13340
rect 24429 13337 24441 13340
rect 24475 13337 24487 13371
rect 24429 13331 24487 13337
rect 23616 13272 23874 13300
rect 14217 13235 14275 13241
rect 14217 13201 14229 13235
rect 14263 13201 14275 13235
rect 21206 13232 21212 13244
rect 21167 13204 21212 13232
rect 14217 13195 14275 13201
rect 21206 13192 21212 13204
rect 21264 13232 21270 13244
rect 22313 13235 22371 13241
rect 22313 13232 22325 13235
rect 21264 13204 22325 13232
rect 21264 13192 21270 13204
rect 22313 13201 22325 13204
rect 22359 13201 22371 13235
rect 22313 13195 22371 13201
rect 23049 13235 23107 13241
rect 23049 13201 23061 13235
rect 23095 13232 23107 13235
rect 23322 13232 23328 13244
rect 23095 13204 23328 13232
rect 23095 13201 23107 13204
rect 23049 13195 23107 13201
rect 23322 13192 23328 13204
rect 23380 13232 23386 13244
rect 23616 13241 23644 13272
rect 23601 13235 23659 13241
rect 23601 13232 23613 13235
rect 23380 13204 23613 13232
rect 23380 13192 23386 13204
rect 23601 13201 23613 13204
rect 23647 13201 23659 13235
rect 23601 13195 23659 13201
rect 23782 13192 23788 13244
rect 23840 13232 23846 13244
rect 23840 13204 25484 13232
rect 23840 13192 23846 13204
rect 11546 13124 11552 13176
rect 11604 13164 11610 13176
rect 11917 13167 11975 13173
rect 11917 13164 11929 13167
rect 11604 13136 11929 13164
rect 11604 13124 11610 13136
rect 11917 13133 11929 13136
rect 11963 13164 11975 13167
rect 12377 13167 12435 13173
rect 12377 13164 12389 13167
rect 11963 13136 12389 13164
rect 11963 13133 11975 13136
rect 11917 13127 11975 13133
rect 12377 13133 12389 13136
rect 12423 13133 12435 13167
rect 13294 13164 13300 13176
rect 12377 13127 12435 13133
rect 12484 13136 13300 13164
rect 11638 13096 11644 13108
rect 11012 13068 11644 13096
rect 9203 13065 9215 13068
rect 9157 13059 9215 13065
rect 11638 13056 11644 13068
rect 11696 13096 11702 13108
rect 11733 13099 11791 13105
rect 11733 13096 11745 13099
rect 11696 13068 11745 13096
rect 11696 13056 11702 13068
rect 11733 13065 11745 13068
rect 11779 13065 11791 13099
rect 11733 13059 11791 13065
rect 1334 13028 1340 13040
rect 1295 13000 1340 13028
rect 1334 12988 1340 13000
rect 1392 12988 1398 13040
rect 1521 13031 1579 13037
rect 1521 12997 1533 13031
rect 1567 13028 1579 13031
rect 1702 13028 1708 13040
rect 1567 13000 1708 13028
rect 1567 12997 1579 13000
rect 1521 12991 1579 12997
rect 1702 12988 1708 13000
rect 1760 12988 1766 13040
rect 3913 13031 3971 13037
rect 3913 12997 3925 13031
rect 3959 13028 3971 13031
rect 4002 13028 4008 13040
rect 3959 13000 4008 13028
rect 3959 12997 3971 13000
rect 3913 12991 3971 12997
rect 4002 12988 4008 13000
rect 4060 12988 4066 13040
rect 5382 12988 5388 13040
rect 5440 13028 5446 13040
rect 5750 13028 5756 13040
rect 5440 13000 5756 13028
rect 5440 12988 5446 13000
rect 5750 12988 5756 13000
rect 5808 13028 5814 13040
rect 6302 13028 6308 13040
rect 5808 13000 6308 13028
rect 5808 12988 5814 13000
rect 6302 12988 6308 13000
rect 6360 12988 6366 13040
rect 6397 13031 6455 13037
rect 6397 12997 6409 13031
rect 6443 13028 6455 13031
rect 6670 13028 6676 13040
rect 6443 13000 6676 13028
rect 6443 12997 6455 13000
rect 6397 12991 6455 12997
rect 6670 12988 6676 13000
rect 6728 12988 6734 13040
rect 7847 13000 7872 13040
rect 7866 12988 7872 13000
rect 7924 12988 7930 13040
rect 8878 13028 8884 13040
rect 8839 13000 8884 13028
rect 8878 12988 8884 13000
rect 8936 12988 8942 13040
rect 9706 13028 9712 13040
rect 9667 13000 9712 13028
rect 9706 12988 9712 13000
rect 9764 12988 9770 13040
rect 10350 13028 10356 13040
rect 10311 13000 10356 13028
rect 10350 12988 10356 13000
rect 10408 12988 10414 13040
rect 11748 13028 11776 13059
rect 12190 13056 12196 13108
rect 12248 13096 12254 13108
rect 12285 13099 12343 13105
rect 12285 13096 12297 13099
rect 12248 13068 12297 13096
rect 12248 13056 12254 13068
rect 12285 13065 12297 13068
rect 12331 13096 12343 13099
rect 12484 13096 12512 13136
rect 13294 13124 13300 13136
rect 13352 13124 13358 13176
rect 14125 13167 14183 13173
rect 14125 13133 14137 13167
rect 14171 13133 14183 13167
rect 14125 13127 14183 13133
rect 17621 13167 17679 13173
rect 17621 13133 17633 13167
rect 17667 13164 17679 13167
rect 17802 13164 17808 13176
rect 17667 13136 17808 13164
rect 17667 13133 17679 13136
rect 17621 13127 17679 13133
rect 13110 13096 13116 13108
rect 12331 13068 12512 13096
rect 13023 13068 13116 13096
rect 12331 13065 12343 13068
rect 12285 13059 12343 13065
rect 13110 13056 13116 13068
rect 13168 13096 13174 13108
rect 14140 13096 14168 13127
rect 17802 13124 17808 13136
rect 17860 13124 17866 13176
rect 19182 13124 19188 13176
rect 19240 13164 19246 13176
rect 19277 13167 19335 13173
rect 19277 13164 19289 13167
rect 19240 13136 19289 13164
rect 19240 13124 19246 13136
rect 19277 13133 19289 13136
rect 19323 13164 19335 13167
rect 20010 13164 20016 13176
rect 19323 13136 20016 13164
rect 19323 13133 19335 13136
rect 19277 13127 19335 13133
rect 20010 13124 20016 13136
rect 20068 13124 20074 13176
rect 20197 13167 20255 13173
rect 20197 13133 20209 13167
rect 20243 13164 20255 13167
rect 20378 13164 20384 13176
rect 20243 13136 20384 13164
rect 20243 13133 20255 13136
rect 20197 13127 20255 13133
rect 20378 13124 20384 13136
rect 20436 13164 20442 13176
rect 21301 13167 21359 13173
rect 21301 13164 21313 13167
rect 20436 13136 21313 13164
rect 20436 13124 20442 13136
rect 21301 13133 21313 13136
rect 21347 13133 21359 13167
rect 21666 13164 21672 13176
rect 21627 13136 21672 13164
rect 21301 13127 21359 13133
rect 13168 13068 14168 13096
rect 13168 13056 13174 13068
rect 17434 13056 17440 13108
rect 17492 13096 17498 13108
rect 17713 13099 17771 13105
rect 17713 13096 17725 13099
rect 17492 13068 17725 13096
rect 17492 13056 17498 13068
rect 17713 13065 17725 13068
rect 17759 13096 17771 13099
rect 17989 13099 18047 13105
rect 17989 13096 18001 13099
rect 17759 13068 18001 13096
rect 17759 13065 17771 13068
rect 17713 13059 17771 13065
rect 17989 13065 18001 13068
rect 18035 13065 18047 13099
rect 20654 13096 20660 13108
rect 20615 13068 20660 13096
rect 17989 13059 18047 13065
rect 20654 13056 20660 13068
rect 20712 13056 20718 13108
rect 21316 13096 21344 13127
rect 21666 13124 21672 13136
rect 21724 13124 21730 13176
rect 21850 13164 21856 13176
rect 21763 13136 21856 13164
rect 21850 13124 21856 13136
rect 21908 13164 21914 13176
rect 22218 13164 22224 13176
rect 21908 13136 22224 13164
rect 21908 13124 21914 13136
rect 22218 13124 22224 13136
rect 22276 13124 22282 13176
rect 23969 13167 24027 13173
rect 23969 13133 23981 13167
rect 24015 13164 24027 13167
rect 24150 13164 24156 13176
rect 24015 13136 24156 13164
rect 24015 13133 24027 13136
rect 23969 13127 24027 13133
rect 24150 13124 24156 13136
rect 24208 13124 24214 13176
rect 25456 13173 25484 13204
rect 25441 13167 25499 13173
rect 25441 13133 25453 13167
rect 25487 13164 25499 13167
rect 25487 13136 25760 13164
rect 25487 13133 25499 13136
rect 25441 13127 25499 13133
rect 21942 13096 21948 13108
rect 21316 13068 21948 13096
rect 21942 13056 21948 13068
rect 22000 13056 22006 13108
rect 23782 13096 23788 13108
rect 23743 13068 23788 13096
rect 23782 13056 23788 13068
rect 23840 13096 23846 13108
rect 24705 13099 24763 13105
rect 24705 13096 24717 13099
rect 23840 13068 24717 13096
rect 23840 13056 23846 13068
rect 24705 13065 24717 13068
rect 24751 13096 24763 13099
rect 25533 13099 25591 13105
rect 25533 13096 25545 13099
rect 24751 13068 25545 13096
rect 24751 13065 24763 13068
rect 24705 13059 24763 13065
rect 25533 13065 25545 13068
rect 25579 13096 25591 13099
rect 25625 13099 25683 13105
rect 25625 13096 25637 13099
rect 25579 13068 25637 13096
rect 25579 13065 25591 13068
rect 25533 13059 25591 13065
rect 25625 13065 25637 13068
rect 25671 13065 25683 13099
rect 25625 13059 25683 13065
rect 25732 13040 25760 13136
rect 12561 13031 12619 13037
rect 12561 13028 12573 13031
rect 11748 13000 12573 13028
rect 12561 12997 12573 13000
rect 12607 12997 12619 13031
rect 12561 12991 12619 12997
rect 20565 13031 20623 13037
rect 20565 12997 20577 13031
rect 20611 13028 20623 13031
rect 21666 13028 21672 13040
rect 20611 13000 21672 13028
rect 20611 12997 20623 13000
rect 20565 12991 20623 12997
rect 21666 12988 21672 13000
rect 21724 12988 21730 13040
rect 25714 12988 25720 13040
rect 25772 13028 25778 13040
rect 25809 13031 25867 13037
rect 25809 13028 25821 13031
rect 25772 13000 25821 13028
rect 25772 12988 25778 13000
rect 25809 12997 25821 13000
rect 25855 12997 25867 13031
rect 25809 12991 25867 12997
rect 400 12938 27264 12960
rect 400 12886 18870 12938
rect 18922 12886 18934 12938
rect 18986 12886 18998 12938
rect 19050 12886 19062 12938
rect 19114 12886 19126 12938
rect 19178 12886 27264 12938
rect 400 12864 27264 12886
rect 1242 12784 1248 12836
rect 1300 12824 1306 12836
rect 1889 12827 1947 12833
rect 1889 12824 1901 12827
rect 1300 12796 1901 12824
rect 1300 12784 1306 12796
rect 1889 12793 1901 12796
rect 1935 12793 1947 12827
rect 7314 12824 7320 12836
rect 1889 12787 1947 12793
rect 3928 12796 7320 12824
rect 2346 12716 2352 12768
rect 2404 12756 2410 12768
rect 3928 12756 3956 12796
rect 7314 12784 7320 12796
rect 7372 12784 7378 12836
rect 7682 12784 7688 12836
rect 7740 12824 7746 12836
rect 8053 12827 8111 12833
rect 8053 12824 8065 12827
rect 7740 12796 8065 12824
rect 7740 12784 7746 12796
rect 8053 12793 8065 12796
rect 8099 12793 8111 12827
rect 8053 12787 8111 12793
rect 8418 12784 8424 12836
rect 8476 12824 8482 12836
rect 9249 12827 9307 12833
rect 9249 12824 9261 12827
rect 8476 12796 9261 12824
rect 8476 12784 8482 12796
rect 9249 12793 9261 12796
rect 9295 12824 9307 12827
rect 9706 12824 9712 12836
rect 9295 12796 9712 12824
rect 9295 12793 9307 12796
rect 9249 12787 9307 12793
rect 9706 12784 9712 12796
rect 9764 12784 9770 12836
rect 12190 12824 12196 12836
rect 12151 12796 12196 12824
rect 12190 12784 12196 12796
rect 12248 12784 12254 12836
rect 13297 12827 13355 12833
rect 13297 12793 13309 12827
rect 13343 12824 13355 12827
rect 13386 12824 13392 12836
rect 13343 12796 13392 12824
rect 13343 12793 13355 12796
rect 13297 12787 13355 12793
rect 13386 12784 13392 12796
rect 13444 12784 13450 12836
rect 20470 12824 20476 12836
rect 20431 12796 20476 12824
rect 20470 12784 20476 12796
rect 20528 12784 20534 12836
rect 20654 12784 20660 12836
rect 20712 12824 20718 12836
rect 20841 12827 20899 12833
rect 20841 12824 20853 12827
rect 20712 12796 20853 12824
rect 20712 12784 20718 12796
rect 20841 12793 20853 12796
rect 20887 12793 20899 12827
rect 20841 12787 20899 12793
rect 2404 12728 3956 12756
rect 4189 12759 4247 12765
rect 2404 12716 2410 12728
rect 4189 12725 4201 12759
rect 4235 12756 4247 12759
rect 4922 12756 4928 12768
rect 4235 12728 4928 12756
rect 4235 12725 4247 12728
rect 4189 12719 4247 12725
rect 4922 12716 4928 12728
rect 4980 12716 4986 12768
rect 5845 12759 5903 12765
rect 5845 12725 5857 12759
rect 5891 12756 5903 12759
rect 6486 12756 6492 12768
rect 5891 12728 6492 12756
rect 5891 12725 5903 12728
rect 5845 12719 5903 12725
rect 6486 12716 6492 12728
rect 6544 12716 6550 12768
rect 7593 12759 7651 12765
rect 7593 12725 7605 12759
rect 7639 12756 7651 12759
rect 7958 12756 7964 12768
rect 7639 12728 7964 12756
rect 7639 12725 7651 12728
rect 7593 12719 7651 12725
rect 7958 12716 7964 12728
rect 8016 12716 8022 12768
rect 12208 12756 12236 12784
rect 17434 12756 17440 12768
rect 11472 12728 12236 12756
rect 17395 12728 17440 12756
rect 11472 12700 11500 12728
rect 17434 12716 17440 12728
rect 17492 12716 17498 12768
rect 1613 12691 1671 12697
rect 1613 12657 1625 12691
rect 1659 12688 1671 12691
rect 1702 12688 1708 12700
rect 1659 12660 1708 12688
rect 1659 12657 1671 12660
rect 1613 12651 1671 12657
rect 1702 12648 1708 12660
rect 1760 12648 1766 12700
rect 1797 12691 1855 12697
rect 1797 12657 1809 12691
rect 1843 12657 1855 12691
rect 1797 12651 1855 12657
rect 4373 12691 4431 12697
rect 4373 12657 4385 12691
rect 4419 12688 4431 12691
rect 4830 12688 4836 12700
rect 4419 12660 4836 12688
rect 4419 12657 4431 12660
rect 4373 12651 4431 12657
rect 1518 12580 1524 12632
rect 1576 12620 1582 12632
rect 1812 12620 1840 12651
rect 4830 12648 4836 12660
rect 4888 12648 4894 12700
rect 5937 12691 5995 12697
rect 5937 12657 5949 12691
rect 5983 12688 5995 12691
rect 7498 12688 7504 12700
rect 5983 12660 7504 12688
rect 5983 12657 5995 12660
rect 5937 12651 5995 12657
rect 7498 12648 7504 12660
rect 7556 12648 7562 12700
rect 7774 12688 7780 12700
rect 7735 12660 7780 12688
rect 7774 12648 7780 12660
rect 7832 12648 7838 12700
rect 9430 12648 9436 12700
rect 9488 12688 9494 12700
rect 10994 12688 11000 12700
rect 9488 12660 11000 12688
rect 9488 12648 9494 12660
rect 10994 12648 11000 12660
rect 11052 12648 11058 12700
rect 11454 12688 11460 12700
rect 11367 12660 11460 12688
rect 11454 12648 11460 12660
rect 11512 12648 11518 12700
rect 11825 12691 11883 12697
rect 11825 12657 11837 12691
rect 11871 12657 11883 12691
rect 11825 12651 11883 12657
rect 15229 12691 15287 12697
rect 15229 12657 15241 12691
rect 15275 12688 15287 12691
rect 15502 12688 15508 12700
rect 15275 12660 15508 12688
rect 15275 12657 15287 12660
rect 15229 12651 15287 12657
rect 4738 12620 4744 12632
rect 1576 12592 1840 12620
rect 4699 12592 4744 12620
rect 1576 12580 1582 12592
rect 4738 12580 4744 12592
rect 4796 12580 4802 12632
rect 5198 12580 5204 12632
rect 5256 12620 5262 12632
rect 6305 12623 6363 12629
rect 6305 12620 6317 12623
rect 5256 12592 6317 12620
rect 5256 12580 5262 12592
rect 6305 12589 6317 12592
rect 6351 12589 6363 12623
rect 6305 12583 6363 12589
rect 6394 12580 6400 12632
rect 6452 12620 6458 12632
rect 7866 12620 7872 12632
rect 6452 12592 7872 12620
rect 6452 12580 6458 12592
rect 7866 12580 7872 12592
rect 7924 12580 7930 12632
rect 8234 12620 8240 12632
rect 8195 12592 8240 12620
rect 8234 12580 8240 12592
rect 8292 12620 8298 12632
rect 8418 12620 8424 12632
rect 8292 12592 8424 12620
rect 8292 12580 8298 12592
rect 8418 12580 8424 12592
rect 8476 12620 8482 12632
rect 9522 12620 9528 12632
rect 8476 12592 9528 12620
rect 8476 12580 8482 12592
rect 9522 12580 9528 12592
rect 9580 12620 9586 12632
rect 9801 12623 9859 12629
rect 9801 12620 9813 12623
rect 9580 12592 9813 12620
rect 9580 12580 9586 12592
rect 9801 12589 9813 12592
rect 9847 12589 9859 12623
rect 9801 12583 9859 12589
rect 10810 12580 10816 12632
rect 10868 12620 10874 12632
rect 11840 12620 11868 12651
rect 15502 12648 15508 12660
rect 15560 12648 15566 12700
rect 17526 12648 17532 12700
rect 17584 12688 17590 12700
rect 17621 12691 17679 12697
rect 17621 12688 17633 12691
rect 17584 12660 17633 12688
rect 17584 12648 17590 12660
rect 17621 12657 17633 12660
rect 17667 12688 17679 12691
rect 18538 12688 18544 12700
rect 17667 12660 18544 12688
rect 17667 12657 17679 12660
rect 17621 12651 17679 12657
rect 18538 12648 18544 12660
rect 18596 12648 18602 12700
rect 20473 12691 20531 12697
rect 20473 12657 20485 12691
rect 20519 12688 20531 12691
rect 20672 12688 20700 12784
rect 23322 12716 23328 12768
rect 23380 12756 23386 12768
rect 24150 12756 24156 12768
rect 23380 12728 24156 12756
rect 23380 12716 23386 12728
rect 21666 12688 21672 12700
rect 20519 12660 20700 12688
rect 21627 12660 21672 12688
rect 20519 12657 20531 12660
rect 20473 12651 20531 12657
rect 21666 12648 21672 12660
rect 21724 12648 21730 12700
rect 21850 12688 21856 12700
rect 21811 12660 21856 12688
rect 21850 12648 21856 12660
rect 21908 12648 21914 12700
rect 22678 12648 22684 12700
rect 22736 12688 22742 12700
rect 23708 12697 23736 12728
rect 24150 12716 24156 12728
rect 24208 12716 24214 12768
rect 23417 12691 23475 12697
rect 23417 12688 23429 12691
rect 22736 12660 23429 12688
rect 22736 12648 22742 12660
rect 23417 12657 23429 12660
rect 23463 12657 23475 12691
rect 23417 12651 23475 12657
rect 23693 12691 23751 12697
rect 23693 12657 23705 12691
rect 23739 12657 23751 12691
rect 24058 12688 24064 12700
rect 24019 12660 24064 12688
rect 23693 12651 23751 12657
rect 24058 12648 24064 12660
rect 24116 12648 24122 12700
rect 10868 12592 11868 12620
rect 11917 12623 11975 12629
rect 10868 12580 10874 12592
rect 11917 12589 11929 12623
rect 11963 12589 11975 12623
rect 15410 12620 15416 12632
rect 15371 12592 15416 12620
rect 11917 12583 11975 12589
rect 3729 12555 3787 12561
rect 3729 12521 3741 12555
rect 3775 12552 3787 12555
rect 4002 12552 4008 12564
rect 3775 12524 4008 12552
rect 3775 12521 3787 12524
rect 3729 12515 3787 12521
rect 4002 12512 4008 12524
rect 4060 12512 4066 12564
rect 6213 12555 6271 12561
rect 6213 12552 6225 12555
rect 4526 12524 6225 12552
rect 4526 12496 4554 12524
rect 6213 12521 6225 12524
rect 6259 12552 6271 12555
rect 6765 12555 6823 12561
rect 6765 12552 6777 12555
rect 6259 12524 6777 12552
rect 6259 12521 6271 12524
rect 6213 12515 6271 12521
rect 6765 12521 6777 12524
rect 6811 12521 6823 12555
rect 7958 12552 7964 12564
rect 6765 12515 6823 12521
rect 7056 12524 7964 12552
rect 2254 12484 2260 12496
rect 2215 12456 2260 12484
rect 2254 12444 2260 12456
rect 2312 12444 2318 12496
rect 4094 12484 4100 12496
rect 4055 12456 4100 12484
rect 4094 12444 4100 12456
rect 4152 12444 4158 12496
rect 4462 12444 4468 12496
rect 4520 12456 4554 12496
rect 6102 12487 6160 12493
rect 4520 12444 4526 12456
rect 6102 12453 6114 12487
rect 6148 12484 6160 12487
rect 6302 12484 6308 12496
rect 6148 12456 6308 12484
rect 6148 12453 6160 12456
rect 6102 12447 6160 12453
rect 6302 12444 6308 12456
rect 6360 12444 6366 12496
rect 6486 12444 6492 12496
rect 6544 12484 6550 12496
rect 6581 12487 6639 12493
rect 6581 12484 6593 12487
rect 6544 12456 6593 12484
rect 6544 12444 6550 12456
rect 6581 12453 6593 12456
rect 6627 12484 6639 12487
rect 7056 12484 7084 12524
rect 7958 12512 7964 12524
rect 8016 12512 8022 12564
rect 11270 12512 11276 12564
rect 11328 12552 11334 12564
rect 11932 12552 11960 12583
rect 15410 12580 15416 12592
rect 15468 12580 15474 12632
rect 20749 12623 20807 12629
rect 20749 12589 20761 12623
rect 20795 12620 20807 12623
rect 21942 12620 21948 12632
rect 20795 12592 21948 12620
rect 20795 12589 20807 12592
rect 20749 12583 20807 12589
rect 21942 12580 21948 12592
rect 22000 12580 22006 12632
rect 22770 12580 22776 12632
rect 22828 12620 22834 12632
rect 23782 12620 23788 12632
rect 22828 12592 23788 12620
rect 22828 12580 22834 12592
rect 23782 12580 23788 12592
rect 23840 12620 23846 12632
rect 23969 12623 24027 12629
rect 23969 12620 23981 12623
rect 23840 12592 23981 12620
rect 23840 12580 23846 12592
rect 23969 12589 23981 12592
rect 24015 12589 24027 12623
rect 23969 12583 24027 12589
rect 23506 12552 23512 12564
rect 11328 12524 11960 12552
rect 23467 12524 23512 12552
rect 11328 12512 11334 12524
rect 23506 12512 23512 12524
rect 23564 12512 23570 12564
rect 6627 12456 7084 12484
rect 6627 12453 6639 12456
rect 6581 12447 6639 12453
rect 7222 12444 7228 12496
rect 7280 12484 7286 12496
rect 7409 12487 7467 12493
rect 7409 12484 7421 12487
rect 7280 12456 7421 12484
rect 7280 12444 7286 12456
rect 7409 12453 7421 12456
rect 7455 12484 7467 12487
rect 8050 12484 8056 12496
rect 7455 12456 8056 12484
rect 7455 12453 7467 12456
rect 7409 12447 7467 12453
rect 8050 12444 8056 12456
rect 8108 12484 8114 12496
rect 9522 12484 9528 12496
rect 8108 12456 9528 12484
rect 8108 12444 8114 12456
rect 9522 12444 9528 12456
rect 9580 12444 9586 12496
rect 14306 12484 14312 12496
rect 14267 12456 14312 12484
rect 14306 12444 14312 12456
rect 14364 12484 14370 12496
rect 15870 12484 15876 12496
rect 14364 12456 15876 12484
rect 14364 12444 14370 12456
rect 15870 12444 15876 12456
rect 15928 12444 15934 12496
rect 17710 12484 17716 12496
rect 17671 12456 17716 12484
rect 17710 12444 17716 12456
rect 17768 12444 17774 12496
rect 400 12394 27264 12416
rect 400 12342 3510 12394
rect 3562 12342 3574 12394
rect 3626 12342 3638 12394
rect 3690 12342 3702 12394
rect 3754 12342 3766 12394
rect 3818 12342 27264 12394
rect 400 12320 27264 12342
rect 1242 12280 1248 12292
rect 1203 12252 1248 12280
rect 1242 12240 1248 12252
rect 1300 12240 1306 12292
rect 1702 12240 1708 12292
rect 1760 12280 1766 12292
rect 1889 12283 1947 12289
rect 1889 12280 1901 12283
rect 1760 12252 1901 12280
rect 1760 12240 1766 12252
rect 1889 12249 1901 12252
rect 1935 12280 1947 12283
rect 1935 12252 4784 12280
rect 1935 12249 1947 12252
rect 1889 12243 1947 12249
rect 4756 12224 4784 12252
rect 5198 12240 5204 12292
rect 5256 12280 5262 12292
rect 5845 12283 5903 12289
rect 5845 12280 5857 12283
rect 5256 12252 5857 12280
rect 5256 12240 5262 12252
rect 5845 12249 5857 12252
rect 5891 12249 5903 12283
rect 6394 12280 6400 12292
rect 6355 12252 6400 12280
rect 5845 12243 5903 12249
rect 6394 12240 6400 12252
rect 6452 12240 6458 12292
rect 6578 12280 6584 12292
rect 6539 12252 6584 12280
rect 6578 12240 6584 12252
rect 6636 12280 6642 12292
rect 7133 12283 7191 12289
rect 7133 12280 7145 12283
rect 6636 12252 7145 12280
rect 6636 12240 6642 12252
rect 7133 12249 7145 12252
rect 7179 12249 7191 12283
rect 7498 12280 7504 12292
rect 7411 12252 7504 12280
rect 7133 12243 7191 12249
rect 7498 12240 7504 12252
rect 7556 12280 7562 12292
rect 8142 12280 8148 12292
rect 7556 12252 8148 12280
rect 7556 12240 7562 12252
rect 8142 12240 8148 12252
rect 8200 12240 8206 12292
rect 8234 12240 8240 12292
rect 8292 12280 8298 12292
rect 9982 12280 9988 12292
rect 8292 12252 9988 12280
rect 8292 12240 8298 12252
rect 9982 12240 9988 12252
rect 10040 12240 10046 12292
rect 11454 12280 11460 12292
rect 11415 12252 11460 12280
rect 11454 12240 11460 12252
rect 11512 12240 11518 12292
rect 17434 12240 17440 12292
rect 17492 12280 17498 12292
rect 17621 12283 17679 12289
rect 17621 12280 17633 12283
rect 17492 12252 17633 12280
rect 17492 12240 17498 12252
rect 17621 12249 17633 12252
rect 17667 12249 17679 12283
rect 17621 12243 17679 12249
rect 17710 12240 17716 12292
rect 17768 12280 17774 12292
rect 17805 12283 17863 12289
rect 17805 12280 17817 12283
rect 17768 12252 17817 12280
rect 17768 12240 17774 12252
rect 17805 12249 17817 12252
rect 17851 12249 17863 12283
rect 17805 12243 17863 12249
rect 20289 12283 20347 12289
rect 20289 12249 20301 12283
rect 20335 12280 20347 12283
rect 20654 12280 20660 12292
rect 20335 12252 20660 12280
rect 20335 12249 20347 12252
rect 20289 12243 20347 12249
rect 20654 12240 20660 12252
rect 20712 12240 20718 12292
rect 21853 12283 21911 12289
rect 21853 12249 21865 12283
rect 21899 12280 21911 12283
rect 21942 12280 21948 12292
rect 21899 12252 21948 12280
rect 21899 12249 21911 12252
rect 21853 12243 21911 12249
rect 21942 12240 21948 12252
rect 22000 12240 22006 12292
rect 22770 12280 22776 12292
rect 22731 12252 22776 12280
rect 22770 12240 22776 12252
rect 22828 12240 22834 12292
rect 23322 12280 23328 12292
rect 23283 12252 23328 12280
rect 23322 12240 23328 12252
rect 23380 12240 23386 12292
rect 23506 12280 23512 12292
rect 23467 12252 23512 12280
rect 23506 12240 23512 12252
rect 23564 12240 23570 12292
rect 1521 12215 1579 12221
rect 1521 12181 1533 12215
rect 1567 12212 1579 12215
rect 2349 12215 2407 12221
rect 2349 12212 2361 12215
rect 1567 12184 2361 12212
rect 1567 12181 1579 12184
rect 1521 12175 1579 12181
rect 2349 12181 2361 12184
rect 2395 12212 2407 12215
rect 2395 12184 3588 12212
rect 2395 12181 2407 12184
rect 2349 12175 2407 12181
rect 2254 12153 2260 12156
rect 2220 12147 2260 12153
rect 2220 12113 2232 12147
rect 2220 12107 2260 12113
rect 2254 12104 2260 12107
rect 2312 12104 2318 12156
rect 2441 12147 2499 12153
rect 2441 12113 2453 12147
rect 2487 12144 2499 12147
rect 2714 12144 2720 12156
rect 2487 12116 2720 12144
rect 2487 12113 2499 12116
rect 2441 12107 2499 12113
rect 2714 12104 2720 12116
rect 2772 12104 2778 12156
rect 3358 12104 3364 12156
rect 3416 12144 3422 12156
rect 3453 12147 3511 12153
rect 3453 12144 3465 12147
rect 3416 12116 3465 12144
rect 3416 12104 3422 12116
rect 3453 12113 3465 12116
rect 3499 12113 3511 12147
rect 3560 12144 3588 12184
rect 4462 12172 4468 12224
rect 4520 12212 4526 12224
rect 4557 12215 4615 12221
rect 4557 12212 4569 12215
rect 4520 12184 4569 12212
rect 4520 12172 4526 12184
rect 4557 12181 4569 12184
rect 4603 12212 4615 12215
rect 4646 12212 4652 12224
rect 4603 12184 4652 12212
rect 4603 12181 4615 12184
rect 4557 12175 4615 12181
rect 4646 12172 4652 12184
rect 4704 12172 4710 12224
rect 4738 12172 4744 12224
rect 4796 12212 4802 12224
rect 5109 12215 5167 12221
rect 5109 12212 5121 12215
rect 4796 12184 5121 12212
rect 4796 12172 4802 12184
rect 5109 12181 5121 12184
rect 5155 12212 5167 12215
rect 5569 12215 5627 12221
rect 5569 12212 5581 12215
rect 5155 12184 5581 12212
rect 5155 12181 5167 12184
rect 5109 12175 5167 12181
rect 5569 12181 5581 12184
rect 5615 12212 5627 12215
rect 6259 12215 6317 12221
rect 6259 12212 6271 12215
rect 5615 12184 6271 12212
rect 5615 12181 5627 12184
rect 5569 12175 5627 12181
rect 6259 12181 6271 12184
rect 6305 12181 6317 12215
rect 6259 12175 6317 12181
rect 3560 12116 3680 12144
rect 3453 12107 3511 12113
rect 2073 12079 2131 12085
rect 2073 12045 2085 12079
rect 2119 12076 2131 12079
rect 2901 12079 2959 12085
rect 2901 12076 2913 12079
rect 2119 12048 2913 12076
rect 2119 12045 2131 12048
rect 2073 12039 2131 12045
rect 2901 12045 2913 12048
rect 2947 12076 2959 12079
rect 2990 12076 2996 12088
rect 2947 12048 2996 12076
rect 2947 12045 2959 12048
rect 2901 12039 2959 12045
rect 2990 12036 2996 12048
rect 3048 12036 3054 12088
rect 3652 12076 3680 12116
rect 3726 12104 3732 12156
rect 3784 12144 3790 12156
rect 4373 12147 4431 12153
rect 4373 12144 4385 12147
rect 3784 12116 4385 12144
rect 3784 12104 3790 12116
rect 4373 12113 4385 12116
rect 4419 12113 4431 12147
rect 4373 12107 4431 12113
rect 5658 12104 5664 12156
rect 5716 12144 5722 12156
rect 5753 12147 5811 12153
rect 5753 12144 5765 12147
rect 5716 12116 5765 12144
rect 5716 12104 5722 12116
rect 5753 12113 5765 12116
rect 5799 12144 5811 12147
rect 6412 12144 6440 12240
rect 7041 12215 7099 12221
rect 7041 12212 7053 12215
rect 6504 12184 7053 12212
rect 6504 12153 6532 12184
rect 7041 12181 7053 12184
rect 7087 12212 7099 12215
rect 7774 12212 7780 12224
rect 7087 12184 7780 12212
rect 7087 12181 7099 12184
rect 7041 12175 7099 12181
rect 7774 12172 7780 12184
rect 7832 12172 7838 12224
rect 10994 12172 11000 12224
rect 11052 12212 11058 12224
rect 11733 12215 11791 12221
rect 11733 12212 11745 12215
rect 11052 12184 11745 12212
rect 11052 12172 11058 12184
rect 11733 12181 11745 12184
rect 11779 12212 11791 12215
rect 12282 12212 12288 12224
rect 11779 12184 12288 12212
rect 11779 12181 11791 12184
rect 11733 12175 11791 12181
rect 12282 12172 12288 12184
rect 12340 12172 12346 12224
rect 17526 12212 17532 12224
rect 17487 12184 17532 12212
rect 17526 12172 17532 12184
rect 17584 12172 17590 12224
rect 20470 12212 20476 12224
rect 20431 12184 20476 12212
rect 20470 12172 20476 12184
rect 20528 12172 20534 12224
rect 22589 12215 22647 12221
rect 22589 12181 22601 12215
rect 22635 12212 22647 12215
rect 22678 12212 22684 12224
rect 22635 12184 22684 12212
rect 22635 12181 22647 12184
rect 22589 12175 22647 12181
rect 22678 12172 22684 12184
rect 22736 12172 22742 12224
rect 5799 12116 6440 12144
rect 6489 12147 6547 12153
rect 5799 12113 5811 12116
rect 5753 12107 5811 12113
rect 6489 12113 6501 12147
rect 6535 12113 6547 12147
rect 14306 12144 14312 12156
rect 14267 12116 14312 12144
rect 6489 12107 6547 12113
rect 14306 12104 14312 12116
rect 14364 12104 14370 12156
rect 21669 12147 21727 12153
rect 21669 12113 21681 12147
rect 21715 12144 21727 12147
rect 21850 12144 21856 12156
rect 21715 12116 21856 12144
rect 21715 12113 21727 12116
rect 21669 12107 21727 12113
rect 21850 12104 21856 12116
rect 21908 12104 21914 12156
rect 23141 12147 23199 12153
rect 23141 12113 23153 12147
rect 23187 12144 23199 12147
rect 23524 12144 23552 12240
rect 23969 12147 24027 12153
rect 23969 12144 23981 12147
rect 23187 12116 23981 12144
rect 23187 12113 23199 12116
rect 23141 12107 23199 12113
rect 23969 12113 23981 12116
rect 24015 12113 24027 12147
rect 23969 12107 24027 12113
rect 4278 12076 4284 12088
rect 3652 12048 4284 12076
rect 4278 12036 4284 12048
rect 4336 12076 4342 12088
rect 6302 12076 6308 12088
rect 4336 12048 6308 12076
rect 4336 12036 4342 12048
rect 6302 12036 6308 12048
rect 6360 12076 6366 12088
rect 7317 12079 7375 12085
rect 7317 12076 7329 12079
rect 6360 12048 7329 12076
rect 6360 12036 6366 12048
rect 7317 12045 7329 12048
rect 7363 12045 7375 12079
rect 7317 12039 7375 12045
rect 7498 12036 7504 12088
rect 7556 12076 7562 12088
rect 7961 12079 8019 12085
rect 7961 12076 7973 12079
rect 7556 12048 7973 12076
rect 7556 12036 7562 12048
rect 7961 12045 7973 12048
rect 8007 12076 8019 12079
rect 11454 12076 11460 12088
rect 8007 12048 11460 12076
rect 8007 12045 8019 12048
rect 7961 12039 8019 12045
rect 3361 12011 3419 12017
rect 3361 11977 3373 12011
rect 3407 12008 3419 12011
rect 4002 12008 4008 12020
rect 3407 11980 3588 12008
rect 3915 11980 4008 12008
rect 3407 11977 3419 11980
rect 3361 11971 3419 11977
rect 1518 11900 1524 11952
rect 1576 11940 1582 11952
rect 1613 11943 1671 11949
rect 1613 11940 1625 11943
rect 1576 11912 1625 11940
rect 1576 11900 1582 11912
rect 1613 11909 1625 11912
rect 1659 11909 1671 11943
rect 1613 11903 1671 11909
rect 2162 11900 2168 11952
rect 2220 11940 2226 11952
rect 2717 11943 2775 11949
rect 2717 11940 2729 11943
rect 2220 11912 2729 11940
rect 2220 11900 2226 11912
rect 2717 11909 2729 11912
rect 2763 11909 2775 11943
rect 3560 11940 3588 11980
rect 4002 11968 4008 11980
rect 4060 12008 4066 12020
rect 4554 12008 4560 12020
rect 4060 11980 4560 12008
rect 4060 11968 4066 11980
rect 4554 11968 4560 11980
rect 4612 11968 4618 12020
rect 5385 12011 5443 12017
rect 4664 11980 5336 12008
rect 4664 11952 4692 11980
rect 3818 11940 3824 11952
rect 3560 11912 3824 11940
rect 2717 11903 2775 11909
rect 3818 11900 3824 11912
rect 3876 11900 3882 11952
rect 3913 11943 3971 11949
rect 3913 11909 3925 11943
rect 3959 11940 3971 11943
rect 4462 11940 4468 11952
rect 3959 11912 4468 11940
rect 3959 11909 3971 11912
rect 3913 11903 3971 11909
rect 4462 11900 4468 11912
rect 4520 11900 4526 11952
rect 4646 11940 4652 11952
rect 4607 11912 4652 11940
rect 4646 11900 4652 11912
rect 4704 11900 4710 11952
rect 4922 11940 4928 11952
rect 4883 11912 4928 11940
rect 4922 11900 4928 11912
rect 4980 11900 4986 11952
rect 5308 11940 5336 11980
rect 5385 11977 5397 12011
rect 5431 12008 5443 12011
rect 5934 12008 5940 12020
rect 5431 11980 5940 12008
rect 5431 11977 5443 11980
rect 5385 11971 5443 11977
rect 5934 11968 5940 11980
rect 5992 12008 5998 12020
rect 6121 12011 6179 12017
rect 6121 12008 6133 12011
rect 5992 11980 6133 12008
rect 5992 11968 5998 11980
rect 6121 11977 6133 11980
rect 6167 11977 6179 12011
rect 6121 11971 6179 11977
rect 7130 11968 7136 12020
rect 7188 12008 7194 12020
rect 8053 12011 8111 12017
rect 8053 12008 8065 12011
rect 7188 11980 8065 12008
rect 7188 11968 7194 11980
rect 8053 11977 8065 11980
rect 8099 11977 8111 12011
rect 8234 12008 8240 12020
rect 8195 11980 8240 12008
rect 8053 11971 8111 11977
rect 8234 11968 8240 11980
rect 8292 11968 8298 12020
rect 8436 12017 8464 12048
rect 11454 12036 11460 12048
rect 11512 12036 11518 12088
rect 23690 12076 23696 12088
rect 23651 12048 23696 12076
rect 23690 12036 23696 12048
rect 23748 12036 23754 12088
rect 8421 12011 8479 12017
rect 8421 11977 8433 12011
rect 8467 11977 8479 12011
rect 8786 12008 8792 12020
rect 8747 11980 8792 12008
rect 8421 11971 8479 11977
rect 8786 11968 8792 11980
rect 8844 11968 8850 12020
rect 14217 12011 14275 12017
rect 14217 11977 14229 12011
rect 14263 12008 14275 12011
rect 14490 12008 14496 12020
rect 14263 11980 14496 12008
rect 14263 11977 14275 11980
rect 14217 11971 14275 11977
rect 14490 11968 14496 11980
rect 14548 12008 14554 12020
rect 14585 12011 14643 12017
rect 14585 12008 14597 12011
rect 14548 11980 14597 12008
rect 14548 11968 14554 11980
rect 14585 11977 14597 11980
rect 14631 11977 14643 12011
rect 14585 11971 14643 11977
rect 15318 11968 15324 12020
rect 15376 11968 15382 12020
rect 16330 12008 16336 12020
rect 16291 11980 16336 12008
rect 16330 11968 16336 11980
rect 16388 11968 16394 12020
rect 21485 12011 21543 12017
rect 21485 11977 21497 12011
rect 21531 12008 21543 12011
rect 21666 12008 21672 12020
rect 21531 11980 21672 12008
rect 21531 11977 21543 11980
rect 21485 11971 21543 11977
rect 21666 11968 21672 11980
rect 21724 12008 21730 12020
rect 21724 11980 23874 12008
rect 21724 11968 21730 11980
rect 6210 11940 6216 11952
rect 5308 11912 6216 11940
rect 6210 11900 6216 11912
rect 6268 11940 6274 11952
rect 7682 11940 7688 11952
rect 6268 11912 7688 11940
rect 6268 11900 6274 11912
rect 7682 11900 7688 11912
rect 7740 11900 7746 11952
rect 8326 11900 8332 11952
rect 8384 11940 8390 11952
rect 8881 11943 8939 11949
rect 8881 11940 8893 11943
rect 8384 11912 8893 11940
rect 8384 11900 8390 11912
rect 8881 11909 8893 11912
rect 8927 11940 8939 11943
rect 10810 11940 10816 11952
rect 8927 11912 10816 11940
rect 8927 11909 8939 11912
rect 8881 11903 8939 11909
rect 10810 11900 10816 11912
rect 10868 11940 10874 11952
rect 10997 11943 11055 11949
rect 10997 11940 11009 11943
rect 10868 11912 11009 11940
rect 10868 11900 10874 11912
rect 10997 11909 11009 11912
rect 11043 11909 11055 11943
rect 11270 11940 11276 11952
rect 11231 11912 11276 11940
rect 10997 11903 11055 11909
rect 11270 11900 11276 11912
rect 11328 11900 11334 11952
rect 14033 11943 14091 11949
rect 14033 11909 14045 11943
rect 14079 11940 14091 11943
rect 15336 11940 15364 11968
rect 14079 11912 15364 11940
rect 23846 11940 23874 11980
rect 24702 11968 24708 12020
rect 24760 11968 24766 12020
rect 25714 12008 25720 12020
rect 25675 11980 25720 12008
rect 25714 11968 25720 11980
rect 25772 11968 25778 12020
rect 24610 11940 24616 11952
rect 23846 11912 24616 11940
rect 14079 11909 14091 11912
rect 14033 11903 14091 11909
rect 24610 11900 24616 11912
rect 24668 11900 24674 11952
rect 400 11850 27264 11872
rect 400 11798 18870 11850
rect 18922 11798 18934 11850
rect 18986 11798 18998 11850
rect 19050 11798 19062 11850
rect 19114 11798 19126 11850
rect 19178 11798 27264 11850
rect 400 11776 27264 11798
rect 2257 11739 2315 11745
rect 2257 11705 2269 11739
rect 2303 11736 2315 11739
rect 2714 11736 2720 11748
rect 2303 11708 2720 11736
rect 2303 11705 2315 11708
rect 2257 11699 2315 11705
rect 2714 11696 2720 11708
rect 2772 11696 2778 11748
rect 3910 11736 3916 11748
rect 3871 11708 3916 11736
rect 3910 11696 3916 11708
rect 3968 11696 3974 11748
rect 4462 11736 4468 11748
rect 4423 11708 4468 11736
rect 4462 11696 4468 11708
rect 4520 11696 4526 11748
rect 7498 11736 7504 11748
rect 4664 11708 7504 11736
rect 1521 11671 1579 11677
rect 1521 11637 1533 11671
rect 1567 11668 1579 11671
rect 1794 11668 1800 11680
rect 1567 11640 1800 11668
rect 1567 11637 1579 11640
rect 1521 11631 1579 11637
rect 1794 11628 1800 11640
rect 1852 11668 1858 11680
rect 3637 11671 3695 11677
rect 3637 11668 3649 11671
rect 1852 11640 3649 11668
rect 1852 11628 1858 11640
rect 3637 11637 3649 11640
rect 3683 11668 3695 11671
rect 3726 11668 3732 11680
rect 3683 11640 3732 11668
rect 3683 11637 3695 11640
rect 3637 11631 3695 11637
rect 3726 11628 3732 11640
rect 3784 11628 3790 11680
rect 4373 11671 4431 11677
rect 4373 11668 4385 11671
rect 4296 11640 4385 11668
rect 1610 11560 1616 11612
rect 1668 11600 1674 11612
rect 1705 11603 1763 11609
rect 1705 11600 1717 11603
rect 1668 11572 1717 11600
rect 1668 11560 1674 11572
rect 1705 11569 1717 11572
rect 1751 11569 1763 11603
rect 1705 11563 1763 11569
rect 3818 11560 3824 11612
rect 3876 11600 3882 11612
rect 4296 11600 4324 11640
rect 4373 11637 4385 11640
rect 4419 11637 4431 11671
rect 4373 11631 4431 11637
rect 4554 11609 4560 11612
rect 3876 11572 4324 11600
rect 3876 11560 3882 11572
rect 4189 11535 4247 11541
rect 4189 11501 4201 11535
rect 4235 11501 4247 11535
rect 4296 11532 4324 11572
rect 4541 11603 4560 11609
rect 4541 11569 4553 11603
rect 4612 11600 4618 11612
rect 4664 11600 4692 11708
rect 7498 11696 7504 11708
rect 7556 11696 7562 11748
rect 7682 11696 7688 11748
rect 7740 11736 7746 11748
rect 8786 11736 8792 11748
rect 7740 11708 8792 11736
rect 7740 11696 7746 11708
rect 8786 11696 8792 11708
rect 8844 11696 8850 11748
rect 9433 11739 9491 11745
rect 9433 11705 9445 11739
rect 9479 11736 9491 11739
rect 10166 11736 10172 11748
rect 9479 11708 10172 11736
rect 9479 11705 9491 11708
rect 9433 11699 9491 11705
rect 10166 11696 10172 11708
rect 10224 11696 10230 11748
rect 10810 11736 10816 11748
rect 10771 11708 10816 11736
rect 10810 11696 10816 11708
rect 10868 11696 10874 11748
rect 15410 11736 15416 11748
rect 15371 11708 15416 11736
rect 15410 11696 15416 11708
rect 15468 11696 15474 11748
rect 23141 11739 23199 11745
rect 23141 11705 23153 11739
rect 23187 11736 23199 11739
rect 23322 11736 23328 11748
rect 23187 11708 23328 11736
rect 23187 11705 23199 11708
rect 23141 11699 23199 11705
rect 23322 11696 23328 11708
rect 23380 11736 23386 11748
rect 24058 11736 24064 11748
rect 23380 11708 24064 11736
rect 23380 11696 23386 11708
rect 24058 11696 24064 11708
rect 24116 11696 24122 11748
rect 24153 11739 24211 11745
rect 24153 11705 24165 11739
rect 24199 11736 24211 11739
rect 25714 11736 25720 11748
rect 24199 11708 25720 11736
rect 24199 11705 24211 11708
rect 24153 11699 24211 11705
rect 25714 11696 25720 11708
rect 25772 11696 25778 11748
rect 5934 11668 5940 11680
rect 5895 11640 5940 11668
rect 5934 11628 5940 11640
rect 5992 11628 5998 11680
rect 6854 11628 6860 11680
rect 6912 11668 6918 11680
rect 7317 11671 7375 11677
rect 7317 11668 7329 11671
rect 6912 11640 7329 11668
rect 6912 11628 6918 11640
rect 7317 11637 7329 11640
rect 7363 11668 7375 11671
rect 7866 11668 7872 11680
rect 7363 11640 7872 11668
rect 7363 11637 7375 11640
rect 7317 11631 7375 11637
rect 7866 11628 7872 11640
rect 7924 11628 7930 11680
rect 9522 11668 9528 11680
rect 9483 11640 9528 11668
rect 9522 11628 9528 11640
rect 9580 11628 9586 11680
rect 13294 11628 13300 11680
rect 13352 11668 13358 11680
rect 14401 11671 14459 11677
rect 14401 11668 14413 11671
rect 13352 11640 14413 11668
rect 13352 11628 13358 11640
rect 14401 11637 14413 11640
rect 14447 11668 14459 11671
rect 15594 11668 15600 11680
rect 14447 11640 15600 11668
rect 14447 11637 14459 11640
rect 14401 11631 14459 11637
rect 15594 11628 15600 11640
rect 15652 11668 15658 11680
rect 16330 11668 16336 11680
rect 15652 11640 16336 11668
rect 15652 11628 15658 11640
rect 16330 11628 16336 11640
rect 16388 11628 16394 11680
rect 23785 11671 23843 11677
rect 23785 11637 23797 11671
rect 23831 11668 23843 11671
rect 24702 11668 24708 11680
rect 23831 11640 24708 11668
rect 23831 11637 23843 11640
rect 23785 11631 23843 11637
rect 24702 11628 24708 11640
rect 24760 11628 24766 11680
rect 5750 11600 5756 11612
rect 4612 11572 4705 11600
rect 4756 11572 5756 11600
rect 4541 11563 4560 11569
rect 4554 11560 4560 11563
rect 4612 11560 4618 11572
rect 4756 11544 4784 11572
rect 5750 11560 5756 11572
rect 5808 11560 5814 11612
rect 6394 11560 6400 11612
rect 6452 11600 6458 11612
rect 6765 11603 6823 11609
rect 6765 11600 6777 11603
rect 6452 11572 6777 11600
rect 6452 11560 6458 11572
rect 6765 11569 6777 11572
rect 6811 11600 6823 11603
rect 7406 11600 7412 11612
rect 6811 11572 7412 11600
rect 6811 11569 6823 11572
rect 6765 11563 6823 11569
rect 7406 11560 7412 11572
rect 7464 11560 7470 11612
rect 9338 11600 9344 11612
rect 9299 11572 9344 11600
rect 9338 11560 9344 11572
rect 9396 11560 9402 11612
rect 10166 11560 10172 11612
rect 10224 11600 10230 11612
rect 10721 11603 10779 11609
rect 10721 11600 10733 11603
rect 10224 11572 10733 11600
rect 10224 11560 10230 11572
rect 10721 11569 10733 11572
rect 10767 11569 10779 11603
rect 12834 11600 12840 11612
rect 12795 11572 12840 11600
rect 10721 11563 10779 11569
rect 12834 11560 12840 11572
rect 12892 11560 12898 11612
rect 15321 11603 15379 11609
rect 15321 11569 15333 11603
rect 15367 11600 15379 11603
rect 15502 11600 15508 11612
rect 15367 11572 15508 11600
rect 15367 11569 15379 11572
rect 15321 11563 15379 11569
rect 15502 11560 15508 11572
rect 15560 11560 15566 11612
rect 23690 11560 23696 11612
rect 23748 11600 23754 11612
rect 23877 11603 23935 11609
rect 23877 11600 23889 11603
rect 23748 11572 23889 11600
rect 23748 11560 23754 11572
rect 23877 11569 23889 11572
rect 23923 11569 23935 11603
rect 24426 11600 24432 11612
rect 24387 11572 24432 11600
rect 23877 11563 23935 11569
rect 24426 11560 24432 11572
rect 24484 11560 24490 11612
rect 4738 11532 4744 11544
rect 4296 11504 4744 11532
rect 4189 11495 4247 11501
rect 2254 11424 2260 11476
rect 2312 11464 2318 11476
rect 4204 11464 4232 11495
rect 4738 11492 4744 11504
rect 4796 11492 4802 11544
rect 4922 11532 4928 11544
rect 4883 11504 4928 11532
rect 4922 11492 4928 11504
rect 4980 11492 4986 11544
rect 6489 11535 6547 11541
rect 6489 11501 6501 11535
rect 6535 11532 6547 11535
rect 6670 11532 6676 11544
rect 6535 11504 6676 11532
rect 6535 11501 6547 11504
rect 6489 11495 6547 11501
rect 6670 11492 6676 11504
rect 6728 11492 6734 11544
rect 6949 11535 7007 11541
rect 6949 11501 6961 11535
rect 6995 11501 7007 11535
rect 6949 11495 7007 11501
rect 5198 11464 5204 11476
rect 2312 11436 3956 11464
rect 4204 11436 5204 11464
rect 2312 11424 2318 11436
rect 1518 11356 1524 11408
rect 1576 11396 1582 11408
rect 1797 11399 1855 11405
rect 1797 11396 1809 11399
rect 1576 11368 1809 11396
rect 1576 11356 1582 11368
rect 1797 11365 1809 11368
rect 1843 11365 1855 11399
rect 1797 11359 1855 11365
rect 2162 11356 2168 11408
rect 2220 11396 2226 11408
rect 2349 11399 2407 11405
rect 2349 11396 2361 11399
rect 2220 11368 2361 11396
rect 2220 11356 2226 11368
rect 2349 11365 2361 11368
rect 2395 11365 2407 11399
rect 3928 11396 3956 11436
rect 5198 11424 5204 11436
rect 5256 11424 5262 11476
rect 5566 11424 5572 11476
rect 5624 11464 5630 11476
rect 6762 11464 6768 11476
rect 5624 11436 6768 11464
rect 5624 11424 5630 11436
rect 6762 11424 6768 11436
rect 6820 11464 6826 11476
rect 6964 11464 6992 11495
rect 8602 11492 8608 11544
rect 8660 11532 8666 11544
rect 9157 11535 9215 11541
rect 9157 11532 9169 11535
rect 8660 11504 9169 11532
rect 8660 11492 8666 11504
rect 9157 11501 9169 11504
rect 9203 11501 9215 11535
rect 9157 11495 9215 11501
rect 9706 11492 9712 11544
rect 9764 11532 9770 11544
rect 9893 11535 9951 11541
rect 9893 11532 9905 11535
rect 9764 11504 9905 11532
rect 9764 11492 9770 11504
rect 9893 11501 9905 11504
rect 9939 11501 9951 11535
rect 9893 11495 9951 11501
rect 6820 11436 6992 11464
rect 6820 11424 6826 11436
rect 12926 11424 12932 11476
rect 12984 11464 12990 11476
rect 14585 11467 14643 11473
rect 14585 11464 14597 11467
rect 12984 11436 14597 11464
rect 12984 11424 12990 11436
rect 14585 11433 14597 11436
rect 14631 11464 14643 11467
rect 14858 11464 14864 11476
rect 14631 11436 14864 11464
rect 14631 11433 14643 11436
rect 14585 11427 14643 11433
rect 14858 11424 14864 11436
rect 14916 11424 14922 11476
rect 4370 11396 4376 11408
rect 3928 11368 4376 11396
rect 2349 11359 2407 11365
rect 4370 11356 4376 11368
rect 4428 11356 4434 11408
rect 6302 11356 6308 11408
rect 6360 11396 6366 11408
rect 8053 11399 8111 11405
rect 8053 11396 8065 11399
rect 6360 11368 8065 11396
rect 6360 11356 6366 11368
rect 8053 11365 8065 11368
rect 8099 11396 8111 11399
rect 8234 11396 8240 11408
rect 8099 11368 8240 11396
rect 8099 11365 8111 11368
rect 8053 11359 8111 11365
rect 8234 11356 8240 11368
rect 8292 11356 8298 11408
rect 11178 11356 11184 11408
rect 11236 11396 11242 11408
rect 11638 11396 11644 11408
rect 11236 11368 11644 11396
rect 11236 11356 11242 11368
rect 11638 11356 11644 11368
rect 11696 11356 11702 11408
rect 13018 11396 13024 11408
rect 12979 11368 13024 11396
rect 13018 11356 13024 11368
rect 13076 11356 13082 11408
rect 13202 11396 13208 11408
rect 13163 11368 13208 11396
rect 13202 11356 13208 11368
rect 13260 11356 13266 11408
rect 13294 11356 13300 11408
rect 13352 11396 13358 11408
rect 13389 11399 13447 11405
rect 13389 11396 13401 11399
rect 13352 11368 13401 11396
rect 13352 11356 13358 11368
rect 13389 11365 13401 11368
rect 13435 11365 13447 11399
rect 13389 11359 13447 11365
rect 13938 11356 13944 11408
rect 13996 11396 14002 11408
rect 14766 11396 14772 11408
rect 13996 11368 14772 11396
rect 13996 11356 14002 11368
rect 14766 11356 14772 11368
rect 14824 11356 14830 11408
rect 400 11306 27264 11328
rect 400 11254 3510 11306
rect 3562 11254 3574 11306
rect 3626 11254 3638 11306
rect 3690 11254 3702 11306
rect 3754 11254 3766 11306
rect 3818 11254 27264 11306
rect 400 11232 27264 11254
rect 1610 11192 1616 11204
rect 1571 11164 1616 11192
rect 1610 11152 1616 11164
rect 1668 11152 1674 11204
rect 1794 11192 1800 11204
rect 1755 11164 1800 11192
rect 1794 11152 1800 11164
rect 1852 11152 1858 11204
rect 2346 11192 2352 11204
rect 2307 11164 2352 11192
rect 2346 11152 2352 11164
rect 2404 11152 2410 11204
rect 2530 11152 2536 11204
rect 2588 11192 2594 11204
rect 3358 11192 3364 11204
rect 2588 11164 3364 11192
rect 2588 11152 2594 11164
rect 3358 11152 3364 11164
rect 3416 11152 3422 11204
rect 3821 11195 3879 11201
rect 3821 11161 3833 11195
rect 3867 11192 3879 11195
rect 4002 11192 4008 11204
rect 3867 11164 4008 11192
rect 3867 11161 3879 11164
rect 3821 11155 3879 11161
rect 4002 11152 4008 11164
rect 4060 11152 4066 11204
rect 4370 11192 4376 11204
rect 4331 11164 4376 11192
rect 4370 11152 4376 11164
rect 4428 11152 4434 11204
rect 4462 11152 4468 11204
rect 4520 11192 4526 11204
rect 4741 11195 4799 11201
rect 4741 11192 4753 11195
rect 4520 11164 4753 11192
rect 4520 11152 4526 11164
rect 4741 11161 4753 11164
rect 4787 11161 4799 11195
rect 4741 11155 4799 11161
rect 5934 11152 5940 11204
rect 5992 11192 5998 11204
rect 6489 11195 6547 11201
rect 6489 11192 6501 11195
rect 5992 11164 6501 11192
rect 5992 11152 5998 11164
rect 6489 11161 6501 11164
rect 6535 11161 6547 11195
rect 6670 11192 6676 11204
rect 6631 11164 6676 11192
rect 6489 11155 6547 11161
rect 6670 11152 6676 11164
rect 6728 11152 6734 11204
rect 7774 11192 7780 11204
rect 7608 11164 7780 11192
rect 3910 11084 3916 11136
rect 3968 11124 3974 11136
rect 4189 11127 4247 11133
rect 4189 11124 4201 11127
rect 3968 11096 4201 11124
rect 3968 11084 3974 11096
rect 4189 11093 4201 11096
rect 4235 11093 4247 11127
rect 4646 11124 4652 11136
rect 4189 11087 4247 11093
rect 4296 11096 4652 11124
rect 2809 11059 2867 11065
rect 2809 11025 2821 11059
rect 2855 11056 2867 11059
rect 2898 11056 2904 11068
rect 2855 11028 2904 11056
rect 2855 11025 2867 11028
rect 2809 11019 2867 11025
rect 2257 10991 2315 10997
rect 2257 10957 2269 10991
rect 2303 10988 2315 10991
rect 2622 10988 2628 11000
rect 2303 10960 2628 10988
rect 2303 10957 2315 10960
rect 2257 10951 2315 10957
rect 2622 10948 2628 10960
rect 2680 10988 2686 11000
rect 2824 10988 2852 11019
rect 2898 11016 2904 11028
rect 2956 11016 2962 11068
rect 4296 11065 4324 11096
rect 4646 11084 4652 11096
rect 4704 11084 4710 11136
rect 5566 11084 5572 11136
rect 5624 11124 5630 11136
rect 6121 11127 6179 11133
rect 6121 11124 6133 11127
rect 5624 11096 6133 11124
rect 5624 11084 5630 11096
rect 6121 11093 6133 11096
rect 6167 11093 6179 11127
rect 6394 11124 6400 11136
rect 6355 11096 6400 11124
rect 6121 11087 6179 11093
rect 6394 11084 6400 11096
rect 6452 11084 6458 11136
rect 7608 11133 7636 11164
rect 7774 11152 7780 11164
rect 7832 11152 7838 11204
rect 9985 11195 10043 11201
rect 9985 11161 9997 11195
rect 10031 11192 10043 11195
rect 10166 11192 10172 11204
rect 10031 11164 10172 11192
rect 10031 11161 10043 11164
rect 9985 11155 10043 11161
rect 10166 11152 10172 11164
rect 10224 11152 10230 11204
rect 10810 11192 10816 11204
rect 10771 11164 10816 11192
rect 10810 11152 10816 11164
rect 10868 11152 10874 11204
rect 13938 11192 13944 11204
rect 13899 11164 13944 11192
rect 13938 11152 13944 11164
rect 13996 11152 14002 11204
rect 14122 11152 14128 11204
rect 14180 11192 14186 11204
rect 14214 11192 14220 11204
rect 14180 11164 14220 11192
rect 14180 11152 14186 11164
rect 14214 11152 14220 11164
rect 14272 11152 14278 11204
rect 14658 11195 14716 11201
rect 14658 11192 14670 11195
rect 14324 11164 14670 11192
rect 7593 11127 7651 11133
rect 7593 11093 7605 11127
rect 7639 11093 7651 11127
rect 9430 11124 9436 11136
rect 7593 11087 7651 11093
rect 7700 11096 9436 11124
rect 3637 11059 3695 11065
rect 3637 11025 3649 11059
rect 3683 11056 3695 11059
rect 4281 11059 4339 11065
rect 4281 11056 4293 11059
rect 3683 11028 4293 11056
rect 3683 11025 3695 11028
rect 3637 11019 3695 11025
rect 4281 11025 4293 11028
rect 4327 11025 4339 11059
rect 7700 11056 7728 11096
rect 9430 11084 9436 11096
rect 9488 11084 9494 11136
rect 9614 11084 9620 11136
rect 9672 11124 9678 11136
rect 13478 11124 13484 11136
rect 9672 11096 13484 11124
rect 9672 11084 9678 11096
rect 13478 11084 13484 11096
rect 13536 11084 13542 11136
rect 13849 11127 13907 11133
rect 13849 11124 13861 11127
rect 13680 11096 13861 11124
rect 8878 11056 8884 11068
rect 4281 11019 4339 11025
rect 4664 11028 7728 11056
rect 7792 11028 8884 11056
rect 4664 11000 4692 11028
rect 3266 10988 3272 11000
rect 2680 10960 2852 10988
rect 3227 10960 3272 10988
rect 2680 10948 2686 10960
rect 3266 10948 3272 10960
rect 3324 10988 3330 11000
rect 4060 10991 4118 10997
rect 4060 10988 4072 10991
rect 3324 10960 4072 10988
rect 3324 10948 3330 10960
rect 4060 10957 4072 10960
rect 4106 10957 4118 10991
rect 4060 10951 4118 10957
rect 4186 10948 4192 11000
rect 4244 10988 4250 11000
rect 4646 10988 4652 11000
rect 4244 10960 4652 10988
rect 4244 10948 4250 10960
rect 4646 10948 4652 10960
rect 4704 10948 4710 11000
rect 4738 10948 4744 11000
rect 4796 10988 4802 11000
rect 7792 10997 7820 11028
rect 8878 11016 8884 11028
rect 8936 11056 8942 11068
rect 9706 11056 9712 11068
rect 8936 11028 9712 11056
rect 8936 11016 8942 11028
rect 9706 11016 9712 11028
rect 9764 11016 9770 11068
rect 10166 11016 10172 11068
rect 10224 11056 10230 11068
rect 10905 11059 10963 11065
rect 10905 11056 10917 11059
rect 10224 11028 10917 11056
rect 10224 11016 10230 11028
rect 10905 11025 10917 11028
rect 10951 11025 10963 11059
rect 10905 11019 10963 11025
rect 11730 11016 11736 11068
rect 11788 11056 11794 11068
rect 12285 11059 12343 11065
rect 12285 11056 12297 11059
rect 11788 11028 12297 11056
rect 11788 11016 11794 11028
rect 12285 11025 12297 11028
rect 12331 11056 12343 11059
rect 12653 11059 12711 11065
rect 12653 11056 12665 11059
rect 12331 11028 12665 11056
rect 12331 11025 12343 11028
rect 12285 11019 12343 11025
rect 12653 11025 12665 11028
rect 12699 11025 12711 11059
rect 12834 11056 12840 11068
rect 12747 11028 12840 11056
rect 12653 11019 12711 11025
rect 12834 11016 12840 11028
rect 12892 11056 12898 11068
rect 13680 11065 13708 11096
rect 13849 11093 13861 11096
rect 13895 11124 13907 11127
rect 14324 11124 14352 11164
rect 14658 11161 14670 11164
rect 14704 11192 14716 11195
rect 15321 11195 15379 11201
rect 15321 11192 15333 11195
rect 14704 11164 15333 11192
rect 14704 11161 14716 11164
rect 14658 11155 14716 11161
rect 15321 11161 15333 11164
rect 15367 11161 15379 11195
rect 24426 11192 24432 11204
rect 24387 11164 24432 11192
rect 15321 11155 15379 11161
rect 24426 11152 24432 11164
rect 24484 11152 24490 11204
rect 24702 11192 24708 11204
rect 24663 11164 24708 11192
rect 24702 11152 24708 11164
rect 24760 11152 24766 11204
rect 14766 11124 14772 11136
rect 13895 11096 14352 11124
rect 14727 11096 14772 11124
rect 13895 11093 13907 11096
rect 13849 11087 13907 11093
rect 14766 11084 14772 11096
rect 14824 11084 14830 11136
rect 18173 11127 18231 11133
rect 18173 11093 18185 11127
rect 18219 11124 18231 11127
rect 18541 11127 18599 11133
rect 18541 11124 18553 11127
rect 18219 11096 18553 11124
rect 18219 11093 18231 11096
rect 18173 11087 18231 11093
rect 18541 11093 18553 11096
rect 18587 11124 18599 11127
rect 19274 11124 19280 11136
rect 18587 11096 19280 11124
rect 18587 11093 18599 11096
rect 18541 11087 18599 11093
rect 19274 11084 19280 11096
rect 19332 11084 19338 11136
rect 13665 11059 13723 11065
rect 13665 11056 13677 11059
rect 12892 11028 13677 11056
rect 12892 11016 12898 11028
rect 13665 11025 13677 11028
rect 13711 11025 13723 11059
rect 13665 11019 13723 11025
rect 14401 11059 14459 11065
rect 14401 11025 14413 11059
rect 14447 11056 14459 11059
rect 14858 11056 14864 11068
rect 14447 11028 14628 11056
rect 14819 11028 14864 11056
rect 14447 11025 14459 11028
rect 14401 11019 14459 11025
rect 4925 10991 4983 10997
rect 4925 10988 4937 10991
rect 4796 10960 4937 10988
rect 4796 10948 4802 10960
rect 4925 10957 4937 10960
rect 4971 10957 4983 10991
rect 4925 10951 4983 10957
rect 7041 10991 7099 10997
rect 7041 10957 7053 10991
rect 7087 10988 7099 10991
rect 7777 10991 7835 10997
rect 7777 10988 7789 10991
rect 7087 10960 7789 10988
rect 7087 10957 7099 10960
rect 7041 10951 7099 10957
rect 7777 10957 7789 10960
rect 7823 10957 7835 10991
rect 7777 10951 7835 10957
rect 7866 10948 7872 11000
rect 7924 10988 7930 11000
rect 7961 10991 8019 10997
rect 7961 10988 7973 10991
rect 7924 10960 7973 10988
rect 7924 10948 7930 10960
rect 7961 10957 7973 10960
rect 8007 10957 8019 10991
rect 7961 10951 8019 10957
rect 8145 10991 8203 10997
rect 8145 10957 8157 10991
rect 8191 10957 8203 10991
rect 8145 10951 8203 10957
rect 1518 10880 1524 10932
rect 1576 10920 1582 10932
rect 1889 10923 1947 10929
rect 1889 10920 1901 10923
rect 1576 10892 1901 10920
rect 1576 10880 1582 10892
rect 1889 10889 1901 10892
rect 1935 10889 1947 10923
rect 1889 10883 1947 10889
rect 2073 10923 2131 10929
rect 2073 10889 2085 10923
rect 2119 10920 2131 10923
rect 2119 10892 3036 10920
rect 2119 10889 2131 10892
rect 2073 10883 2131 10889
rect 3008 10864 3036 10892
rect 3358 10880 3364 10932
rect 3416 10920 3422 10932
rect 3913 10923 3971 10929
rect 3913 10920 3925 10923
rect 3416 10892 3925 10920
rect 3416 10880 3422 10892
rect 3913 10889 3925 10892
rect 3959 10889 3971 10923
rect 3913 10883 3971 10889
rect 2990 10852 2996 10864
rect 2951 10824 2996 10852
rect 2990 10812 2996 10824
rect 3048 10812 3054 10864
rect 5198 10852 5204 10864
rect 5159 10824 5204 10852
rect 5198 10812 5204 10824
rect 5256 10812 5262 10864
rect 7222 10852 7228 10864
rect 7183 10824 7228 10852
rect 7222 10812 7228 10824
rect 7280 10852 7286 10864
rect 8160 10852 8188 10951
rect 8602 10948 8608 11000
rect 8660 10988 8666 11000
rect 9157 10991 9215 10997
rect 9157 10988 9169 10991
rect 8660 10960 9169 10988
rect 8660 10948 8666 10960
rect 9157 10957 9169 10960
rect 9203 10957 9215 10991
rect 9157 10951 9215 10957
rect 9522 10948 9528 11000
rect 9580 10988 9586 11000
rect 9617 10991 9675 10997
rect 9617 10988 9629 10991
rect 9580 10960 9629 10988
rect 9580 10948 9586 10960
rect 9617 10957 9629 10960
rect 9663 10988 9675 10991
rect 11270 10988 11276 11000
rect 9663 10960 11276 10988
rect 9663 10957 9675 10960
rect 9617 10951 9675 10957
rect 11270 10948 11276 10960
rect 11328 10948 11334 11000
rect 11917 10991 11975 10997
rect 11917 10957 11929 10991
rect 11963 10988 11975 10991
rect 12377 10991 12435 10997
rect 12377 10988 12389 10991
rect 11963 10960 12389 10988
rect 11963 10957 11975 10960
rect 11917 10951 11975 10957
rect 12377 10957 12389 10960
rect 12423 10988 12435 10991
rect 12558 10988 12564 11000
rect 12423 10960 12564 10988
rect 12423 10957 12435 10960
rect 12377 10951 12435 10957
rect 12558 10948 12564 10960
rect 12616 10948 12622 11000
rect 13113 10991 13171 10997
rect 13113 10957 13125 10991
rect 13159 10988 13171 10991
rect 13202 10988 13208 11000
rect 13159 10960 13208 10988
rect 13159 10957 13171 10960
rect 13113 10951 13171 10957
rect 8694 10880 8700 10932
rect 8752 10920 8758 10932
rect 9338 10920 9344 10932
rect 8752 10892 9344 10920
rect 8752 10880 8758 10892
rect 9338 10880 9344 10892
rect 9396 10880 9402 10932
rect 11178 10880 11184 10932
rect 11236 10920 11242 10932
rect 11549 10923 11607 10929
rect 11549 10920 11561 10923
rect 11236 10892 11561 10920
rect 11236 10880 11242 10892
rect 11549 10889 11561 10892
rect 11595 10920 11607 10923
rect 11733 10923 11791 10929
rect 11733 10920 11745 10923
rect 11595 10892 11745 10920
rect 11595 10889 11607 10892
rect 11549 10883 11607 10889
rect 11733 10889 11745 10892
rect 11779 10920 11791 10923
rect 13128 10920 13156 10951
rect 13202 10948 13208 10960
rect 13260 10948 13266 11000
rect 13294 10948 13300 11000
rect 13352 10988 13358 11000
rect 13352 10960 13397 10988
rect 13352 10948 13358 10960
rect 11779 10892 13156 10920
rect 11779 10889 11791 10892
rect 11733 10883 11791 10889
rect 14214 10880 14220 10932
rect 14272 10920 14278 10932
rect 14493 10923 14551 10929
rect 14272 10892 14444 10920
rect 14272 10880 14278 10892
rect 9062 10852 9068 10864
rect 7280 10824 9068 10852
rect 7280 10812 7286 10824
rect 9062 10812 9068 10824
rect 9120 10812 9126 10864
rect 12282 10812 12288 10864
rect 12340 10852 12346 10864
rect 12929 10855 12987 10861
rect 12929 10852 12941 10855
rect 12340 10824 12941 10852
rect 12340 10812 12346 10824
rect 12929 10821 12941 10824
rect 12975 10852 12987 10855
rect 13018 10852 13024 10864
rect 12975 10824 13024 10852
rect 12975 10821 12987 10824
rect 12929 10815 12987 10821
rect 13018 10812 13024 10824
rect 13076 10812 13082 10864
rect 14416 10852 14444 10892
rect 14493 10889 14505 10923
rect 14539 10920 14551 10923
rect 14600 10920 14628 11028
rect 14858 11016 14864 11028
rect 14916 11016 14922 11068
rect 15502 11016 15508 11068
rect 15560 11056 15566 11068
rect 21669 11059 21727 11065
rect 21669 11056 21681 11059
rect 15560 11028 21681 11056
rect 15560 11016 15566 11028
rect 18357 10991 18415 10997
rect 18357 10957 18369 10991
rect 18403 10988 18415 10991
rect 18722 10988 18728 11000
rect 18403 10960 18728 10988
rect 18403 10957 18415 10960
rect 18357 10951 18415 10957
rect 18722 10948 18728 10960
rect 18780 10948 18786 11000
rect 19185 10991 19243 10997
rect 19185 10957 19197 10991
rect 19231 10988 19243 10991
rect 19277 10991 19335 10997
rect 19277 10988 19289 10991
rect 19231 10960 19289 10988
rect 19231 10957 19243 10960
rect 19185 10951 19243 10957
rect 19277 10957 19289 10960
rect 19323 10988 19335 10991
rect 19366 10988 19372 11000
rect 19323 10960 19372 10988
rect 19323 10957 19335 10960
rect 19277 10951 19335 10957
rect 19366 10948 19372 10960
rect 19424 10948 19430 11000
rect 21132 10997 21160 11028
rect 21669 11025 21681 11028
rect 21715 11056 21727 11059
rect 24426 11056 24432 11068
rect 21715 11028 24432 11056
rect 21715 11025 21727 11028
rect 21669 11019 21727 11025
rect 24426 11016 24432 11028
rect 24484 11016 24490 11068
rect 21117 10991 21175 10997
rect 21117 10957 21129 10991
rect 21163 10957 21175 10991
rect 21117 10951 21175 10957
rect 17986 10920 17992 10932
rect 14539 10892 17992 10920
rect 14539 10889 14551 10892
rect 14493 10883 14551 10889
rect 17986 10880 17992 10892
rect 18044 10880 18050 10932
rect 20930 10880 20936 10932
rect 20988 10920 20994 10932
rect 21393 10923 21451 10929
rect 21393 10920 21405 10923
rect 20988 10892 21405 10920
rect 20988 10880 20994 10892
rect 21393 10889 21405 10892
rect 21439 10920 21451 10923
rect 21853 10923 21911 10929
rect 21853 10920 21865 10923
rect 21439 10892 21865 10920
rect 21439 10889 21451 10892
rect 21393 10883 21451 10889
rect 21853 10889 21865 10892
rect 21899 10889 21911 10923
rect 21853 10883 21911 10889
rect 15137 10855 15195 10861
rect 15137 10852 15149 10855
rect 14416 10824 15149 10852
rect 15137 10821 15149 10824
rect 15183 10821 15195 10855
rect 15137 10815 15195 10821
rect 400 10762 27264 10784
rect 400 10710 18870 10762
rect 18922 10710 18934 10762
rect 18986 10710 18998 10762
rect 19050 10710 19062 10762
rect 19114 10710 19126 10762
rect 19178 10710 27264 10762
rect 400 10688 27264 10710
rect 1797 10651 1855 10657
rect 1797 10617 1809 10651
rect 1843 10648 1855 10651
rect 2070 10648 2076 10660
rect 1843 10620 2076 10648
rect 1843 10617 1855 10620
rect 1797 10611 1855 10617
rect 2070 10608 2076 10620
rect 2128 10608 2134 10660
rect 2165 10651 2223 10657
rect 2165 10617 2177 10651
rect 2211 10648 2223 10651
rect 2346 10648 2352 10660
rect 2211 10620 2352 10648
rect 2211 10617 2223 10620
rect 2165 10611 2223 10617
rect 2346 10608 2352 10620
rect 2404 10608 2410 10660
rect 2990 10608 2996 10660
rect 3048 10648 3054 10660
rect 4278 10648 4284 10660
rect 3048 10620 4284 10648
rect 3048 10608 3054 10620
rect 4278 10608 4284 10620
rect 4336 10608 4342 10660
rect 4462 10608 4468 10660
rect 4520 10648 4526 10660
rect 4557 10651 4615 10657
rect 4557 10648 4569 10651
rect 4520 10620 4569 10648
rect 4520 10608 4526 10620
rect 4557 10617 4569 10620
rect 4603 10617 4615 10651
rect 4557 10611 4615 10617
rect 7409 10651 7467 10657
rect 7409 10617 7421 10651
rect 7455 10648 7467 10651
rect 7774 10648 7780 10660
rect 7455 10620 7780 10648
rect 7455 10617 7467 10620
rect 7409 10611 7467 10617
rect 7774 10608 7780 10620
rect 7832 10608 7838 10660
rect 8510 10608 8516 10660
rect 8568 10648 8574 10660
rect 8568 10620 9752 10648
rect 8568 10608 8574 10620
rect 4373 10583 4431 10589
rect 4373 10580 4385 10583
rect 3744 10552 4385 10580
rect 3174 10472 3180 10524
rect 3232 10512 3238 10524
rect 3744 10521 3772 10552
rect 4373 10549 4385 10552
rect 4419 10580 4431 10583
rect 4922 10580 4928 10592
rect 4419 10552 4928 10580
rect 4419 10549 4431 10552
rect 4373 10543 4431 10549
rect 4922 10540 4928 10552
rect 4980 10540 4986 10592
rect 5658 10580 5664 10592
rect 5619 10552 5664 10580
rect 5658 10540 5664 10552
rect 5716 10540 5722 10592
rect 8326 10540 8332 10592
rect 8384 10580 8390 10592
rect 8786 10580 8792 10592
rect 8384 10552 8792 10580
rect 8384 10540 8390 10552
rect 8786 10540 8792 10552
rect 8844 10580 8850 10592
rect 8973 10583 9031 10589
rect 8973 10580 8985 10583
rect 8844 10552 8985 10580
rect 8844 10540 8850 10552
rect 8973 10549 8985 10552
rect 9019 10549 9031 10583
rect 8973 10543 9031 10549
rect 9062 10540 9068 10592
rect 9120 10580 9126 10592
rect 9157 10583 9215 10589
rect 9157 10580 9169 10583
rect 9120 10552 9169 10580
rect 9120 10540 9126 10552
rect 9157 10549 9169 10552
rect 9203 10549 9215 10583
rect 9157 10543 9215 10549
rect 9341 10583 9399 10589
rect 9341 10549 9353 10583
rect 9387 10580 9399 10583
rect 9430 10580 9436 10592
rect 9387 10552 9436 10580
rect 9387 10549 9399 10552
rect 9341 10543 9399 10549
rect 9430 10540 9436 10552
rect 9488 10540 9494 10592
rect 9724 10589 9752 10620
rect 14766 10608 14772 10660
rect 14824 10648 14830 10660
rect 19274 10648 19280 10660
rect 14824 10620 15824 10648
rect 19235 10620 19280 10648
rect 14824 10608 14830 10620
rect 9709 10583 9767 10589
rect 9709 10549 9721 10583
rect 9755 10549 9767 10583
rect 14214 10580 14220 10592
rect 9709 10543 9767 10549
rect 13404 10552 14220 10580
rect 3729 10515 3787 10521
rect 3729 10512 3741 10515
rect 3232 10484 3741 10512
rect 3232 10472 3238 10484
rect 3729 10481 3741 10484
rect 3775 10481 3787 10515
rect 3910 10512 3916 10524
rect 3871 10484 3916 10512
rect 3729 10475 3787 10481
rect 3910 10472 3916 10484
rect 3968 10472 3974 10524
rect 4278 10512 4284 10524
rect 4239 10484 4284 10512
rect 4278 10472 4284 10484
rect 4336 10472 4342 10524
rect 4462 10472 4468 10524
rect 4520 10512 4526 10524
rect 5109 10515 5167 10521
rect 5109 10512 5121 10515
rect 4520 10484 5121 10512
rect 4520 10472 4526 10484
rect 5109 10481 5121 10484
rect 5155 10481 5167 10515
rect 5290 10512 5296 10524
rect 5251 10484 5296 10512
rect 5109 10475 5167 10481
rect 5290 10472 5296 10484
rect 5348 10472 5354 10524
rect 9246 10512 9252 10524
rect 9207 10484 9252 10512
rect 9246 10472 9252 10484
rect 9304 10472 9310 10524
rect 12282 10512 12288 10524
rect 12243 10484 12288 10512
rect 12282 10472 12288 10484
rect 12340 10472 12346 10524
rect 12742 10512 12748 10524
rect 12703 10484 12748 10512
rect 12742 10472 12748 10484
rect 12800 10472 12806 10524
rect 13113 10515 13171 10521
rect 13113 10481 13125 10515
rect 13159 10512 13171 10515
rect 13404 10512 13432 10552
rect 14214 10540 14220 10552
rect 14272 10580 14278 10592
rect 14272 10552 15732 10580
rect 14272 10540 14278 10552
rect 13159 10484 13432 10512
rect 13159 10481 13171 10484
rect 13113 10475 13171 10481
rect 13846 10472 13852 10524
rect 13904 10512 13910 10524
rect 15229 10515 15287 10521
rect 15229 10512 15241 10515
rect 13904 10484 15241 10512
rect 13904 10472 13910 10484
rect 15229 10481 15241 10484
rect 15275 10481 15287 10515
rect 15594 10512 15600 10524
rect 15555 10484 15600 10512
rect 15229 10475 15287 10481
rect 15594 10472 15600 10484
rect 15652 10472 15658 10524
rect 15704 10521 15732 10552
rect 15689 10515 15747 10521
rect 15689 10481 15701 10515
rect 15735 10481 15747 10515
rect 15796 10512 15824 10620
rect 19274 10608 19280 10620
rect 19332 10608 19338 10660
rect 20212 10620 21804 10648
rect 15870 10540 15876 10592
rect 15928 10580 15934 10592
rect 20212 10580 20240 10620
rect 15928 10552 20240 10580
rect 15928 10540 15934 10552
rect 17805 10515 17863 10521
rect 17805 10512 17817 10515
rect 15796 10484 17817 10512
rect 15689 10475 15747 10481
rect 17805 10481 17817 10484
rect 17851 10481 17863 10515
rect 17986 10512 17992 10524
rect 17947 10484 17992 10512
rect 17805 10475 17863 10481
rect 4738 10404 4744 10456
rect 4796 10444 4802 10456
rect 8605 10447 8663 10453
rect 8605 10444 8617 10447
rect 4796 10416 8617 10444
rect 4796 10404 4802 10416
rect 8605 10413 8617 10416
rect 8651 10444 8663 10447
rect 8694 10444 8700 10456
rect 8651 10416 8700 10444
rect 8651 10413 8663 10416
rect 8605 10407 8663 10413
rect 8694 10404 8700 10416
rect 8752 10404 8758 10456
rect 15318 10444 15324 10456
rect 13128 10416 15324 10444
rect 13128 10388 13156 10416
rect 15318 10404 15324 10416
rect 15376 10404 15382 10456
rect 17820 10444 17848 10475
rect 17986 10472 17992 10484
rect 18044 10472 18050 10524
rect 18354 10512 18360 10524
rect 18315 10484 18360 10512
rect 18354 10472 18360 10484
rect 18412 10472 18418 10524
rect 18538 10512 18544 10524
rect 18499 10484 18544 10512
rect 18538 10472 18544 10484
rect 18596 10472 18602 10524
rect 20212 10521 20240 10552
rect 20930 10540 20936 10592
rect 20988 10540 20994 10592
rect 21776 10580 21804 10620
rect 22678 10608 22684 10660
rect 22736 10648 22742 10660
rect 23141 10651 23199 10657
rect 23141 10648 23153 10651
rect 22736 10620 23153 10648
rect 22736 10608 22742 10620
rect 23141 10617 23153 10620
rect 23187 10648 23199 10651
rect 23230 10648 23236 10660
rect 23187 10620 23236 10648
rect 23187 10617 23199 10620
rect 23141 10611 23199 10617
rect 23230 10608 23236 10620
rect 23288 10608 23294 10660
rect 23782 10648 23788 10660
rect 23743 10620 23788 10648
rect 23782 10608 23788 10620
rect 23840 10608 23846 10660
rect 23800 10580 23828 10608
rect 21776 10552 23828 10580
rect 20197 10515 20255 10521
rect 20197 10481 20209 10515
rect 20243 10481 20255 10515
rect 20197 10475 20255 10481
rect 23046 10472 23052 10524
rect 23104 10512 23110 10524
rect 23322 10512 23328 10524
rect 23104 10484 23328 10512
rect 23104 10472 23110 10484
rect 23322 10472 23328 10484
rect 23380 10472 23386 10524
rect 23782 10472 23788 10524
rect 23840 10512 23846 10524
rect 24426 10512 24432 10524
rect 23840 10484 24432 10512
rect 23840 10472 23846 10484
rect 24426 10472 24432 10484
rect 24484 10472 24490 10524
rect 18078 10444 18084 10456
rect 17820 10416 18084 10444
rect 18078 10404 18084 10416
rect 18136 10404 18142 10456
rect 20470 10444 20476 10456
rect 20431 10416 20476 10444
rect 20470 10404 20476 10416
rect 20528 10404 20534 10456
rect 22218 10444 22224 10456
rect 22179 10416 22224 10444
rect 22218 10404 22224 10416
rect 22276 10404 22282 10456
rect 23506 10404 23512 10456
rect 23564 10444 23570 10456
rect 24702 10444 24708 10456
rect 23564 10416 24708 10444
rect 23564 10404 23570 10416
rect 24702 10404 24708 10416
rect 24760 10404 24766 10456
rect 4646 10376 4652 10388
rect 4526 10348 4652 10376
rect 3910 10268 3916 10320
rect 3968 10308 3974 10320
rect 4526 10308 4554 10348
rect 4646 10336 4652 10348
rect 4704 10336 4710 10388
rect 8234 10336 8240 10388
rect 8292 10376 8298 10388
rect 9522 10376 9528 10388
rect 8292 10348 9528 10376
rect 8292 10336 8298 10348
rect 9522 10336 9528 10348
rect 9580 10336 9586 10388
rect 13110 10376 13116 10388
rect 13071 10348 13116 10376
rect 13110 10336 13116 10348
rect 13168 10336 13174 10388
rect 18096 10376 18124 10404
rect 19461 10379 19519 10385
rect 19461 10376 19473 10379
rect 18096 10348 19473 10376
rect 19461 10345 19473 10348
rect 19507 10376 19519 10379
rect 19507 10348 19734 10376
rect 19507 10345 19519 10348
rect 19461 10339 19519 10345
rect 14398 10308 14404 10320
rect 3968 10280 4554 10308
rect 14359 10280 14404 10308
rect 3968 10268 3974 10280
rect 14398 10268 14404 10280
rect 14456 10268 14462 10320
rect 14677 10311 14735 10317
rect 14677 10277 14689 10311
rect 14723 10308 14735 10311
rect 15134 10308 15140 10320
rect 14723 10280 15140 10308
rect 14723 10277 14735 10280
rect 14677 10271 14735 10277
rect 15134 10268 15140 10280
rect 15192 10268 15198 10320
rect 16974 10268 16980 10320
rect 17032 10308 17038 10320
rect 17621 10311 17679 10317
rect 17621 10308 17633 10311
rect 17032 10280 17633 10308
rect 17032 10268 17038 10280
rect 17621 10277 17633 10280
rect 17667 10308 17679 10311
rect 18722 10308 18728 10320
rect 17667 10280 18728 10308
rect 17667 10277 17679 10280
rect 17621 10271 17679 10277
rect 18722 10268 18728 10280
rect 18780 10268 18786 10320
rect 19090 10308 19096 10320
rect 19051 10280 19096 10308
rect 19090 10268 19096 10280
rect 19148 10268 19154 10320
rect 19706 10308 19734 10348
rect 20286 10308 20292 10320
rect 19706 10280 20292 10308
rect 20286 10268 20292 10280
rect 20344 10268 20350 10320
rect 24058 10308 24064 10320
rect 24019 10280 24064 10308
rect 24058 10268 24064 10280
rect 24116 10268 24122 10320
rect 400 10218 27264 10240
rect 400 10166 3510 10218
rect 3562 10166 3574 10218
rect 3626 10166 3638 10218
rect 3690 10166 3702 10218
rect 3754 10166 3766 10218
rect 3818 10166 27264 10218
rect 400 10144 27264 10166
rect 1334 10064 1340 10116
rect 1392 10104 1398 10116
rect 1429 10107 1487 10113
rect 1429 10104 1441 10107
rect 1392 10076 1441 10104
rect 1392 10064 1398 10076
rect 1429 10073 1441 10076
rect 1475 10104 1487 10107
rect 1843 10107 1901 10113
rect 1843 10104 1855 10107
rect 1475 10076 1855 10104
rect 1475 10073 1487 10076
rect 1429 10067 1487 10073
rect 1843 10073 1855 10076
rect 1889 10073 1901 10107
rect 2622 10104 2628 10116
rect 2583 10076 2628 10104
rect 1843 10067 1901 10073
rect 2622 10064 2628 10076
rect 2680 10064 2686 10116
rect 2990 10104 2996 10116
rect 2951 10076 2996 10104
rect 2990 10064 2996 10076
rect 3048 10064 3054 10116
rect 3174 10104 3180 10116
rect 3135 10076 3180 10104
rect 3174 10064 3180 10076
rect 3232 10064 3238 10116
rect 4186 10104 4192 10116
rect 4147 10076 4192 10104
rect 4186 10064 4192 10076
rect 4244 10064 4250 10116
rect 4557 10107 4615 10113
rect 4557 10073 4569 10107
rect 4603 10104 4615 10107
rect 4646 10104 4652 10116
rect 4603 10076 4652 10104
rect 4603 10073 4615 10076
rect 4557 10067 4615 10073
rect 4646 10064 4652 10076
rect 4704 10064 4710 10116
rect 5201 10107 5259 10113
rect 5201 10073 5213 10107
rect 5247 10104 5259 10107
rect 5290 10104 5296 10116
rect 5247 10076 5296 10104
rect 5247 10073 5259 10076
rect 5201 10067 5259 10073
rect 5290 10064 5296 10076
rect 5348 10064 5354 10116
rect 5569 10107 5627 10113
rect 5569 10073 5581 10107
rect 5615 10104 5627 10107
rect 5658 10104 5664 10116
rect 5615 10076 5664 10104
rect 5615 10073 5627 10076
rect 5569 10067 5627 10073
rect 5658 10064 5664 10076
rect 5716 10064 5722 10116
rect 6762 10104 6768 10116
rect 6723 10076 6768 10104
rect 6762 10064 6768 10076
rect 6820 10104 6826 10116
rect 7130 10104 7136 10116
rect 6820 10076 7136 10104
rect 6820 10064 6826 10076
rect 7130 10064 7136 10076
rect 7188 10104 7194 10116
rect 7225 10107 7283 10113
rect 7225 10104 7237 10107
rect 7188 10076 7237 10104
rect 7188 10064 7194 10076
rect 7225 10073 7237 10076
rect 7271 10073 7283 10107
rect 7225 10067 7283 10073
rect 8145 10107 8203 10113
rect 8145 10073 8157 10107
rect 8191 10104 8203 10107
rect 8510 10104 8516 10116
rect 8191 10076 8516 10104
rect 8191 10073 8203 10076
rect 8145 10067 8203 10073
rect 8510 10064 8516 10076
rect 8568 10064 8574 10116
rect 9062 10064 9068 10116
rect 9120 10104 9126 10116
rect 9801 10107 9859 10113
rect 9801 10104 9813 10107
rect 9120 10076 9813 10104
rect 9120 10064 9126 10076
rect 9801 10073 9813 10076
rect 9847 10073 9859 10107
rect 11454 10104 11460 10116
rect 11415 10076 11460 10104
rect 9801 10067 9859 10073
rect 11454 10064 11460 10076
rect 11512 10104 11518 10116
rect 11825 10107 11883 10113
rect 11825 10104 11837 10107
rect 11512 10076 11837 10104
rect 11512 10064 11518 10076
rect 11825 10073 11837 10076
rect 11871 10104 11883 10107
rect 12653 10107 12711 10113
rect 12653 10104 12665 10107
rect 11871 10076 12665 10104
rect 11871 10073 11883 10076
rect 11825 10067 11883 10073
rect 12653 10073 12665 10076
rect 12699 10104 12711 10107
rect 12742 10104 12748 10116
rect 12699 10076 12748 10104
rect 12699 10073 12711 10076
rect 12653 10067 12711 10073
rect 12742 10064 12748 10076
rect 12800 10064 12806 10116
rect 13110 10104 13116 10116
rect 13071 10076 13116 10104
rect 13110 10064 13116 10076
rect 13168 10064 13174 10116
rect 13846 10104 13852 10116
rect 13807 10076 13852 10104
rect 13846 10064 13852 10076
rect 13904 10064 13910 10116
rect 14401 10107 14459 10113
rect 14401 10073 14413 10107
rect 14447 10104 14459 10107
rect 14490 10104 14496 10116
rect 14447 10076 14496 10104
rect 14447 10073 14459 10076
rect 14401 10067 14459 10073
rect 14490 10064 14496 10076
rect 14548 10064 14554 10116
rect 16974 10104 16980 10116
rect 16935 10076 16980 10104
rect 16974 10064 16980 10076
rect 17032 10064 17038 10116
rect 17342 10064 17348 10116
rect 17400 10104 17406 10116
rect 18538 10104 18544 10116
rect 17400 10076 18544 10104
rect 17400 10064 17406 10076
rect 18538 10064 18544 10076
rect 18596 10064 18602 10116
rect 19001 10107 19059 10113
rect 19001 10073 19013 10107
rect 19047 10104 19059 10107
rect 20470 10104 20476 10116
rect 19047 10076 20476 10104
rect 19047 10073 19059 10076
rect 19001 10067 19059 10073
rect 1613 10039 1671 10045
rect 1613 10005 1625 10039
rect 1659 10036 1671 10039
rect 1981 10039 2039 10045
rect 1981 10036 1993 10039
rect 1659 10008 1993 10036
rect 1659 10005 1671 10008
rect 1613 9999 1671 10005
rect 1981 10005 1993 10008
rect 2027 10036 2039 10039
rect 3082 10036 3088 10048
rect 2027 10008 3088 10036
rect 2027 10005 2039 10008
rect 1981 9999 2039 10005
rect 3082 9996 3088 10008
rect 3140 9996 3146 10048
rect 7869 10039 7927 10045
rect 7869 10005 7881 10039
rect 7915 10036 7927 10039
rect 8234 10036 8240 10048
rect 7915 10008 8240 10036
rect 7915 10005 7927 10008
rect 7869 9999 7927 10005
rect 2073 9971 2131 9977
rect 2073 9937 2085 9971
rect 2119 9968 2131 9971
rect 2622 9968 2628 9980
rect 2119 9940 2628 9968
rect 2119 9937 2131 9940
rect 2073 9931 2131 9937
rect 2622 9928 2628 9940
rect 2680 9928 2686 9980
rect 4281 9971 4339 9977
rect 4281 9968 4293 9971
rect 3468 9940 4293 9968
rect 2640 9900 2668 9928
rect 3468 9909 3496 9940
rect 4281 9937 4293 9940
rect 4327 9937 4339 9971
rect 7222 9968 7228 9980
rect 4281 9931 4339 9937
rect 6964 9940 7228 9968
rect 3453 9903 3511 9909
rect 3453 9900 3465 9903
rect 2640 9872 3465 9900
rect 3453 9869 3465 9872
rect 3499 9869 3511 9903
rect 3453 9863 3511 9869
rect 3637 9903 3695 9909
rect 3637 9869 3649 9903
rect 3683 9900 3695 9903
rect 4554 9900 4560 9912
rect 3683 9872 4560 9900
rect 3683 9869 3695 9872
rect 3637 9863 3695 9869
rect 4554 9860 4560 9872
rect 4612 9860 4618 9912
rect 6118 9860 6124 9912
rect 6176 9900 6182 9912
rect 6964 9909 6992 9940
rect 7222 9928 7228 9940
rect 7280 9968 7286 9980
rect 7593 9971 7651 9977
rect 7593 9968 7605 9971
rect 7280 9940 7605 9968
rect 7280 9928 7286 9940
rect 7593 9937 7605 9940
rect 7639 9937 7651 9971
rect 7593 9931 7651 9937
rect 6949 9903 7007 9909
rect 6949 9900 6961 9903
rect 6176 9872 6961 9900
rect 6176 9860 6182 9872
rect 6949 9869 6961 9872
rect 6995 9869 7007 9903
rect 6949 9863 7007 9869
rect 7041 9903 7099 9909
rect 7041 9869 7053 9903
rect 7087 9900 7099 9903
rect 7884 9900 7912 9999
rect 8234 9996 8240 10008
rect 8292 9996 8298 10048
rect 8786 9996 8792 10048
rect 8844 10036 8850 10048
rect 9617 10039 9675 10045
rect 9617 10036 9629 10039
rect 8844 10008 9629 10036
rect 8844 9996 8850 10008
rect 9617 10005 9629 10008
rect 9663 10005 9675 10039
rect 9617 9999 9675 10005
rect 14033 10039 14091 10045
rect 14033 10005 14045 10039
rect 14079 10036 14091 10039
rect 14306 10036 14312 10048
rect 14079 10008 14312 10036
rect 14079 10005 14091 10008
rect 14033 9999 14091 10005
rect 14306 9996 14312 10008
rect 14364 9996 14370 10048
rect 9062 9928 9068 9980
rect 9120 9968 9126 9980
rect 10350 9968 10356 9980
rect 9120 9940 10356 9968
rect 9120 9928 9126 9940
rect 10350 9928 10356 9940
rect 10408 9968 10414 9980
rect 12282 9968 12288 9980
rect 10408 9940 12288 9968
rect 10408 9928 10414 9940
rect 12282 9928 12288 9940
rect 12340 9928 12346 9980
rect 14508 9977 14536 10064
rect 17161 10039 17219 10045
rect 17161 10005 17173 10039
rect 17207 10036 17219 10039
rect 17897 10039 17955 10045
rect 17897 10036 17909 10039
rect 17207 10008 17909 10036
rect 17207 10005 17219 10008
rect 17161 9999 17219 10005
rect 17897 10005 17909 10008
rect 17943 10036 17955 10039
rect 18354 10036 18360 10048
rect 17943 10008 18360 10036
rect 17943 10005 17955 10008
rect 17897 9999 17955 10005
rect 18354 9996 18360 10008
rect 18412 10036 18418 10048
rect 18449 10039 18507 10045
rect 18449 10036 18461 10039
rect 18412 10008 18461 10036
rect 18412 9996 18418 10008
rect 18449 10005 18461 10008
rect 18495 10005 18507 10039
rect 18449 9999 18507 10005
rect 19108 9977 19136 10076
rect 20470 10064 20476 10076
rect 20528 10104 20534 10116
rect 20657 10107 20715 10113
rect 20657 10104 20669 10107
rect 20528 10076 20669 10104
rect 20528 10064 20534 10076
rect 20657 10073 20669 10076
rect 20703 10073 20715 10107
rect 20930 10104 20936 10116
rect 20891 10076 20936 10104
rect 20657 10067 20715 10073
rect 20930 10064 20936 10076
rect 20988 10064 20994 10116
rect 23230 10104 23236 10116
rect 23191 10076 23236 10104
rect 23230 10064 23236 10076
rect 23288 10064 23294 10116
rect 23506 10104 23512 10116
rect 23467 10076 23512 10104
rect 23506 10064 23512 10076
rect 23564 10064 23570 10116
rect 23874 10064 23880 10116
rect 23932 10064 23938 10116
rect 14493 9971 14551 9977
rect 14493 9937 14505 9971
rect 14539 9937 14551 9971
rect 16057 9971 16115 9977
rect 16057 9968 16069 9971
rect 14493 9931 14551 9937
rect 15152 9940 16069 9968
rect 15152 9912 15180 9940
rect 16057 9937 16069 9940
rect 16103 9968 16115 9971
rect 16241 9971 16299 9977
rect 16241 9968 16253 9971
rect 16103 9940 16253 9968
rect 16103 9937 16115 9940
rect 16057 9931 16115 9937
rect 16241 9937 16253 9940
rect 16287 9937 16299 9971
rect 18633 9971 18691 9977
rect 18633 9968 18645 9971
rect 16241 9931 16299 9937
rect 16348 9940 18645 9968
rect 7087 9872 7912 9900
rect 7087 9869 7099 9872
rect 7041 9863 7099 9869
rect 1705 9835 1763 9841
rect 1705 9801 1717 9835
rect 1751 9832 1763 9835
rect 2070 9832 2076 9844
rect 1751 9804 2076 9832
rect 1751 9801 1763 9804
rect 1705 9795 1763 9801
rect 2070 9792 2076 9804
rect 2128 9792 2134 9844
rect 4005 9835 4063 9841
rect 4005 9801 4017 9835
rect 4051 9832 4063 9835
rect 4094 9832 4100 9844
rect 4051 9804 4100 9832
rect 4051 9801 4063 9804
rect 4005 9795 4063 9801
rect 1794 9724 1800 9776
rect 1852 9764 1858 9776
rect 2349 9767 2407 9773
rect 2349 9764 2361 9767
rect 1852 9736 2361 9764
rect 1852 9724 1858 9736
rect 2349 9733 2361 9736
rect 2395 9733 2407 9767
rect 2349 9727 2407 9733
rect 3361 9767 3419 9773
rect 3361 9733 3373 9767
rect 3407 9764 3419 9767
rect 4020 9764 4048 9795
rect 4094 9792 4100 9804
rect 4152 9792 4158 9844
rect 5293 9835 5351 9841
rect 5293 9832 5305 9835
rect 4526 9804 5305 9832
rect 3407 9736 4048 9764
rect 3407 9733 3419 9736
rect 3361 9727 3419 9733
rect 4370 9724 4376 9776
rect 4428 9764 4434 9776
rect 4526 9764 4554 9804
rect 5293 9801 5305 9804
rect 5339 9801 5351 9835
rect 5293 9795 5351 9801
rect 6486 9792 6492 9844
rect 6544 9832 6550 9844
rect 7056 9832 7084 9863
rect 8694 9860 8700 9912
rect 8752 9900 8758 9912
rect 8789 9903 8847 9909
rect 8789 9900 8801 9903
rect 8752 9872 8801 9900
rect 8752 9860 8758 9872
rect 8789 9869 8801 9872
rect 8835 9869 8847 9903
rect 8789 9863 8847 9869
rect 8878 9860 8884 9912
rect 8936 9900 8942 9912
rect 9246 9900 9252 9912
rect 8936 9872 9252 9900
rect 8936 9860 8942 9872
rect 9246 9860 9252 9872
rect 9304 9900 9310 9912
rect 9985 9903 10043 9909
rect 9985 9900 9997 9903
rect 9304 9872 9997 9900
rect 9304 9860 9310 9872
rect 9985 9869 9997 9872
rect 10031 9900 10043 9903
rect 10169 9903 10227 9909
rect 10169 9900 10181 9903
rect 10031 9872 10181 9900
rect 10031 9869 10043 9872
rect 9985 9863 10043 9869
rect 10169 9869 10181 9872
rect 10215 9869 10227 9903
rect 12006 9900 12012 9912
rect 11919 9872 12012 9900
rect 10169 9863 10227 9869
rect 12006 9860 12012 9872
rect 12064 9900 12070 9912
rect 12469 9903 12527 9909
rect 12469 9900 12481 9903
rect 12064 9872 12481 9900
rect 12064 9860 12070 9872
rect 12469 9869 12481 9872
rect 12515 9869 12527 9903
rect 12469 9863 12527 9869
rect 13386 9860 13392 9912
rect 13444 9900 13450 9912
rect 14953 9903 15011 9909
rect 14953 9900 14965 9903
rect 13444 9872 14965 9900
rect 13444 9860 13450 9872
rect 14953 9869 14965 9872
rect 14999 9869 15011 9903
rect 15134 9900 15140 9912
rect 15095 9872 15140 9900
rect 14953 9863 15011 9869
rect 15134 9860 15140 9872
rect 15192 9860 15198 9912
rect 15321 9903 15379 9909
rect 15321 9869 15333 9903
rect 15367 9869 15379 9903
rect 15594 9900 15600 9912
rect 15555 9872 15600 9900
rect 15321 9863 15379 9869
rect 8602 9832 8608 9844
rect 6544 9804 7084 9832
rect 8252 9804 8608 9832
rect 6544 9792 6550 9804
rect 8252 9776 8280 9804
rect 8602 9792 8608 9804
rect 8660 9792 8666 9844
rect 8973 9835 9031 9841
rect 8973 9832 8985 9835
rect 8712 9804 8985 9832
rect 8234 9764 8240 9776
rect 4428 9736 4554 9764
rect 8195 9736 8240 9764
rect 4428 9724 4434 9736
rect 8234 9724 8240 9736
rect 8292 9724 8298 9776
rect 8510 9764 8516 9776
rect 8471 9736 8516 9764
rect 8510 9724 8516 9736
rect 8568 9764 8574 9776
rect 8712 9764 8740 9804
rect 8973 9801 8985 9804
rect 9019 9801 9031 9835
rect 9338 9832 9344 9844
rect 9299 9804 9344 9832
rect 8973 9795 9031 9801
rect 8878 9764 8884 9776
rect 8568 9736 8740 9764
rect 8839 9736 8884 9764
rect 8568 9724 8574 9736
rect 8878 9724 8884 9736
rect 8936 9724 8942 9776
rect 8988 9764 9016 9795
rect 9338 9792 9344 9804
rect 9396 9792 9402 9844
rect 12929 9835 12987 9841
rect 12929 9801 12941 9835
rect 12975 9832 12987 9835
rect 14214 9832 14220 9844
rect 12975 9804 14220 9832
rect 12975 9801 12987 9804
rect 12929 9795 12987 9801
rect 14214 9792 14220 9804
rect 14272 9792 14278 9844
rect 14306 9792 14312 9844
rect 14364 9832 14370 9844
rect 15336 9832 15364 9863
rect 15594 9860 15600 9872
rect 15652 9860 15658 9912
rect 15686 9860 15692 9912
rect 15744 9900 15750 9912
rect 15965 9903 16023 9909
rect 15965 9900 15977 9903
rect 15744 9872 15977 9900
rect 15744 9860 15750 9872
rect 15965 9869 15977 9872
rect 16011 9900 16023 9903
rect 16348 9900 16376 9940
rect 18633 9937 18645 9940
rect 18679 9937 18691 9971
rect 18633 9931 18691 9937
rect 19093 9971 19151 9977
rect 19093 9937 19105 9971
rect 19139 9937 19151 9971
rect 19093 9931 19151 9937
rect 19844 9940 20056 9968
rect 16011 9872 16376 9900
rect 17713 9903 17771 9909
rect 16011 9869 16023 9872
rect 15965 9863 16023 9869
rect 17713 9869 17725 9903
rect 17759 9900 17771 9903
rect 17805 9903 17863 9909
rect 17805 9900 17817 9903
rect 17759 9872 17817 9900
rect 17759 9869 17771 9872
rect 17713 9863 17771 9869
rect 17805 9869 17817 9872
rect 17851 9869 17863 9903
rect 17805 9863 17863 9869
rect 19274 9860 19280 9912
rect 19332 9900 19338 9912
rect 19553 9903 19611 9909
rect 19553 9900 19565 9903
rect 19332 9872 19565 9900
rect 19332 9860 19338 9872
rect 19553 9869 19565 9872
rect 19599 9869 19611 9903
rect 19734 9900 19740 9912
rect 19695 9872 19740 9900
rect 19553 9863 19611 9869
rect 19734 9860 19740 9872
rect 19792 9860 19798 9912
rect 19090 9832 19096 9844
rect 14364 9804 19096 9832
rect 14364 9792 14370 9804
rect 19090 9792 19096 9804
rect 19148 9832 19154 9844
rect 19844 9832 19872 9940
rect 20028 9909 20056 9940
rect 20286 9928 20292 9980
rect 20344 9968 20350 9980
rect 20381 9971 20439 9977
rect 20381 9968 20393 9971
rect 20344 9940 20393 9968
rect 20344 9928 20350 9940
rect 20381 9937 20393 9940
rect 20427 9968 20439 9971
rect 22218 9968 22224 9980
rect 20427 9940 22224 9968
rect 20427 9937 20439 9940
rect 20381 9931 20439 9937
rect 22218 9928 22224 9940
rect 22276 9928 22282 9980
rect 23892 9968 23920 10064
rect 23800 9940 23920 9968
rect 20013 9903 20071 9909
rect 20013 9869 20025 9903
rect 20059 9900 20071 9903
rect 20470 9900 20476 9912
rect 20059 9872 20476 9900
rect 20059 9869 20071 9872
rect 20013 9863 20071 9869
rect 20470 9860 20476 9872
rect 20528 9860 20534 9912
rect 23800 9909 23828 9940
rect 24058 9928 24064 9980
rect 24116 9968 24122 9980
rect 25438 9968 25444 9980
rect 24116 9940 25444 9968
rect 24116 9928 24122 9940
rect 25438 9928 25444 9940
rect 25496 9968 25502 9980
rect 25809 9971 25867 9977
rect 25809 9968 25821 9971
rect 25496 9940 25821 9968
rect 25496 9928 25502 9940
rect 25809 9937 25821 9940
rect 25855 9937 25867 9971
rect 25809 9931 25867 9937
rect 20565 9903 20623 9909
rect 20565 9869 20577 9903
rect 20611 9869 20623 9903
rect 20565 9863 20623 9869
rect 21117 9903 21175 9909
rect 21117 9869 21129 9903
rect 21163 9900 21175 9903
rect 23785 9903 23843 9909
rect 23785 9900 23797 9903
rect 21163 9872 23797 9900
rect 21163 9869 21175 9872
rect 21117 9863 21175 9869
rect 23785 9869 23797 9872
rect 23831 9869 23843 9903
rect 23785 9863 23843 9869
rect 19148 9804 19872 9832
rect 20580 9832 20608 9863
rect 21298 9832 21304 9844
rect 20580 9804 21304 9832
rect 19148 9792 19154 9804
rect 9430 9764 9436 9776
rect 8988 9736 9436 9764
rect 9430 9724 9436 9736
rect 9488 9724 9494 9776
rect 13386 9724 13392 9776
rect 13444 9764 13450 9776
rect 13573 9767 13631 9773
rect 13573 9764 13585 9767
rect 13444 9736 13585 9764
rect 13444 9724 13450 9736
rect 13573 9733 13585 9736
rect 13619 9733 13631 9767
rect 13573 9727 13631 9733
rect 14125 9767 14183 9773
rect 14125 9733 14137 9767
rect 14171 9764 14183 9767
rect 15686 9764 15692 9776
rect 14171 9736 15692 9764
rect 14171 9733 14183 9736
rect 14125 9727 14183 9733
rect 15686 9724 15692 9736
rect 15744 9724 15750 9776
rect 15778 9724 15784 9776
rect 15836 9764 15842 9776
rect 17342 9764 17348 9776
rect 15836 9736 17348 9764
rect 15836 9724 15842 9736
rect 17342 9724 17348 9736
rect 17400 9724 17406 9776
rect 17434 9724 17440 9776
rect 17492 9764 17498 9776
rect 17529 9767 17587 9773
rect 17529 9764 17541 9767
rect 17492 9736 17541 9764
rect 17492 9724 17498 9736
rect 17529 9733 17541 9736
rect 17575 9764 17587 9767
rect 17713 9767 17771 9773
rect 17713 9764 17725 9767
rect 17575 9736 17725 9764
rect 17575 9733 17587 9736
rect 17529 9727 17587 9733
rect 17713 9733 17725 9736
rect 17759 9764 17771 9767
rect 17986 9764 17992 9776
rect 17759 9736 17992 9764
rect 17759 9733 17771 9736
rect 17713 9727 17771 9733
rect 17986 9724 17992 9736
rect 18044 9764 18050 9776
rect 18265 9767 18323 9773
rect 18265 9764 18277 9767
rect 18044 9736 18277 9764
rect 18044 9724 18050 9736
rect 18265 9733 18277 9736
rect 18311 9733 18323 9767
rect 18265 9727 18323 9733
rect 18633 9767 18691 9773
rect 18633 9733 18645 9767
rect 18679 9764 18691 9767
rect 18817 9767 18875 9773
rect 18817 9764 18829 9767
rect 18679 9736 18829 9764
rect 18679 9733 18691 9736
rect 18633 9727 18691 9733
rect 18817 9733 18829 9736
rect 18863 9764 18875 9767
rect 20580 9764 20608 9804
rect 21298 9792 21304 9804
rect 21356 9792 21362 9844
rect 24061 9835 24119 9841
rect 24061 9832 24073 9835
rect 23616 9804 24073 9832
rect 23616 9776 23644 9804
rect 24061 9801 24073 9804
rect 24107 9801 24119 9835
rect 24061 9795 24119 9801
rect 24702 9792 24708 9844
rect 24760 9792 24766 9844
rect 18863 9736 20608 9764
rect 18863 9733 18875 9736
rect 18817 9727 18875 9733
rect 22218 9724 22224 9776
rect 22276 9764 22282 9776
rect 23046 9764 23052 9776
rect 22276 9736 23052 9764
rect 22276 9724 22282 9736
rect 23046 9724 23052 9736
rect 23104 9724 23110 9776
rect 23598 9764 23604 9776
rect 23559 9736 23604 9764
rect 23598 9724 23604 9736
rect 23656 9724 23662 9776
rect 400 9674 27264 9696
rect 400 9622 18870 9674
rect 18922 9622 18934 9674
rect 18986 9622 18998 9674
rect 19050 9622 19062 9674
rect 19114 9622 19126 9674
rect 19178 9622 27264 9674
rect 400 9600 27264 9622
rect 506 9520 512 9572
rect 564 9560 570 9572
rect 693 9563 751 9569
rect 693 9560 705 9563
rect 564 9532 705 9560
rect 564 9520 570 9532
rect 693 9529 705 9532
rect 739 9529 751 9563
rect 693 9523 751 9529
rect 708 9492 736 9523
rect 782 9520 788 9572
rect 840 9560 846 9572
rect 969 9563 1027 9569
rect 969 9560 981 9563
rect 840 9532 981 9560
rect 840 9520 846 9532
rect 969 9529 981 9532
rect 1015 9560 1027 9563
rect 1794 9560 1800 9572
rect 1015 9532 1800 9560
rect 1015 9529 1027 9532
rect 969 9523 1027 9529
rect 1794 9520 1800 9532
rect 1852 9520 1858 9572
rect 2070 9560 2076 9572
rect 1904 9532 2076 9560
rect 1610 9492 1616 9504
rect 708 9464 1616 9492
rect 1610 9452 1616 9464
rect 1668 9452 1674 9504
rect 1904 9501 1932 9532
rect 2070 9520 2076 9532
rect 2128 9520 2134 9572
rect 3266 9520 3272 9572
rect 3324 9560 3330 9572
rect 3324 9532 6164 9560
rect 3324 9520 3330 9532
rect 1889 9495 1947 9501
rect 1889 9461 1901 9495
rect 1935 9461 1947 9495
rect 1889 9455 1947 9461
rect 3174 9452 3180 9504
rect 3232 9492 3238 9504
rect 5198 9492 5204 9504
rect 3232 9464 5204 9492
rect 3232 9452 3238 9464
rect 5198 9452 5204 9464
rect 5256 9452 5262 9504
rect 6136 9501 6164 9532
rect 7406 9520 7412 9572
rect 7464 9560 7470 9572
rect 8605 9563 8663 9569
rect 8605 9560 8617 9563
rect 7464 9532 8617 9560
rect 7464 9520 7470 9532
rect 8605 9529 8617 9532
rect 8651 9560 8663 9563
rect 9338 9560 9344 9572
rect 8651 9532 9344 9560
rect 8651 9529 8663 9532
rect 8605 9523 8663 9529
rect 9338 9520 9344 9532
rect 9396 9520 9402 9572
rect 12558 9560 12564 9572
rect 12519 9532 12564 9560
rect 12558 9520 12564 9532
rect 12616 9520 12622 9572
rect 15318 9520 15324 9572
rect 15376 9560 15382 9572
rect 15413 9563 15471 9569
rect 15413 9560 15425 9563
rect 15376 9532 15425 9560
rect 15376 9520 15382 9532
rect 15413 9529 15425 9532
rect 15459 9529 15471 9563
rect 15413 9523 15471 9529
rect 17437 9563 17495 9569
rect 17437 9529 17449 9563
rect 17483 9560 17495 9563
rect 18078 9560 18084 9572
rect 17483 9532 18084 9560
rect 17483 9529 17495 9532
rect 17437 9523 17495 9529
rect 18078 9520 18084 9532
rect 18136 9520 18142 9572
rect 19461 9563 19519 9569
rect 19461 9560 19473 9563
rect 19292 9532 19473 9560
rect 19292 9504 19320 9532
rect 19461 9529 19473 9532
rect 19507 9560 19519 9563
rect 19734 9560 19740 9572
rect 19507 9532 19740 9560
rect 19507 9529 19519 9532
rect 19461 9523 19519 9529
rect 19734 9520 19740 9532
rect 19792 9520 19798 9572
rect 20286 9560 20292 9572
rect 20247 9532 20292 9560
rect 20286 9520 20292 9532
rect 20344 9520 20350 9572
rect 23782 9520 23788 9572
rect 23840 9560 23846 9572
rect 24521 9563 24579 9569
rect 24521 9560 24533 9563
rect 23840 9532 24533 9560
rect 23840 9520 23846 9532
rect 24521 9529 24533 9532
rect 24567 9529 24579 9563
rect 24702 9560 24708 9572
rect 24663 9532 24708 9560
rect 24521 9523 24579 9529
rect 6121 9495 6179 9501
rect 6121 9461 6133 9495
rect 6167 9492 6179 9495
rect 6394 9492 6400 9504
rect 6167 9464 6400 9492
rect 6167 9461 6179 9464
rect 6121 9455 6179 9461
rect 6394 9452 6400 9464
rect 6452 9452 6458 9504
rect 14398 9492 14404 9504
rect 13312 9464 14404 9492
rect 13312 9436 13340 9464
rect 14398 9452 14404 9464
rect 14456 9492 14462 9504
rect 15594 9492 15600 9504
rect 14456 9464 15600 9492
rect 14456 9452 14462 9464
rect 15594 9452 15600 9464
rect 15652 9452 15658 9504
rect 19274 9492 19280 9504
rect 19187 9464 19280 9492
rect 19274 9452 19280 9464
rect 19332 9452 19338 9504
rect 23046 9452 23052 9504
rect 23104 9492 23110 9504
rect 24536 9492 24564 9523
rect 24702 9520 24708 9532
rect 24760 9520 24766 9572
rect 25070 9492 25076 9504
rect 23104 9464 23874 9492
rect 24536 9464 25076 9492
rect 23104 9452 23110 9464
rect 2073 9427 2131 9433
rect 2073 9393 2085 9427
rect 2119 9424 2131 9427
rect 2346 9424 2352 9436
rect 2119 9396 2352 9424
rect 2119 9393 2131 9396
rect 2073 9387 2131 9393
rect 2346 9384 2352 9396
rect 2404 9384 2410 9436
rect 3358 9384 3364 9436
rect 3416 9424 3422 9436
rect 3821 9427 3879 9433
rect 3821 9424 3833 9427
rect 3416 9396 3833 9424
rect 3416 9384 3422 9396
rect 3821 9393 3833 9396
rect 3867 9393 3879 9427
rect 3821 9387 3879 9393
rect 4186 9384 4192 9436
rect 4244 9424 4250 9436
rect 4281 9427 4339 9433
rect 4281 9424 4293 9427
rect 4244 9396 4293 9424
rect 4244 9384 4250 9396
rect 4281 9393 4293 9396
rect 4327 9393 4339 9427
rect 4281 9387 4339 9393
rect 4554 9384 4560 9436
rect 4612 9424 4618 9436
rect 4741 9427 4799 9433
rect 4612 9396 4657 9424
rect 4612 9384 4618 9396
rect 4741 9393 4753 9427
rect 4787 9424 4799 9427
rect 6670 9424 6676 9436
rect 4787 9396 6676 9424
rect 4787 9393 4799 9396
rect 4741 9387 4799 9393
rect 2441 9359 2499 9365
rect 2441 9325 2453 9359
rect 2487 9356 2499 9359
rect 2530 9356 2536 9368
rect 2487 9328 2536 9356
rect 2487 9325 2499 9328
rect 2441 9319 2499 9325
rect 2530 9316 2536 9328
rect 2588 9316 2594 9368
rect 2990 9316 2996 9368
rect 3048 9356 3054 9368
rect 4756 9356 4784 9387
rect 6670 9384 6676 9396
rect 6728 9384 6734 9436
rect 6946 9424 6952 9436
rect 6907 9396 6952 9424
rect 6946 9384 6952 9396
rect 7004 9384 7010 9436
rect 9062 9424 9068 9436
rect 9023 9396 9068 9424
rect 9062 9384 9068 9396
rect 9120 9384 9126 9436
rect 11178 9424 11184 9436
rect 11139 9396 11184 9424
rect 11178 9384 11184 9396
rect 11236 9384 11242 9436
rect 12466 9424 12472 9436
rect 12427 9396 12472 9424
rect 12466 9384 12472 9396
rect 12524 9424 12530 9436
rect 13294 9424 13300 9436
rect 12524 9396 13300 9424
rect 12524 9384 12530 9396
rect 13294 9384 13300 9396
rect 13352 9384 13358 9436
rect 14122 9384 14128 9436
rect 14180 9424 14186 9436
rect 14677 9427 14735 9433
rect 14677 9424 14689 9427
rect 14180 9396 14689 9424
rect 14180 9384 14186 9396
rect 14677 9393 14689 9396
rect 14723 9424 14735 9427
rect 14766 9424 14772 9436
rect 14723 9396 14772 9424
rect 14723 9393 14735 9396
rect 14677 9387 14735 9393
rect 14766 9384 14772 9396
rect 14824 9384 14830 9436
rect 16422 9384 16428 9436
rect 16480 9424 16486 9436
rect 16609 9427 16667 9433
rect 16609 9424 16621 9427
rect 16480 9396 16621 9424
rect 16480 9384 16486 9396
rect 16609 9393 16621 9396
rect 16655 9424 16667 9427
rect 17710 9424 17716 9436
rect 16655 9396 17716 9424
rect 16655 9393 16667 9396
rect 16609 9387 16667 9393
rect 17710 9384 17716 9396
rect 17768 9384 17774 9436
rect 18722 9424 18728 9436
rect 18683 9396 18728 9424
rect 18722 9384 18728 9396
rect 18780 9384 18786 9436
rect 18906 9424 18912 9436
rect 18819 9396 18912 9424
rect 18906 9384 18912 9396
rect 18964 9424 18970 9436
rect 19366 9424 19372 9436
rect 18964 9396 19372 9424
rect 18964 9384 18970 9396
rect 19366 9384 19372 9396
rect 19424 9384 19430 9436
rect 23414 9424 23420 9436
rect 23375 9396 23420 9424
rect 23414 9384 23420 9396
rect 23472 9384 23478 9436
rect 23690 9424 23696 9436
rect 23651 9396 23696 9424
rect 23690 9384 23696 9396
rect 23748 9384 23754 9436
rect 23846 9424 23874 9464
rect 25070 9452 25076 9464
rect 25128 9452 25134 9504
rect 24150 9424 24156 9436
rect 23846 9396 24156 9424
rect 24150 9384 24156 9396
rect 24208 9384 24214 9436
rect 5106 9356 5112 9368
rect 3048 9328 4784 9356
rect 5067 9328 5112 9356
rect 3048 9316 3054 9328
rect 5106 9316 5112 9328
rect 5164 9316 5170 9368
rect 5201 9359 5259 9365
rect 5201 9325 5213 9359
rect 5247 9325 5259 9359
rect 5201 9319 5259 9325
rect 3910 9248 3916 9300
rect 3968 9288 3974 9300
rect 4370 9288 4376 9300
rect 3968 9260 4376 9288
rect 3968 9248 3974 9260
rect 4370 9248 4376 9260
rect 4428 9288 4434 9300
rect 4428 9260 4968 9288
rect 4428 9248 4434 9260
rect 4940 9232 4968 9260
rect 3082 9180 3088 9232
rect 3140 9220 3146 9232
rect 4278 9220 4284 9232
rect 3140 9192 4284 9220
rect 3140 9180 3146 9192
rect 4278 9180 4284 9192
rect 4336 9180 4342 9232
rect 4922 9180 4928 9232
rect 4980 9220 4986 9232
rect 5216 9220 5244 9319
rect 6762 9316 6768 9368
rect 6820 9356 6826 9368
rect 7130 9356 7136 9368
rect 6820 9328 7136 9356
rect 6820 9316 6826 9328
rect 7130 9316 7136 9328
rect 7188 9316 7194 9368
rect 8973 9359 9031 9365
rect 8973 9325 8985 9359
rect 9019 9325 9031 9359
rect 11086 9356 11092 9368
rect 11047 9328 11092 9356
rect 8973 9319 9031 9325
rect 6670 9248 6676 9300
rect 6728 9288 6734 9300
rect 8602 9288 8608 9300
rect 6728 9260 8608 9288
rect 6728 9248 6734 9260
rect 8602 9248 8608 9260
rect 8660 9288 8666 9300
rect 8988 9288 9016 9319
rect 11086 9316 11092 9328
rect 11144 9316 11150 9368
rect 13846 9316 13852 9368
rect 13904 9356 13910 9368
rect 14585 9359 14643 9365
rect 14585 9356 14597 9359
rect 13904 9328 14597 9356
rect 13904 9316 13910 9328
rect 14585 9325 14597 9328
rect 14631 9356 14643 9359
rect 15318 9356 15324 9368
rect 14631 9328 15324 9356
rect 14631 9325 14643 9328
rect 14585 9319 14643 9325
rect 15318 9316 15324 9328
rect 15376 9356 15382 9368
rect 15376 9328 16468 9356
rect 15376 9316 15382 9328
rect 9338 9288 9344 9300
rect 8660 9260 9344 9288
rect 8660 9248 8666 9260
rect 9338 9248 9344 9260
rect 9396 9248 9402 9300
rect 16440 9297 16468 9328
rect 23322 9316 23328 9368
rect 23380 9356 23386 9368
rect 24337 9359 24395 9365
rect 24337 9356 24349 9359
rect 23380 9328 24349 9356
rect 23380 9316 23386 9328
rect 24337 9325 24349 9328
rect 24383 9356 24395 9359
rect 25162 9356 25168 9368
rect 24383 9328 25168 9356
rect 24383 9325 24395 9328
rect 24337 9319 24395 9325
rect 25162 9316 25168 9328
rect 25220 9316 25226 9368
rect 16425 9291 16483 9297
rect 16425 9257 16437 9291
rect 16471 9288 16483 9291
rect 16514 9288 16520 9300
rect 16471 9260 16520 9288
rect 16471 9257 16483 9260
rect 16425 9251 16483 9257
rect 16514 9248 16520 9260
rect 16572 9248 16578 9300
rect 23046 9248 23052 9300
rect 23104 9288 23110 9300
rect 23417 9291 23475 9297
rect 23417 9288 23429 9291
rect 23104 9260 23429 9288
rect 23104 9248 23110 9260
rect 23417 9257 23429 9260
rect 23463 9288 23475 9291
rect 23598 9288 23604 9300
rect 23463 9260 23604 9288
rect 23463 9257 23475 9260
rect 23417 9251 23475 9257
rect 23598 9248 23604 9260
rect 23656 9248 23662 9300
rect 6578 9220 6584 9232
rect 4980 9192 6584 9220
rect 4980 9180 4986 9192
rect 6578 9180 6584 9192
rect 6636 9220 6642 9232
rect 7866 9220 7872 9232
rect 6636 9192 7872 9220
rect 6636 9180 6642 9192
rect 7866 9180 7872 9192
rect 7924 9220 7930 9232
rect 9246 9220 9252 9232
rect 7924 9192 9252 9220
rect 7924 9180 7930 9192
rect 9246 9180 9252 9192
rect 9304 9180 9310 9232
rect 11270 9180 11276 9232
rect 11328 9220 11334 9232
rect 11365 9223 11423 9229
rect 11365 9220 11377 9223
rect 11328 9192 11377 9220
rect 11328 9180 11334 9192
rect 11365 9189 11377 9192
rect 11411 9189 11423 9223
rect 14858 9220 14864 9232
rect 14819 9192 14864 9220
rect 11365 9183 11423 9189
rect 14858 9180 14864 9192
rect 14916 9180 14922 9232
rect 15226 9220 15232 9232
rect 15187 9192 15232 9220
rect 15226 9180 15232 9192
rect 15284 9180 15290 9232
rect 22770 9180 22776 9232
rect 22828 9220 22834 9232
rect 23690 9220 23696 9232
rect 22828 9192 23696 9220
rect 22828 9180 22834 9192
rect 23690 9180 23696 9192
rect 23748 9180 23754 9232
rect 400 9130 27264 9152
rect 400 9078 3510 9130
rect 3562 9078 3574 9130
rect 3626 9078 3638 9130
rect 3690 9078 3702 9130
rect 3754 9078 3766 9130
rect 3818 9078 27264 9130
rect 400 9056 27264 9078
rect 2070 9016 2076 9028
rect 2031 8988 2076 9016
rect 2070 8976 2076 8988
rect 2128 8976 2134 9028
rect 2990 9016 2996 9028
rect 2951 8988 2996 9016
rect 2990 8976 2996 8988
rect 3048 8976 3054 9028
rect 3174 9016 3180 9028
rect 3135 8988 3180 9016
rect 3174 8976 3180 8988
rect 3232 8976 3238 9028
rect 3545 9019 3603 9025
rect 3545 8985 3557 9019
rect 3591 9016 3603 9019
rect 3910 9016 3916 9028
rect 3591 8988 3916 9016
rect 3591 8985 3603 8988
rect 3545 8979 3603 8985
rect 3910 8976 3916 8988
rect 3968 8976 3974 9028
rect 4278 8976 4284 9028
rect 4336 9016 4342 9028
rect 4922 9016 4928 9028
rect 4336 8988 4381 9016
rect 4883 8988 4928 9016
rect 4336 8976 4342 8988
rect 4922 8976 4928 8988
rect 4980 8976 4986 9028
rect 5569 9019 5627 9025
rect 5569 8985 5581 9019
rect 5615 9016 5627 9019
rect 6946 9016 6952 9028
rect 5615 8988 6952 9016
rect 5615 8985 5627 8988
rect 5569 8979 5627 8985
rect 6946 8976 6952 8988
rect 7004 9016 7010 9028
rect 7593 9019 7651 9025
rect 7593 9016 7605 9019
rect 7004 8988 7605 9016
rect 7004 8976 7010 8988
rect 7593 8985 7605 8988
rect 7639 9016 7651 9019
rect 8053 9019 8111 9025
rect 8053 9016 8065 9019
rect 7639 8988 8065 9016
rect 7639 8985 7651 8988
rect 7593 8979 7651 8985
rect 8053 8985 8065 8988
rect 8099 8985 8111 9019
rect 9062 9016 9068 9028
rect 9023 8988 9068 9016
rect 8053 8979 8111 8985
rect 9062 8976 9068 8988
rect 9120 8976 9126 9028
rect 9246 9016 9252 9028
rect 9207 8988 9252 9016
rect 9246 8976 9252 8988
rect 9304 8976 9310 9028
rect 9338 8976 9344 9028
rect 9396 9016 9402 9028
rect 9396 8988 9441 9016
rect 9396 8976 9402 8988
rect 11086 8976 11092 9028
rect 11144 9016 11150 9028
rect 11181 9019 11239 9025
rect 11181 9016 11193 9019
rect 11144 8988 11193 9016
rect 11144 8976 11150 8988
rect 11181 8985 11193 8988
rect 11227 9016 11239 9019
rect 11454 9016 11460 9028
rect 11227 8988 11460 9016
rect 11227 8985 11239 8988
rect 11181 8979 11239 8985
rect 11454 8976 11460 8988
rect 11512 9016 11518 9028
rect 12285 9019 12343 9025
rect 12285 9016 12297 9019
rect 11512 8988 12297 9016
rect 11512 8976 11518 8988
rect 12285 8985 12297 8988
rect 12331 9016 12343 9019
rect 12377 9019 12435 9025
rect 12377 9016 12389 9019
rect 12331 8988 12389 9016
rect 12331 8985 12343 8988
rect 12285 8979 12343 8985
rect 12377 8985 12389 8988
rect 12423 9016 12435 9019
rect 12558 9016 12564 9028
rect 12423 8988 12564 9016
rect 12423 8985 12435 8988
rect 12377 8979 12435 8985
rect 12558 8976 12564 8988
rect 12616 8976 12622 9028
rect 14858 9016 14864 9028
rect 13956 8988 14864 9016
rect 1981 8951 2039 8957
rect 1981 8917 1993 8951
rect 2027 8948 2039 8951
rect 2346 8948 2352 8960
rect 2027 8920 2352 8948
rect 2027 8917 2039 8920
rect 1981 8911 2039 8917
rect 2346 8908 2352 8920
rect 2404 8908 2410 8960
rect 3082 8908 3088 8960
rect 3140 8948 3146 8960
rect 3269 8951 3327 8957
rect 3269 8948 3281 8951
rect 3140 8920 3281 8948
rect 3140 8908 3146 8920
rect 3269 8917 3281 8920
rect 3315 8917 3327 8951
rect 3269 8911 3327 8917
rect 3729 8951 3787 8957
rect 3729 8917 3741 8951
rect 3775 8948 3787 8951
rect 4554 8948 4560 8960
rect 3775 8920 4560 8948
rect 3775 8917 3787 8920
rect 3729 8911 3787 8917
rect 4554 8908 4560 8920
rect 4612 8948 4618 8960
rect 5753 8951 5811 8957
rect 4612 8920 4705 8948
rect 4612 8908 4618 8920
rect 690 8840 696 8892
rect 748 8880 754 8892
rect 1705 8883 1763 8889
rect 1705 8880 1717 8883
rect 748 8852 1717 8880
rect 748 8840 754 8852
rect 1705 8849 1717 8852
rect 1751 8849 1763 8883
rect 1705 8843 1763 8849
rect 3913 8883 3971 8889
rect 3913 8849 3925 8883
rect 3959 8880 3971 8883
rect 4186 8880 4192 8892
rect 3959 8852 4192 8880
rect 3959 8849 3971 8852
rect 3913 8843 3971 8849
rect 4186 8840 4192 8852
rect 4244 8840 4250 8892
rect 4664 8880 4692 8920
rect 5753 8917 5765 8951
rect 5799 8948 5811 8951
rect 6762 8948 6768 8960
rect 5799 8920 6768 8948
rect 5799 8917 5811 8920
rect 5753 8911 5811 8917
rect 6762 8908 6768 8920
rect 6820 8908 6826 8960
rect 8878 8908 8884 8960
rect 8936 8948 8942 8960
rect 11825 8951 11883 8957
rect 11825 8948 11837 8951
rect 8936 8920 11837 8948
rect 8936 8908 8942 8920
rect 11825 8917 11837 8920
rect 11871 8948 11883 8951
rect 12466 8948 12472 8960
rect 11871 8920 12472 8948
rect 11871 8917 11883 8920
rect 11825 8911 11883 8917
rect 12466 8908 12472 8920
rect 12524 8908 12530 8960
rect 4664 8852 5980 8880
rect 782 8812 788 8824
rect 743 8784 788 8812
rect 782 8772 788 8784
rect 840 8772 846 8824
rect 1610 8812 1616 8824
rect 1571 8784 1616 8812
rect 1610 8772 1616 8784
rect 1668 8772 1674 8824
rect 4005 8815 4063 8821
rect 4005 8781 4017 8815
rect 4051 8781 4063 8815
rect 4005 8775 4063 8781
rect 4097 8815 4155 8821
rect 4097 8781 4109 8815
rect 4143 8812 4155 8815
rect 4370 8812 4376 8824
rect 4143 8784 4376 8812
rect 4143 8781 4155 8784
rect 4097 8775 4155 8781
rect 874 8744 880 8756
rect 835 8716 880 8744
rect 874 8704 880 8716
rect 932 8704 938 8756
rect 2349 8679 2407 8685
rect 2349 8645 2361 8679
rect 2395 8676 2407 8679
rect 2530 8676 2536 8688
rect 2395 8648 2536 8676
rect 2395 8645 2407 8648
rect 2349 8639 2407 8645
rect 2530 8636 2536 8648
rect 2588 8636 2594 8688
rect 4020 8676 4048 8775
rect 4370 8772 4376 8784
rect 4428 8772 4434 8824
rect 5952 8821 5980 8852
rect 6210 8840 6216 8892
rect 6268 8880 6274 8892
rect 6949 8883 7007 8889
rect 6949 8880 6961 8883
rect 6268 8852 6961 8880
rect 6268 8840 6274 8852
rect 6949 8849 6961 8852
rect 6995 8880 7007 8883
rect 8234 8880 8240 8892
rect 6995 8852 8240 8880
rect 6995 8849 7007 8852
rect 6949 8843 7007 8849
rect 7884 8821 7912 8852
rect 8234 8840 8240 8852
rect 8292 8880 8298 8892
rect 8605 8883 8663 8889
rect 8605 8880 8617 8883
rect 8292 8852 8617 8880
rect 8292 8840 8298 8852
rect 8605 8849 8617 8852
rect 8651 8880 8663 8883
rect 9062 8880 9068 8892
rect 8651 8852 9068 8880
rect 8651 8849 8663 8852
rect 8605 8843 8663 8849
rect 9062 8840 9068 8852
rect 9120 8840 9126 8892
rect 11178 8840 11184 8892
rect 11236 8880 11242 8892
rect 11457 8883 11515 8889
rect 11457 8880 11469 8883
rect 11236 8852 11469 8880
rect 11236 8840 11242 8852
rect 11457 8849 11469 8852
rect 11503 8849 11515 8883
rect 12576 8880 12604 8976
rect 13386 8948 13392 8960
rect 13347 8920 13392 8948
rect 13386 8908 13392 8920
rect 13444 8908 13450 8960
rect 12653 8883 12711 8889
rect 12653 8880 12665 8883
rect 12576 8852 12665 8880
rect 11457 8843 11515 8849
rect 12653 8849 12665 8852
rect 12699 8849 12711 8883
rect 12653 8843 12711 8849
rect 5937 8815 5995 8821
rect 5937 8781 5949 8815
rect 5983 8812 5995 8815
rect 7777 8815 7835 8821
rect 5983 8784 6532 8812
rect 5983 8781 5995 8784
rect 5937 8775 5995 8781
rect 6504 8756 6532 8784
rect 7777 8781 7789 8815
rect 7823 8781 7835 8815
rect 7777 8775 7835 8781
rect 7869 8815 7927 8821
rect 7869 8781 7881 8815
rect 7915 8781 7927 8815
rect 11270 8812 11276 8824
rect 11231 8784 11276 8812
rect 7869 8775 7927 8781
rect 4186 8704 4192 8756
rect 4244 8744 4250 8756
rect 6121 8747 6179 8753
rect 6121 8744 6133 8747
rect 4244 8716 6133 8744
rect 4244 8704 4250 8716
rect 6121 8713 6133 8716
rect 6167 8744 6179 8747
rect 6210 8744 6216 8756
rect 6167 8716 6216 8744
rect 6167 8713 6179 8716
rect 6121 8707 6179 8713
rect 6210 8704 6216 8716
rect 6268 8704 6274 8756
rect 6486 8744 6492 8756
rect 6447 8716 6492 8744
rect 6486 8704 6492 8716
rect 6544 8704 6550 8756
rect 6854 8744 6860 8756
rect 6815 8716 6860 8744
rect 6854 8704 6860 8716
rect 6912 8704 6918 8756
rect 7792 8744 7820 8775
rect 11270 8772 11276 8784
rect 11328 8772 11334 8824
rect 13110 8812 13116 8824
rect 13071 8784 13116 8812
rect 13110 8772 13116 8784
rect 13168 8772 13174 8824
rect 13389 8815 13447 8821
rect 13389 8781 13401 8815
rect 13435 8781 13447 8815
rect 13389 8775 13447 8781
rect 8510 8744 8516 8756
rect 7792 8716 8516 8744
rect 8510 8704 8516 8716
rect 8568 8744 8574 8756
rect 11362 8744 11368 8756
rect 8568 8716 11368 8744
rect 8568 8704 8574 8716
rect 11362 8704 11368 8716
rect 11420 8704 11426 8756
rect 12101 8747 12159 8753
rect 12101 8713 12113 8747
rect 12147 8744 12159 8747
rect 13018 8744 13024 8756
rect 12147 8716 13024 8744
rect 12147 8713 12159 8716
rect 12101 8707 12159 8713
rect 13018 8704 13024 8716
rect 13076 8744 13082 8756
rect 13404 8744 13432 8775
rect 13956 8753 13984 8988
rect 14858 8976 14864 8988
rect 14916 8976 14922 9028
rect 15318 9016 15324 9028
rect 15279 8988 15324 9016
rect 15318 8976 15324 8988
rect 15376 8976 15382 9028
rect 16422 9016 16428 9028
rect 16383 8988 16428 9016
rect 16422 8976 16428 8988
rect 16480 8976 16486 9028
rect 16514 8976 16520 9028
rect 16572 9016 16578 9028
rect 16572 8988 16617 9016
rect 16572 8976 16578 8988
rect 18722 8976 18728 9028
rect 18780 9016 18786 9028
rect 19093 9019 19151 9025
rect 19093 9016 19105 9019
rect 18780 8988 19105 9016
rect 18780 8976 18786 8988
rect 19093 8985 19105 8988
rect 19139 8985 19151 9019
rect 19274 9016 19280 9028
rect 19235 8988 19280 9016
rect 19093 8979 19151 8985
rect 19274 8976 19280 8988
rect 19332 8976 19338 9028
rect 20470 8976 20476 9028
rect 20528 9016 20534 9028
rect 21117 9019 21175 9025
rect 21117 9016 21129 9019
rect 20528 8988 21129 9016
rect 20528 8976 20534 8988
rect 21117 8985 21129 8988
rect 21163 9016 21175 9019
rect 21482 9016 21488 9028
rect 21163 8988 21488 9016
rect 21163 8985 21175 8988
rect 21117 8979 21175 8985
rect 21482 8976 21488 8988
rect 21540 9016 21546 9028
rect 21669 9019 21727 9025
rect 21669 9016 21681 9019
rect 21540 8988 21681 9016
rect 21540 8976 21546 8988
rect 21669 8985 21681 8988
rect 21715 8985 21727 9019
rect 22218 9016 22224 9028
rect 22179 8988 22224 9016
rect 21669 8979 21727 8985
rect 22218 8976 22224 8988
rect 22276 8976 22282 9028
rect 22589 9019 22647 9025
rect 22589 8985 22601 9019
rect 22635 9016 22647 9019
rect 22770 9016 22776 9028
rect 22635 8988 22776 9016
rect 22635 8985 22647 8988
rect 22589 8979 22647 8985
rect 22770 8976 22776 8988
rect 22828 8976 22834 9028
rect 23046 9016 23052 9028
rect 23007 8988 23052 9016
rect 23046 8976 23052 8988
rect 23104 8976 23110 9028
rect 23414 9016 23420 9028
rect 23375 8988 23420 9016
rect 23414 8976 23420 8988
rect 23472 9016 23478 9028
rect 24153 9019 24211 9025
rect 24153 9016 24165 9019
rect 23472 8988 24165 9016
rect 23472 8976 23478 8988
rect 24153 8985 24165 8988
rect 24199 9016 24211 9019
rect 24337 9019 24395 9025
rect 24337 9016 24349 9019
rect 24199 8988 24349 9016
rect 24199 8985 24211 8988
rect 24153 8979 24211 8985
rect 24337 8985 24349 8988
rect 24383 8985 24395 9019
rect 25438 9016 25444 9028
rect 25399 8988 25444 9016
rect 24337 8979 24395 8985
rect 25438 8976 25444 8988
rect 25496 8976 25502 9028
rect 14214 8908 14220 8960
rect 14272 8948 14278 8960
rect 17805 8951 17863 8957
rect 14272 8920 14317 8948
rect 14272 8908 14278 8920
rect 17805 8917 17817 8951
rect 17851 8948 17863 8951
rect 18906 8948 18912 8960
rect 17851 8920 18912 8948
rect 17851 8917 17863 8920
rect 17805 8911 17863 8917
rect 18906 8908 18912 8920
rect 18964 8908 18970 8960
rect 14232 8880 14260 8908
rect 14953 8883 15011 8889
rect 14953 8880 14965 8883
rect 14232 8852 14965 8880
rect 14953 8849 14965 8852
rect 14999 8880 15011 8883
rect 15226 8880 15232 8892
rect 14999 8852 15232 8880
rect 14999 8849 15011 8852
rect 14953 8843 15011 8849
rect 15226 8840 15232 8852
rect 15284 8840 15290 8892
rect 18262 8880 18268 8892
rect 17912 8852 18268 8880
rect 14674 8812 14680 8824
rect 14587 8784 14680 8812
rect 14674 8772 14680 8784
rect 14732 8812 14738 8824
rect 15137 8815 15195 8821
rect 15137 8812 15149 8815
rect 14732 8784 15149 8812
rect 14732 8772 14738 8784
rect 15137 8781 15149 8784
rect 15183 8781 15195 8815
rect 15137 8775 15195 8781
rect 16514 8772 16520 8824
rect 16572 8812 16578 8824
rect 17710 8812 17716 8824
rect 16572 8784 17716 8812
rect 16572 8772 16578 8784
rect 17710 8772 17716 8784
rect 17768 8812 17774 8824
rect 17912 8821 17940 8852
rect 18262 8840 18268 8852
rect 18320 8840 18326 8892
rect 17897 8815 17955 8821
rect 17897 8812 17909 8815
rect 17768 8784 17909 8812
rect 17768 8772 17774 8784
rect 17897 8781 17909 8784
rect 17943 8781 17955 8815
rect 17897 8775 17955 8781
rect 18081 8815 18139 8821
rect 18081 8781 18093 8815
rect 18127 8812 18139 8815
rect 18127 8784 18308 8812
rect 18127 8781 18139 8784
rect 18081 8775 18139 8781
rect 13941 8747 13999 8753
rect 13941 8744 13953 8747
rect 13076 8716 13953 8744
rect 13076 8704 13082 8716
rect 13941 8713 13953 8716
rect 13987 8713 13999 8747
rect 13941 8707 13999 8713
rect 14401 8747 14459 8753
rect 14401 8713 14413 8747
rect 14447 8744 14459 8747
rect 14490 8744 14496 8756
rect 14447 8716 14496 8744
rect 14447 8713 14459 8716
rect 14401 8707 14459 8713
rect 14490 8704 14496 8716
rect 14548 8704 14554 8756
rect 18280 8688 18308 8784
rect 18446 8772 18452 8824
rect 18504 8812 18510 8824
rect 18924 8812 18952 8908
rect 22788 8880 22816 8976
rect 23306 8951 23364 8957
rect 23306 8917 23318 8951
rect 23352 8917 23364 8951
rect 23306 8911 23364 8917
rect 23321 8880 23349 8911
rect 22788 8852 23349 8880
rect 23509 8883 23567 8889
rect 23509 8849 23521 8883
rect 23555 8849 23567 8883
rect 23509 8843 23567 8849
rect 23877 8883 23935 8889
rect 23877 8849 23889 8883
rect 23923 8880 23935 8883
rect 24521 8883 24579 8889
rect 24521 8880 24533 8883
rect 23923 8852 24533 8880
rect 23923 8849 23935 8852
rect 23877 8843 23935 8849
rect 21298 8812 21304 8824
rect 18504 8784 18952 8812
rect 21211 8784 21304 8812
rect 18504 8772 18510 8784
rect 21298 8772 21304 8784
rect 21356 8812 21362 8824
rect 22405 8815 22463 8821
rect 21356 8784 21620 8812
rect 21356 8772 21362 8784
rect 18354 8704 18360 8756
rect 18412 8744 18418 8756
rect 18725 8747 18783 8753
rect 18725 8744 18737 8747
rect 18412 8716 18737 8744
rect 18412 8704 18418 8716
rect 18725 8713 18737 8716
rect 18771 8713 18783 8747
rect 18725 8707 18783 8713
rect 4738 8676 4744 8688
rect 4020 8648 4744 8676
rect 4738 8636 4744 8648
rect 4796 8636 4802 8688
rect 5385 8679 5443 8685
rect 5385 8645 5397 8679
rect 5431 8676 5443 8679
rect 6302 8676 6308 8688
rect 5431 8648 6308 8676
rect 5431 8645 5443 8648
rect 5385 8639 5443 8645
rect 6302 8636 6308 8648
rect 6360 8636 6366 8688
rect 6397 8679 6455 8685
rect 6397 8645 6409 8679
rect 6443 8676 6455 8679
rect 6670 8676 6676 8688
rect 6443 8648 6676 8676
rect 6443 8645 6455 8648
rect 6397 8639 6455 8645
rect 6670 8636 6676 8648
rect 6728 8676 6734 8688
rect 7133 8679 7191 8685
rect 7133 8676 7145 8679
rect 6728 8648 7145 8676
rect 6728 8636 6734 8648
rect 7133 8645 7145 8648
rect 7179 8645 7191 8679
rect 7133 8639 7191 8645
rect 18262 8636 18268 8688
rect 18320 8676 18326 8688
rect 21592 8685 21620 8784
rect 22405 8781 22417 8815
rect 22451 8812 22463 8815
rect 23141 8815 23199 8821
rect 23141 8812 23153 8815
rect 22451 8784 23153 8812
rect 22451 8781 22463 8784
rect 22405 8775 22463 8781
rect 23141 8781 23153 8784
rect 23187 8812 23199 8815
rect 23322 8812 23328 8824
rect 23187 8784 23328 8812
rect 23187 8781 23199 8784
rect 23141 8775 23199 8781
rect 23322 8772 23328 8784
rect 23380 8772 23386 8824
rect 23524 8756 23552 8843
rect 23969 8815 24027 8821
rect 23969 8812 23981 8815
rect 23846 8784 23981 8812
rect 23506 8704 23512 8756
rect 23564 8744 23570 8756
rect 23846 8744 23874 8784
rect 23969 8781 23981 8784
rect 24015 8781 24027 8815
rect 23969 8775 24027 8781
rect 23564 8716 23874 8744
rect 23564 8704 23570 8716
rect 18541 8679 18599 8685
rect 18541 8676 18553 8679
rect 18320 8648 18553 8676
rect 18320 8636 18326 8648
rect 18541 8645 18553 8648
rect 18587 8645 18599 8679
rect 18541 8639 18599 8645
rect 21577 8679 21635 8685
rect 21577 8645 21589 8679
rect 21623 8676 21635 8679
rect 24076 8676 24104 8852
rect 24521 8849 24533 8852
rect 24567 8849 24579 8883
rect 25162 8880 25168 8892
rect 25075 8852 25168 8880
rect 24521 8843 24579 8849
rect 25162 8840 25168 8852
rect 25220 8880 25226 8892
rect 25257 8883 25315 8889
rect 25257 8880 25269 8883
rect 25220 8852 25269 8880
rect 25220 8840 25226 8852
rect 25257 8849 25269 8852
rect 25303 8849 25315 8883
rect 25257 8843 25315 8849
rect 25073 8815 25131 8821
rect 25073 8781 25085 8815
rect 25119 8812 25131 8815
rect 25438 8812 25444 8824
rect 25119 8784 25444 8812
rect 25119 8781 25131 8784
rect 25073 8775 25131 8781
rect 25438 8772 25444 8784
rect 25496 8772 25502 8824
rect 21623 8648 24104 8676
rect 21623 8645 21635 8648
rect 21577 8639 21635 8645
rect 400 8586 27264 8608
rect 400 8534 18870 8586
rect 18922 8534 18934 8586
rect 18986 8534 18998 8586
rect 19050 8534 19062 8586
rect 19114 8534 19126 8586
rect 19178 8534 27264 8586
rect 400 8512 27264 8534
rect 690 8472 696 8484
rect 651 8444 696 8472
rect 690 8432 696 8444
rect 748 8432 754 8484
rect 874 8472 880 8484
rect 835 8444 880 8472
rect 874 8432 880 8444
rect 932 8432 938 8484
rect 3358 8432 3364 8484
rect 3416 8472 3422 8484
rect 3821 8475 3879 8481
rect 3821 8472 3833 8475
rect 3416 8444 3833 8472
rect 3416 8432 3422 8444
rect 3821 8441 3833 8444
rect 3867 8441 3879 8475
rect 4646 8472 4652 8484
rect 3821 8435 3879 8441
rect 4526 8444 4652 8472
rect 4097 8407 4155 8413
rect 4097 8373 4109 8407
rect 4143 8404 4155 8407
rect 4370 8404 4376 8416
rect 4143 8376 4376 8404
rect 4143 8373 4155 8376
rect 4097 8367 4155 8373
rect 4370 8364 4376 8376
rect 4428 8404 4434 8416
rect 4526 8404 4554 8444
rect 4646 8432 4652 8444
rect 4704 8432 4710 8484
rect 5290 8432 5296 8484
rect 5348 8472 5354 8484
rect 6213 8475 6271 8481
rect 6213 8472 6225 8475
rect 5348 8444 6225 8472
rect 5348 8432 5354 8444
rect 6213 8441 6225 8444
rect 6259 8472 6271 8475
rect 6854 8472 6860 8484
rect 6259 8444 6860 8472
rect 6259 8441 6271 8444
rect 6213 8435 6271 8441
rect 6854 8432 6860 8444
rect 6912 8432 6918 8484
rect 9062 8472 9068 8484
rect 9023 8444 9068 8472
rect 9062 8432 9068 8444
rect 9120 8432 9126 8484
rect 12837 8475 12895 8481
rect 12837 8441 12849 8475
rect 12883 8472 12895 8475
rect 13386 8472 13392 8484
rect 12883 8444 13392 8472
rect 12883 8441 12895 8444
rect 12837 8435 12895 8441
rect 13386 8432 13392 8444
rect 13444 8432 13450 8484
rect 14677 8475 14735 8481
rect 14677 8441 14689 8475
rect 14723 8472 14735 8475
rect 14766 8472 14772 8484
rect 14723 8444 14772 8472
rect 14723 8441 14735 8444
rect 14677 8435 14735 8441
rect 14766 8432 14772 8444
rect 14824 8432 14830 8484
rect 23141 8475 23199 8481
rect 23141 8441 23153 8475
rect 23187 8472 23199 8475
rect 23322 8472 23328 8484
rect 23187 8444 23328 8472
rect 23187 8441 23199 8444
rect 23141 8435 23199 8441
rect 23322 8432 23328 8444
rect 23380 8432 23386 8484
rect 6394 8404 6400 8416
rect 4428 8376 4554 8404
rect 6355 8376 6400 8404
rect 4428 8364 4434 8376
rect 6394 8364 6400 8376
rect 6452 8364 6458 8416
rect 6670 8404 6676 8416
rect 6631 8376 6676 8404
rect 6670 8364 6676 8376
rect 6728 8364 6734 8416
rect 11273 8407 11331 8413
rect 11273 8373 11285 8407
rect 11319 8404 11331 8407
rect 11362 8404 11368 8416
rect 11319 8376 11368 8404
rect 11319 8373 11331 8376
rect 11273 8367 11331 8373
rect 11362 8364 11368 8376
rect 11420 8364 11426 8416
rect 11825 8407 11883 8413
rect 11825 8373 11837 8407
rect 11871 8404 11883 8407
rect 12006 8404 12012 8416
rect 11871 8376 12012 8404
rect 11871 8373 11883 8376
rect 11825 8367 11883 8373
rect 12006 8364 12012 8376
rect 12064 8364 12070 8416
rect 1429 8339 1487 8345
rect 1429 8305 1441 8339
rect 1475 8336 1487 8339
rect 1518 8336 1524 8348
rect 1475 8308 1524 8336
rect 1475 8305 1487 8308
rect 1429 8299 1487 8305
rect 1518 8296 1524 8308
rect 1576 8296 1582 8348
rect 1610 8296 1616 8348
rect 1668 8336 1674 8348
rect 4002 8336 4008 8348
rect 1668 8308 4008 8336
rect 1668 8296 1674 8308
rect 4002 8296 4008 8308
rect 4060 8296 4066 8348
rect 4186 8296 4192 8348
rect 4244 8336 4250 8348
rect 4281 8339 4339 8345
rect 4281 8336 4293 8339
rect 4244 8308 4293 8336
rect 4244 8296 4250 8308
rect 4281 8305 4293 8308
rect 4327 8305 4339 8339
rect 4281 8299 4339 8305
rect 4649 8339 4707 8345
rect 4649 8305 4661 8339
rect 4695 8336 4707 8339
rect 4738 8336 4744 8348
rect 4695 8308 4744 8336
rect 4695 8305 4707 8308
rect 4649 8299 4707 8305
rect 4738 8296 4744 8308
rect 4796 8336 4802 8348
rect 5750 8336 5756 8348
rect 4796 8308 5756 8336
rect 4796 8296 4802 8308
rect 5750 8296 5756 8308
rect 5808 8296 5814 8348
rect 8418 8296 8424 8348
rect 8476 8336 8482 8348
rect 8970 8336 8976 8348
rect 8476 8308 8976 8336
rect 8476 8296 8482 8308
rect 8970 8296 8976 8308
rect 9028 8296 9034 8348
rect 11454 8336 11460 8348
rect 11415 8308 11460 8336
rect 11454 8296 11460 8308
rect 11512 8296 11518 8348
rect 15229 8339 15287 8345
rect 15229 8305 15241 8339
rect 15275 8305 15287 8339
rect 15229 8299 15287 8305
rect 9062 8228 9068 8280
rect 9120 8268 9126 8280
rect 14674 8268 14680 8280
rect 9120 8240 14680 8268
rect 9120 8228 9126 8240
rect 14674 8228 14680 8240
rect 14732 8228 14738 8280
rect 14766 8228 14772 8280
rect 14824 8268 14830 8280
rect 15244 8268 15272 8299
rect 15318 8296 15324 8348
rect 15376 8336 15382 8348
rect 15413 8339 15471 8345
rect 15413 8336 15425 8339
rect 15376 8308 15425 8336
rect 15376 8296 15382 8308
rect 15413 8305 15425 8308
rect 15459 8305 15471 8339
rect 15594 8336 15600 8348
rect 15507 8308 15600 8336
rect 15413 8299 15471 8305
rect 15594 8296 15600 8308
rect 15652 8336 15658 8348
rect 16422 8336 16428 8348
rect 15652 8308 16428 8336
rect 15652 8296 15658 8308
rect 16422 8296 16428 8308
rect 16480 8296 16486 8348
rect 17710 8336 17716 8348
rect 17671 8308 17716 8336
rect 17710 8296 17716 8308
rect 17768 8296 17774 8348
rect 18262 8336 18268 8348
rect 18223 8308 18268 8336
rect 18262 8296 18268 8308
rect 18320 8296 18326 8348
rect 23414 8296 23420 8348
rect 23472 8336 23478 8348
rect 23601 8339 23659 8345
rect 23601 8336 23613 8339
rect 23472 8308 23613 8336
rect 23472 8296 23478 8308
rect 23601 8305 23613 8308
rect 23647 8305 23659 8339
rect 24242 8336 24248 8348
rect 24203 8308 24248 8336
rect 23601 8299 23659 8305
rect 24242 8296 24248 8308
rect 24300 8296 24306 8348
rect 26085 8339 26143 8345
rect 26085 8305 26097 8339
rect 26131 8336 26143 8339
rect 26174 8336 26180 8348
rect 26131 8308 26180 8336
rect 26131 8305 26143 8308
rect 26085 8299 26143 8305
rect 26174 8296 26180 8308
rect 26232 8296 26238 8348
rect 15686 8268 15692 8280
rect 14824 8240 14869 8268
rect 15244 8240 15692 8268
rect 14824 8228 14830 8240
rect 15686 8228 15692 8240
rect 15744 8228 15750 8280
rect 23506 8268 23512 8280
rect 23467 8240 23512 8268
rect 23506 8228 23512 8240
rect 23564 8228 23570 8280
rect 23966 8268 23972 8280
rect 23927 8240 23972 8268
rect 23966 8228 23972 8240
rect 24024 8228 24030 8280
rect 24521 8271 24579 8277
rect 24521 8237 24533 8271
rect 24567 8268 24579 8271
rect 24567 8240 26128 8268
rect 24567 8237 24579 8240
rect 24521 8231 24579 8237
rect 12653 8203 12711 8209
rect 12653 8169 12665 8203
rect 12699 8200 12711 8203
rect 13110 8200 13116 8212
rect 12699 8172 13116 8200
rect 12699 8169 12711 8172
rect 12653 8163 12711 8169
rect 13110 8160 13116 8172
rect 13168 8160 13174 8212
rect 23690 8160 23696 8212
rect 23748 8200 23754 8212
rect 24536 8200 24564 8231
rect 23748 8172 24564 8200
rect 23748 8160 23754 8172
rect 1702 8132 1708 8144
rect 1663 8104 1708 8132
rect 1702 8092 1708 8104
rect 1760 8092 1766 8144
rect 6029 8135 6087 8141
rect 6029 8101 6041 8135
rect 6075 8132 6087 8135
rect 6118 8132 6124 8144
rect 6075 8104 6124 8132
rect 6075 8101 6087 8104
rect 6029 8095 6087 8101
rect 6118 8092 6124 8104
rect 6176 8092 6182 8144
rect 12469 8135 12527 8141
rect 12469 8101 12481 8135
rect 12515 8132 12527 8135
rect 12926 8132 12932 8144
rect 12515 8104 12932 8132
rect 12515 8101 12527 8104
rect 12469 8095 12527 8101
rect 12926 8092 12932 8104
rect 12984 8092 12990 8144
rect 17802 8132 17808 8144
rect 17763 8104 17808 8132
rect 17802 8092 17808 8104
rect 17860 8132 17866 8144
rect 18541 8135 18599 8141
rect 18541 8132 18553 8135
rect 17860 8104 18553 8132
rect 17860 8092 17866 8104
rect 18541 8101 18553 8104
rect 18587 8132 18599 8135
rect 18630 8132 18636 8144
rect 18587 8104 18636 8132
rect 18587 8101 18599 8104
rect 18541 8095 18599 8101
rect 18630 8092 18636 8104
rect 18688 8092 18694 8144
rect 18814 8132 18820 8144
rect 18775 8104 18820 8132
rect 18814 8092 18820 8104
rect 18872 8092 18878 8144
rect 26100 8141 26128 8240
rect 26085 8135 26143 8141
rect 26085 8101 26097 8135
rect 26131 8132 26143 8135
rect 26266 8132 26272 8144
rect 26131 8104 26272 8132
rect 26131 8101 26143 8104
rect 26085 8095 26143 8101
rect 26266 8092 26272 8104
rect 26324 8092 26330 8144
rect 400 8042 27264 8064
rect 400 7990 3510 8042
rect 3562 7990 3574 8042
rect 3626 7990 3638 8042
rect 3690 7990 3702 8042
rect 3754 7990 3766 8042
rect 3818 7990 27264 8042
rect 400 7968 27264 7990
rect 1518 7888 1524 7940
rect 1576 7928 1582 7940
rect 1613 7931 1671 7937
rect 1613 7928 1625 7931
rect 1576 7900 1625 7928
rect 1576 7888 1582 7900
rect 1613 7897 1625 7900
rect 1659 7897 1671 7931
rect 1613 7891 1671 7897
rect 1702 7888 1708 7940
rect 1760 7928 1766 7940
rect 1797 7931 1855 7937
rect 1797 7928 1809 7931
rect 1760 7900 1809 7928
rect 1760 7888 1766 7900
rect 1797 7897 1809 7900
rect 1843 7897 1855 7931
rect 4186 7928 4192 7940
rect 4147 7900 4192 7928
rect 1797 7891 1855 7897
rect 4186 7888 4192 7900
rect 4244 7888 4250 7940
rect 4370 7928 4376 7940
rect 4331 7900 4376 7928
rect 4370 7888 4376 7900
rect 4428 7888 4434 7940
rect 4557 7931 4615 7937
rect 4557 7897 4569 7931
rect 4603 7928 4615 7931
rect 5750 7928 5756 7940
rect 4603 7900 5756 7928
rect 4603 7897 4615 7900
rect 4557 7891 4615 7897
rect 5750 7888 5756 7900
rect 5808 7888 5814 7940
rect 6118 7928 6124 7940
rect 6079 7900 6124 7928
rect 6118 7888 6124 7900
rect 6176 7888 6182 7940
rect 9062 7928 9068 7940
rect 9023 7900 9068 7928
rect 9062 7888 9068 7900
rect 9120 7888 9126 7940
rect 11365 7931 11423 7937
rect 11365 7897 11377 7931
rect 11411 7928 11423 7931
rect 11454 7928 11460 7940
rect 11411 7900 11460 7928
rect 11411 7897 11423 7900
rect 11365 7891 11423 7897
rect 11454 7888 11460 7900
rect 11512 7888 11518 7940
rect 11825 7931 11883 7937
rect 11825 7897 11837 7931
rect 11871 7928 11883 7931
rect 12006 7928 12012 7940
rect 11871 7900 12012 7928
rect 11871 7897 11883 7900
rect 11825 7891 11883 7897
rect 12006 7888 12012 7900
rect 12064 7928 12070 7940
rect 12193 7931 12251 7937
rect 12193 7928 12205 7931
rect 12064 7900 12205 7928
rect 12064 7888 12070 7900
rect 12193 7897 12205 7900
rect 12239 7928 12251 7931
rect 13386 7928 13392 7940
rect 12239 7900 13392 7928
rect 12239 7897 12251 7900
rect 12193 7891 12251 7897
rect 13386 7888 13392 7900
rect 13444 7888 13450 7940
rect 15226 7928 15232 7940
rect 15187 7900 15232 7928
rect 15226 7888 15232 7900
rect 15284 7888 15290 7940
rect 16977 7931 17035 7937
rect 16977 7897 16989 7931
rect 17023 7928 17035 7931
rect 17802 7928 17808 7940
rect 17023 7900 17808 7928
rect 17023 7897 17035 7900
rect 16977 7891 17035 7897
rect 17802 7888 17808 7900
rect 17860 7888 17866 7940
rect 20565 7931 20623 7937
rect 20565 7897 20577 7931
rect 20611 7928 20623 7931
rect 20930 7928 20936 7940
rect 20611 7900 20936 7928
rect 20611 7897 20623 7900
rect 20565 7891 20623 7897
rect 20930 7888 20936 7900
rect 20988 7888 20994 7940
rect 21482 7928 21488 7940
rect 21443 7900 21488 7928
rect 21482 7888 21488 7900
rect 21540 7888 21546 7940
rect 23141 7931 23199 7937
rect 23141 7897 23153 7931
rect 23187 7928 23199 7931
rect 23414 7928 23420 7940
rect 23187 7900 23420 7928
rect 23187 7897 23199 7900
rect 23141 7891 23199 7897
rect 23414 7888 23420 7900
rect 23472 7888 23478 7940
rect 23690 7928 23696 7940
rect 23651 7900 23696 7928
rect 23690 7888 23696 7900
rect 23748 7888 23754 7940
rect 23966 7928 23972 7940
rect 23927 7900 23972 7928
rect 23966 7888 23972 7900
rect 24024 7888 24030 7940
rect 26266 7928 26272 7940
rect 26227 7900 26272 7928
rect 26266 7888 26272 7900
rect 26324 7888 26330 7940
rect 8970 7820 8976 7872
rect 9028 7860 9034 7872
rect 9157 7863 9215 7869
rect 9157 7860 9169 7863
rect 9028 7832 9169 7860
rect 9028 7820 9034 7832
rect 9157 7829 9169 7832
rect 9203 7829 9215 7863
rect 9157 7823 9215 7829
rect 12101 7863 12159 7869
rect 12101 7829 12113 7863
rect 12147 7860 12159 7863
rect 14401 7863 14459 7869
rect 14401 7860 14413 7863
rect 12147 7832 14413 7860
rect 12147 7829 12159 7832
rect 12101 7823 12159 7829
rect 14401 7829 14413 7832
rect 14447 7860 14459 7863
rect 15045 7863 15103 7869
rect 15045 7860 15057 7863
rect 14447 7832 15057 7860
rect 14447 7829 14459 7832
rect 14401 7823 14459 7829
rect 15045 7829 15057 7832
rect 15091 7860 15103 7863
rect 15594 7860 15600 7872
rect 15091 7832 15600 7860
rect 15091 7829 15103 7832
rect 15045 7823 15103 7829
rect 15594 7820 15600 7832
rect 15652 7820 15658 7872
rect 23325 7863 23383 7869
rect 23325 7829 23337 7863
rect 23371 7860 23383 7863
rect 23984 7860 24012 7888
rect 23371 7832 24012 7860
rect 23371 7829 23383 7832
rect 23325 7823 23383 7829
rect 1521 7795 1579 7801
rect 1521 7761 1533 7795
rect 1567 7792 1579 7795
rect 1610 7792 1616 7804
rect 1567 7764 1616 7792
rect 1567 7761 1579 7764
rect 1521 7755 1579 7761
rect 1610 7752 1616 7764
rect 1668 7752 1674 7804
rect 12926 7792 12932 7804
rect 12887 7764 12932 7792
rect 12926 7752 12932 7764
rect 12984 7752 12990 7804
rect 13478 7752 13484 7804
rect 13536 7792 13542 7804
rect 17618 7792 17624 7804
rect 13536 7764 17624 7792
rect 13536 7752 13542 7764
rect 17618 7752 17624 7764
rect 17676 7752 17682 7804
rect 18354 7752 18360 7804
rect 18412 7792 18418 7804
rect 18814 7792 18820 7804
rect 18412 7764 18820 7792
rect 18412 7752 18418 7764
rect 18814 7752 18820 7764
rect 18872 7792 18878 7804
rect 19093 7795 19151 7801
rect 19093 7792 19105 7795
rect 18872 7764 19105 7792
rect 18872 7752 18878 7764
rect 19093 7761 19105 7764
rect 19139 7761 19151 7795
rect 19093 7755 19151 7761
rect 20010 7752 20016 7804
rect 20068 7792 20074 7804
rect 20657 7795 20715 7801
rect 20657 7792 20669 7795
rect 20068 7764 20669 7792
rect 20068 7752 20074 7764
rect 20657 7761 20669 7764
rect 20703 7792 20715 7795
rect 21301 7795 21359 7801
rect 21301 7792 21313 7795
rect 20703 7764 21313 7792
rect 20703 7761 20715 7764
rect 20657 7755 20715 7761
rect 21301 7761 21313 7764
rect 21347 7761 21359 7795
rect 23984 7792 24012 7832
rect 24429 7795 24487 7801
rect 24429 7792 24441 7795
rect 23984 7764 24441 7792
rect 21301 7755 21359 7761
rect 24429 7761 24441 7764
rect 24475 7761 24487 7795
rect 24429 7755 24487 7761
rect 12377 7659 12435 7665
rect 12377 7625 12389 7659
rect 12423 7656 12435 7659
rect 12558 7656 12564 7668
rect 12423 7628 12564 7656
rect 12423 7625 12435 7628
rect 12377 7619 12435 7625
rect 12558 7616 12564 7628
rect 12616 7616 12622 7668
rect 12944 7656 12972 7752
rect 13018 7684 13024 7736
rect 13076 7724 13082 7736
rect 13386 7724 13392 7736
rect 13076 7696 13121 7724
rect 13347 7696 13392 7724
rect 13076 7684 13082 7696
rect 13386 7684 13392 7696
rect 13444 7684 13450 7736
rect 13573 7727 13631 7733
rect 13573 7693 13585 7727
rect 13619 7724 13631 7727
rect 14401 7727 14459 7733
rect 14401 7724 14413 7727
rect 13619 7696 14413 7724
rect 13619 7693 13631 7696
rect 13573 7687 13631 7693
rect 14401 7693 14413 7696
rect 14447 7693 14459 7727
rect 14401 7687 14459 7693
rect 15689 7727 15747 7733
rect 15689 7693 15701 7727
rect 15735 7724 15747 7727
rect 15870 7724 15876 7736
rect 15735 7696 15876 7724
rect 15735 7693 15747 7696
rect 15689 7687 15747 7693
rect 15870 7684 15876 7696
rect 15928 7684 15934 7736
rect 17161 7727 17219 7733
rect 17161 7693 17173 7727
rect 17207 7724 17219 7727
rect 18446 7724 18452 7736
rect 17207 7696 18452 7724
rect 17207 7693 17219 7696
rect 17161 7687 17219 7693
rect 18446 7684 18452 7696
rect 18504 7684 18510 7736
rect 18630 7724 18636 7736
rect 18591 7696 18636 7724
rect 18630 7684 18636 7696
rect 18688 7684 18694 7736
rect 18909 7727 18967 7733
rect 18909 7693 18921 7727
rect 18955 7693 18967 7727
rect 19458 7724 19464 7736
rect 19419 7696 19464 7724
rect 18909 7687 18967 7693
rect 14585 7659 14643 7665
rect 14585 7656 14597 7659
rect 12944 7628 14597 7656
rect 14585 7625 14597 7628
rect 14631 7656 14643 7659
rect 14766 7656 14772 7668
rect 14631 7628 14772 7656
rect 14631 7625 14643 7628
rect 14585 7619 14643 7625
rect 14766 7616 14772 7628
rect 14824 7616 14830 7668
rect 15778 7656 15784 7668
rect 15691 7628 15784 7656
rect 15778 7616 15784 7628
rect 15836 7656 15842 7668
rect 16057 7659 16115 7665
rect 16057 7656 16069 7659
rect 15836 7628 16069 7656
rect 15836 7616 15842 7628
rect 16057 7625 16069 7628
rect 16103 7625 16115 7659
rect 17894 7656 17900 7668
rect 17807 7628 17900 7656
rect 16057 7619 16115 7625
rect 17894 7616 17900 7628
rect 17952 7656 17958 7668
rect 17989 7659 18047 7665
rect 17989 7656 18001 7659
rect 17952 7628 18001 7656
rect 17952 7616 17958 7628
rect 17989 7625 18001 7628
rect 18035 7625 18047 7659
rect 17989 7619 18047 7625
rect 18078 7616 18084 7668
rect 18136 7656 18142 7668
rect 18924 7656 18952 7687
rect 19458 7684 19464 7696
rect 19516 7684 19522 7736
rect 20749 7727 20807 7733
rect 20749 7724 20761 7727
rect 19706 7696 20761 7724
rect 19706 7656 19734 7696
rect 20749 7693 20761 7696
rect 20795 7724 20807 7727
rect 21482 7724 21488 7736
rect 20795 7696 21488 7724
rect 20795 7693 20807 7696
rect 20749 7687 20807 7693
rect 21482 7684 21488 7696
rect 21540 7684 21546 7736
rect 23874 7684 23880 7736
rect 23932 7724 23938 7736
rect 24153 7727 24211 7733
rect 24153 7724 24165 7727
rect 23932 7696 24165 7724
rect 23932 7684 23938 7696
rect 24153 7693 24165 7696
rect 24199 7693 24211 7727
rect 24153 7687 24211 7693
rect 18136 7628 19734 7656
rect 18136 7616 18142 7628
rect 24886 7616 24892 7668
rect 24944 7616 24950 7668
rect 26174 7656 26180 7668
rect 26135 7628 26180 7656
rect 26174 7616 26180 7628
rect 26232 7656 26238 7668
rect 26453 7659 26511 7665
rect 26453 7656 26465 7659
rect 26232 7628 26465 7656
rect 26232 7616 26238 7628
rect 26453 7625 26465 7628
rect 26499 7625 26511 7659
rect 26453 7619 26511 7625
rect 11362 7548 11368 7600
rect 11420 7588 11426 7600
rect 11457 7591 11515 7597
rect 11457 7588 11469 7591
rect 11420 7560 11469 7588
rect 11420 7548 11426 7560
rect 11457 7557 11469 7560
rect 11503 7557 11515 7591
rect 14858 7588 14864 7600
rect 14771 7560 14864 7588
rect 11457 7551 11515 7557
rect 14858 7548 14864 7560
rect 14916 7588 14922 7600
rect 15686 7588 15692 7600
rect 14916 7560 15692 7588
rect 14916 7548 14922 7560
rect 15686 7548 15692 7560
rect 15744 7548 15750 7600
rect 17526 7588 17532 7600
rect 17487 7560 17532 7588
rect 17526 7548 17532 7560
rect 17584 7548 17590 7600
rect 17618 7548 17624 7600
rect 17676 7588 17682 7600
rect 17713 7591 17771 7597
rect 17713 7588 17725 7591
rect 17676 7560 17725 7588
rect 17676 7548 17682 7560
rect 17713 7557 17725 7560
rect 17759 7588 17771 7591
rect 19458 7588 19464 7600
rect 17759 7560 19464 7588
rect 17759 7557 17771 7560
rect 17713 7551 17771 7557
rect 19458 7548 19464 7560
rect 19516 7548 19522 7600
rect 23506 7588 23512 7600
rect 23467 7560 23512 7588
rect 23506 7548 23512 7560
rect 23564 7548 23570 7600
rect 23877 7591 23935 7597
rect 23877 7557 23889 7591
rect 23923 7588 23935 7591
rect 24242 7588 24248 7600
rect 23923 7560 24248 7588
rect 23923 7557 23935 7560
rect 23877 7551 23935 7557
rect 24242 7548 24248 7560
rect 24300 7548 24306 7600
rect 400 7498 27264 7520
rect 400 7446 18870 7498
rect 18922 7446 18934 7498
rect 18986 7446 18998 7498
rect 19050 7446 19062 7498
rect 19114 7446 19126 7498
rect 19178 7446 27264 7498
rect 400 7424 27264 7446
rect 9890 7384 9896 7396
rect 9632 7356 9896 7384
rect 6578 7316 6584 7328
rect 6504 7288 6584 7316
rect 874 7208 880 7260
rect 932 7248 938 7260
rect 1334 7248 1340 7260
rect 932 7220 1340 7248
rect 932 7208 938 7220
rect 1334 7208 1340 7220
rect 1392 7248 1398 7260
rect 1613 7251 1671 7257
rect 1613 7248 1625 7251
rect 1392 7220 1625 7248
rect 1392 7208 1398 7220
rect 1613 7217 1625 7220
rect 1659 7217 1671 7251
rect 1613 7211 1671 7217
rect 5842 7208 5848 7260
rect 5900 7248 5906 7260
rect 6504 7257 6532 7288
rect 6578 7276 6584 7288
rect 6636 7276 6642 7328
rect 8418 7316 8424 7328
rect 6688 7288 8424 7316
rect 6688 7260 6716 7288
rect 8418 7276 8424 7288
rect 8476 7276 8482 7328
rect 9632 7260 9660 7356
rect 9890 7344 9896 7356
rect 9948 7344 9954 7396
rect 12469 7387 12527 7393
rect 12469 7353 12481 7387
rect 12515 7384 12527 7387
rect 13018 7384 13024 7396
rect 12515 7356 13024 7384
rect 12515 7353 12527 7356
rect 12469 7347 12527 7353
rect 13018 7344 13024 7356
rect 13076 7344 13082 7396
rect 15594 7344 15600 7396
rect 15652 7344 15658 7396
rect 17710 7384 17716 7396
rect 17671 7356 17716 7384
rect 17710 7344 17716 7356
rect 17768 7344 17774 7396
rect 18078 7384 18084 7396
rect 18039 7356 18084 7384
rect 18078 7344 18084 7356
rect 18136 7344 18142 7396
rect 19458 7344 19464 7396
rect 19516 7384 19522 7396
rect 20933 7387 20991 7393
rect 20933 7384 20945 7387
rect 19516 7356 20945 7384
rect 19516 7344 19522 7356
rect 20933 7353 20945 7356
rect 20979 7384 20991 7387
rect 21298 7384 21304 7396
rect 20979 7356 21304 7384
rect 20979 7353 20991 7356
rect 20933 7347 20991 7353
rect 21298 7344 21304 7356
rect 21356 7344 21362 7396
rect 23874 7344 23880 7396
rect 23932 7384 23938 7396
rect 24337 7387 24395 7393
rect 24337 7384 24349 7387
rect 23932 7356 24349 7384
rect 23932 7344 23938 7356
rect 24337 7353 24349 7356
rect 24383 7353 24395 7387
rect 24337 7347 24395 7353
rect 24613 7387 24671 7393
rect 24613 7353 24625 7387
rect 24659 7384 24671 7387
rect 26174 7384 26180 7396
rect 24659 7356 26180 7384
rect 24659 7353 24671 7356
rect 24613 7347 24671 7353
rect 26174 7344 26180 7356
rect 26232 7344 26238 7396
rect 12558 7316 12564 7328
rect 12519 7288 12564 7316
rect 12558 7276 12564 7288
rect 12616 7276 12622 7328
rect 15612 7316 15640 7344
rect 15612 7288 16008 7316
rect 6305 7251 6363 7257
rect 6305 7248 6317 7251
rect 5900 7220 6317 7248
rect 5900 7208 5906 7220
rect 6305 7217 6317 7220
rect 6351 7217 6363 7251
rect 6305 7211 6363 7217
rect 6489 7251 6547 7257
rect 6489 7217 6501 7251
rect 6535 7217 6547 7251
rect 6670 7248 6676 7260
rect 6583 7220 6676 7248
rect 6489 7211 6547 7217
rect 6670 7208 6676 7220
rect 6728 7208 6734 7260
rect 8878 7208 8884 7260
rect 8936 7248 8942 7260
rect 9433 7251 9491 7257
rect 9433 7248 9445 7251
rect 8936 7220 9445 7248
rect 8936 7208 8942 7220
rect 9433 7217 9445 7220
rect 9479 7217 9491 7251
rect 9614 7248 9620 7260
rect 9527 7220 9620 7248
rect 9433 7211 9491 7217
rect 9614 7208 9620 7220
rect 9672 7208 9678 7260
rect 9890 7248 9896 7260
rect 9851 7220 9896 7248
rect 9890 7208 9896 7220
rect 9948 7208 9954 7260
rect 11178 7208 11184 7260
rect 11236 7248 11242 7260
rect 11273 7251 11331 7257
rect 11273 7248 11285 7251
rect 11236 7220 11285 7248
rect 11236 7208 11242 7220
rect 11273 7217 11285 7220
rect 11319 7217 11331 7251
rect 12834 7248 12840 7260
rect 12795 7220 12840 7248
rect 11273 7211 11331 7217
rect 12834 7208 12840 7220
rect 12892 7208 12898 7260
rect 14214 7208 14220 7260
rect 14272 7248 14278 7260
rect 15980 7257 16008 7288
rect 17434 7276 17440 7328
rect 17492 7316 17498 7328
rect 24245 7319 24303 7325
rect 17492 7288 18860 7316
rect 17492 7276 17498 7288
rect 15597 7251 15655 7257
rect 15597 7248 15609 7251
rect 14272 7220 15609 7248
rect 14272 7208 14278 7220
rect 15597 7217 15609 7220
rect 15643 7217 15655 7251
rect 15597 7211 15655 7217
rect 15965 7251 16023 7257
rect 15965 7217 15977 7251
rect 16011 7217 16023 7251
rect 16146 7248 16152 7260
rect 16107 7220 16152 7248
rect 15965 7211 16023 7217
rect 16146 7208 16152 7220
rect 16204 7208 16210 7260
rect 17618 7248 17624 7260
rect 17452 7220 17624 7248
rect 966 7140 972 7192
rect 1024 7180 1030 7192
rect 2165 7183 2223 7189
rect 2165 7180 2177 7183
rect 1024 7152 2177 7180
rect 1024 7140 1030 7152
rect 2165 7149 2177 7152
rect 2211 7180 2223 7183
rect 3358 7180 3364 7192
rect 2211 7152 3364 7180
rect 2211 7149 2223 7152
rect 2165 7143 2223 7149
rect 3358 7140 3364 7152
rect 3416 7140 3422 7192
rect 8973 7183 9031 7189
rect 8973 7149 8985 7183
rect 9019 7180 9031 7183
rect 9522 7180 9528 7192
rect 9019 7152 9528 7180
rect 9019 7149 9031 7152
rect 8973 7143 9031 7149
rect 9522 7140 9528 7152
rect 9580 7140 9586 7192
rect 10074 7180 10080 7192
rect 10035 7152 10080 7180
rect 10074 7140 10080 7152
rect 10132 7140 10138 7192
rect 10353 7183 10411 7189
rect 10353 7149 10365 7183
rect 10399 7149 10411 7183
rect 12742 7180 12748 7192
rect 12703 7152 12748 7180
rect 10353 7143 10411 7149
rect 1521 7115 1579 7121
rect 1521 7081 1533 7115
rect 1567 7112 1579 7115
rect 2070 7112 2076 7124
rect 1567 7084 2076 7112
rect 1567 7081 1579 7084
rect 1521 7075 1579 7081
rect 2070 7072 2076 7084
rect 2128 7072 2134 7124
rect 6121 7115 6179 7121
rect 6121 7081 6133 7115
rect 6167 7112 6179 7115
rect 6578 7112 6584 7124
rect 6167 7084 6584 7112
rect 6167 7081 6179 7084
rect 6121 7075 6179 7081
rect 6578 7072 6584 7084
rect 6636 7072 6642 7124
rect 9246 7072 9252 7124
rect 9304 7112 9310 7124
rect 10368 7112 10396 7143
rect 12742 7140 12748 7152
rect 12800 7140 12806 7192
rect 15686 7180 15692 7192
rect 15599 7152 15692 7180
rect 15686 7140 15692 7152
rect 15744 7180 15750 7192
rect 17452 7180 17480 7220
rect 17618 7208 17624 7220
rect 17676 7208 17682 7260
rect 18832 7257 18860 7288
rect 24245 7285 24257 7319
rect 24291 7316 24303 7319
rect 24886 7316 24892 7328
rect 24291 7288 24892 7316
rect 24291 7285 24303 7288
rect 24245 7279 24303 7285
rect 24886 7276 24892 7288
rect 24944 7276 24950 7328
rect 18817 7251 18875 7257
rect 18817 7217 18829 7251
rect 18863 7248 18875 7251
rect 19093 7251 19151 7257
rect 18863 7220 18952 7248
rect 18863 7217 18875 7220
rect 18817 7211 18875 7217
rect 15744 7152 17480 7180
rect 15744 7140 15750 7152
rect 17526 7140 17532 7192
rect 17584 7180 17590 7192
rect 18262 7180 18268 7192
rect 17584 7152 18268 7180
rect 17584 7140 17590 7152
rect 18262 7140 18268 7152
rect 18320 7180 18326 7192
rect 18630 7180 18636 7192
rect 18320 7152 18636 7180
rect 18320 7140 18326 7152
rect 18630 7140 18636 7152
rect 18688 7140 18694 7192
rect 18170 7112 18176 7124
rect 9304 7084 18176 7112
rect 9304 7072 9310 7084
rect 18170 7072 18176 7084
rect 18228 7072 18234 7124
rect 18924 7112 18952 7220
rect 19093 7217 19105 7251
rect 19139 7248 19151 7251
rect 19642 7248 19648 7260
rect 19139 7220 19648 7248
rect 19139 7217 19151 7220
rect 19093 7211 19151 7217
rect 19642 7208 19648 7220
rect 19700 7208 19706 7260
rect 20010 7208 20016 7260
rect 20068 7248 20074 7260
rect 20289 7251 20347 7257
rect 20289 7248 20301 7251
rect 20068 7220 20301 7248
rect 20068 7208 20074 7220
rect 20289 7217 20301 7220
rect 20335 7217 20347 7251
rect 21577 7251 21635 7257
rect 21577 7248 21589 7251
rect 20289 7211 20347 7217
rect 20488 7220 21589 7248
rect 19274 7180 19280 7192
rect 19235 7152 19280 7180
rect 19274 7140 19280 7152
rect 19332 7140 19338 7192
rect 20102 7140 20108 7192
rect 20160 7180 20166 7192
rect 20197 7183 20255 7189
rect 20197 7180 20209 7183
rect 20160 7152 20209 7180
rect 20160 7140 20166 7152
rect 20197 7149 20209 7152
rect 20243 7149 20255 7183
rect 20197 7143 20255 7149
rect 20378 7112 20384 7124
rect 18924 7084 20384 7112
rect 20378 7072 20384 7084
rect 20436 7072 20442 7124
rect 11362 7044 11368 7056
rect 11323 7016 11368 7044
rect 11362 7004 11368 7016
rect 11420 7004 11426 7056
rect 13021 7047 13079 7053
rect 13021 7013 13033 7047
rect 13067 7044 13079 7047
rect 13110 7044 13116 7056
rect 13067 7016 13116 7044
rect 13067 7013 13079 7016
rect 13021 7007 13079 7013
rect 13110 7004 13116 7016
rect 13168 7004 13174 7056
rect 15042 7044 15048 7056
rect 15003 7016 15048 7044
rect 15042 7004 15048 7016
rect 15100 7004 15106 7056
rect 19642 7004 19648 7056
rect 19700 7044 19706 7056
rect 20488 7053 20516 7220
rect 21577 7217 21589 7220
rect 21623 7248 21635 7251
rect 22034 7248 22040 7260
rect 21623 7220 22040 7248
rect 21623 7217 21635 7220
rect 21577 7211 21635 7217
rect 22034 7208 22040 7220
rect 22092 7208 22098 7260
rect 20473 7047 20531 7053
rect 20473 7044 20485 7047
rect 19700 7016 20485 7044
rect 19700 7004 19706 7016
rect 20473 7013 20485 7016
rect 20519 7013 20531 7047
rect 20473 7007 20531 7013
rect 21117 7047 21175 7053
rect 21117 7013 21129 7047
rect 21163 7044 21175 7047
rect 21666 7044 21672 7056
rect 21163 7016 21672 7044
rect 21163 7013 21175 7016
rect 21117 7007 21175 7013
rect 21666 7004 21672 7016
rect 21724 7004 21730 7056
rect 400 6954 27264 6976
rect 400 6902 3510 6954
rect 3562 6902 3574 6954
rect 3626 6902 3638 6954
rect 3690 6902 3702 6954
rect 3754 6902 3766 6954
rect 3818 6902 27264 6954
rect 400 6880 27264 6902
rect 966 6840 972 6852
rect 927 6812 972 6840
rect 966 6800 972 6812
rect 1024 6800 1030 6852
rect 1334 6840 1340 6852
rect 1295 6812 1340 6840
rect 1334 6800 1340 6812
rect 1392 6840 1398 6852
rect 2441 6843 2499 6849
rect 2441 6840 2453 6843
rect 1392 6812 2453 6840
rect 1392 6800 1398 6812
rect 2441 6809 2453 6812
rect 2487 6809 2499 6843
rect 2441 6803 2499 6809
rect 5842 6800 5848 6852
rect 5900 6840 5906 6852
rect 6121 6843 6179 6849
rect 6121 6840 6133 6843
rect 5900 6812 6133 6840
rect 5900 6800 5906 6812
rect 6121 6809 6133 6812
rect 6167 6809 6179 6843
rect 6121 6803 6179 6809
rect 6581 6843 6639 6849
rect 6581 6809 6593 6843
rect 6627 6840 6639 6843
rect 6670 6840 6676 6852
rect 6627 6812 6676 6840
rect 6627 6809 6639 6812
rect 6581 6803 6639 6809
rect 6670 6800 6676 6812
rect 6728 6800 6734 6852
rect 8602 6840 8608 6852
rect 8563 6812 8608 6840
rect 8602 6800 8608 6812
rect 8660 6800 8666 6852
rect 8878 6840 8884 6852
rect 8839 6812 8884 6840
rect 8878 6800 8884 6812
rect 8936 6800 8942 6852
rect 9246 6840 9252 6852
rect 9207 6812 9252 6840
rect 9246 6800 9252 6812
rect 9304 6800 9310 6852
rect 9522 6840 9528 6852
rect 9483 6812 9528 6840
rect 9522 6800 9528 6812
rect 9580 6800 9586 6852
rect 10350 6800 10356 6852
rect 10408 6840 10414 6852
rect 10445 6843 10503 6849
rect 10445 6840 10457 6843
rect 10408 6812 10457 6840
rect 10408 6800 10414 6812
rect 10445 6809 10457 6812
rect 10491 6840 10503 6843
rect 12558 6840 12564 6852
rect 10491 6812 12564 6840
rect 10491 6809 10503 6812
rect 10445 6803 10503 6809
rect 12558 6800 12564 6812
rect 12616 6800 12622 6852
rect 13110 6840 13116 6852
rect 13071 6812 13116 6840
rect 13110 6800 13116 6812
rect 13168 6800 13174 6852
rect 14490 6800 14496 6852
rect 14548 6840 14554 6852
rect 14585 6843 14643 6849
rect 14585 6840 14597 6843
rect 14548 6812 14597 6840
rect 14548 6800 14554 6812
rect 14585 6809 14597 6812
rect 14631 6840 14643 6843
rect 16146 6840 16152 6852
rect 14631 6812 16152 6840
rect 14631 6809 14643 6812
rect 14585 6803 14643 6809
rect 16146 6800 16152 6812
rect 16204 6800 16210 6852
rect 19093 6843 19151 6849
rect 19093 6809 19105 6843
rect 19139 6840 19151 6843
rect 19274 6840 19280 6852
rect 19139 6812 19280 6840
rect 19139 6809 19151 6812
rect 19093 6803 19151 6809
rect 5937 6775 5995 6781
rect 5937 6741 5949 6775
rect 5983 6772 5995 6775
rect 6486 6772 6492 6784
rect 5983 6744 6492 6772
rect 5983 6741 5995 6744
rect 5937 6735 5995 6741
rect 6486 6732 6492 6744
rect 6544 6732 6550 6784
rect 9433 6775 9491 6781
rect 9433 6741 9445 6775
rect 9479 6772 9491 6775
rect 9614 6772 9620 6784
rect 9479 6744 9620 6772
rect 9479 6741 9491 6744
rect 9433 6735 9491 6741
rect 9614 6732 9620 6744
rect 9672 6732 9678 6784
rect 11178 6732 11184 6784
rect 11236 6772 11242 6784
rect 11457 6775 11515 6781
rect 11457 6772 11469 6775
rect 11236 6744 11469 6772
rect 11236 6732 11242 6744
rect 11457 6741 11469 6744
rect 11503 6741 11515 6775
rect 11457 6735 11515 6741
rect 14769 6775 14827 6781
rect 14769 6741 14781 6775
rect 14815 6772 14827 6775
rect 15594 6772 15600 6784
rect 14815 6744 15600 6772
rect 14815 6741 14827 6744
rect 14769 6735 14827 6741
rect 15594 6732 15600 6744
rect 15652 6732 15658 6784
rect 15686 6732 15692 6784
rect 15744 6772 15750 6784
rect 17986 6772 17992 6784
rect 15744 6744 17992 6772
rect 15744 6732 15750 6744
rect 9065 6707 9123 6713
rect 9065 6673 9077 6707
rect 9111 6704 9123 6707
rect 10074 6704 10080 6716
rect 9111 6676 10080 6704
rect 9111 6673 9123 6676
rect 9065 6667 9123 6673
rect 10074 6664 10080 6676
rect 10132 6664 10138 6716
rect 14401 6707 14459 6713
rect 14401 6673 14413 6707
rect 14447 6704 14459 6707
rect 15505 6707 15563 6713
rect 15505 6704 15517 6707
rect 14447 6676 15517 6704
rect 14447 6673 14459 6676
rect 14401 6667 14459 6673
rect 15505 6673 15517 6676
rect 15551 6704 15563 6707
rect 16054 6704 16060 6716
rect 15551 6676 16060 6704
rect 15551 6673 15563 6676
rect 15505 6667 15563 6673
rect 16054 6664 16060 6676
rect 16112 6664 16118 6716
rect 16164 6713 16192 6744
rect 17986 6732 17992 6744
rect 18044 6732 18050 6784
rect 16149 6707 16207 6713
rect 16149 6673 16161 6707
rect 16195 6673 16207 6707
rect 19108 6704 19136 6803
rect 19274 6800 19280 6812
rect 19332 6800 19338 6852
rect 19921 6843 19979 6849
rect 19921 6809 19933 6843
rect 19967 6840 19979 6843
rect 20010 6840 20016 6852
rect 19967 6812 20016 6840
rect 19967 6809 19979 6812
rect 19921 6803 19979 6809
rect 20010 6800 20016 6812
rect 20068 6800 20074 6852
rect 22034 6840 22040 6852
rect 21995 6812 22040 6840
rect 22034 6800 22040 6812
rect 22092 6800 22098 6852
rect 20473 6775 20531 6781
rect 20473 6741 20485 6775
rect 20519 6772 20531 6775
rect 20933 6775 20991 6781
rect 20933 6772 20945 6775
rect 20519 6744 20945 6772
rect 20519 6741 20531 6744
rect 20473 6735 20531 6741
rect 20933 6741 20945 6744
rect 20979 6772 20991 6775
rect 21206 6772 21212 6784
rect 20979 6744 21212 6772
rect 20979 6741 20991 6744
rect 20933 6735 20991 6741
rect 21206 6732 21212 6744
rect 21264 6732 21270 6784
rect 16149 6667 16207 6673
rect 18004 6676 19136 6704
rect 1334 6596 1340 6648
rect 1392 6636 1398 6648
rect 1429 6639 1487 6645
rect 1429 6636 1441 6639
rect 1392 6608 1441 6636
rect 1392 6596 1398 6608
rect 1429 6605 1441 6608
rect 1475 6605 1487 6639
rect 2070 6636 2076 6648
rect 2031 6608 2076 6636
rect 1429 6599 1487 6605
rect 2070 6596 2076 6608
rect 2128 6636 2134 6648
rect 3177 6639 3235 6645
rect 3177 6636 3189 6639
rect 2128 6608 3189 6636
rect 2128 6596 2134 6608
rect 3177 6605 3189 6608
rect 3223 6636 3235 6639
rect 3453 6639 3511 6645
rect 3453 6636 3465 6639
rect 3223 6608 3465 6636
rect 3223 6605 3235 6608
rect 3177 6599 3235 6605
rect 3453 6605 3465 6608
rect 3499 6605 3511 6639
rect 3453 6599 3511 6605
rect 6026 6596 6032 6648
rect 6084 6636 6090 6648
rect 7041 6639 7099 6645
rect 7041 6636 7053 6639
rect 6084 6608 7053 6636
rect 6084 6596 6090 6608
rect 7041 6605 7053 6608
rect 7087 6636 7099 6639
rect 7314 6636 7320 6648
rect 7087 6608 7320 6636
rect 7087 6605 7099 6608
rect 7041 6599 7099 6605
rect 7314 6596 7320 6608
rect 7372 6596 7378 6648
rect 8602 6596 8608 6648
rect 8660 6636 8666 6648
rect 9890 6636 9896 6648
rect 8660 6608 9896 6636
rect 8660 6596 8666 6608
rect 9890 6596 9896 6608
rect 9948 6636 9954 6648
rect 10718 6636 10724 6648
rect 9948 6608 10724 6636
rect 9948 6596 9954 6608
rect 10718 6596 10724 6608
rect 10776 6596 10782 6648
rect 12834 6596 12840 6648
rect 12892 6636 12898 6648
rect 13021 6639 13079 6645
rect 13021 6636 13033 6639
rect 12892 6608 13033 6636
rect 12892 6596 12898 6608
rect 13021 6605 13033 6608
rect 13067 6636 13079 6639
rect 15045 6639 15103 6645
rect 15045 6636 15057 6639
rect 13067 6608 15057 6636
rect 13067 6605 13079 6608
rect 13021 6599 13079 6605
rect 15045 6605 15057 6608
rect 15091 6605 15103 6639
rect 15045 6599 15103 6605
rect 1153 6571 1211 6577
rect 1153 6537 1165 6571
rect 1199 6568 1211 6571
rect 2346 6568 2352 6580
rect 1199 6540 2352 6568
rect 1199 6537 1211 6540
rect 1153 6531 1211 6537
rect 2346 6528 2352 6540
rect 2404 6528 2410 6580
rect 2990 6528 2996 6580
rect 3048 6568 3054 6580
rect 3361 6571 3419 6577
rect 3361 6568 3373 6571
rect 3048 6540 3373 6568
rect 3048 6528 3054 6540
rect 3361 6537 3373 6540
rect 3407 6568 3419 6571
rect 3637 6571 3695 6577
rect 3637 6568 3649 6571
rect 3407 6540 3649 6568
rect 3407 6537 3419 6540
rect 3361 6531 3419 6537
rect 3637 6537 3649 6540
rect 3683 6537 3695 6571
rect 3637 6531 3695 6537
rect 6397 6571 6455 6577
rect 6397 6537 6409 6571
rect 6443 6568 6455 6571
rect 6578 6568 6584 6580
rect 6443 6540 6584 6568
rect 6443 6537 6455 6540
rect 6397 6531 6455 6537
rect 6578 6528 6584 6540
rect 6636 6528 6642 6580
rect 9709 6571 9767 6577
rect 9709 6537 9721 6571
rect 9755 6537 9767 6571
rect 9709 6531 9767 6537
rect 6857 6503 6915 6509
rect 6857 6469 6869 6503
rect 6903 6500 6915 6503
rect 7133 6503 7191 6509
rect 7133 6500 7145 6503
rect 6903 6472 7145 6500
rect 6903 6469 6915 6472
rect 6857 6463 6915 6469
rect 7133 6469 7145 6472
rect 7179 6500 7191 6503
rect 7222 6500 7228 6512
rect 7179 6472 7228 6500
rect 7179 6469 7191 6472
rect 7133 6463 7191 6469
rect 7222 6460 7228 6472
rect 7280 6460 7286 6512
rect 9724 6500 9752 6531
rect 9798 6528 9804 6580
rect 9856 6568 9862 6580
rect 10261 6571 10319 6577
rect 10261 6568 10273 6571
rect 9856 6540 10273 6568
rect 9856 6528 9862 6540
rect 10261 6537 10273 6540
rect 10307 6568 10319 6571
rect 10537 6571 10595 6577
rect 10537 6568 10549 6571
rect 10307 6540 10549 6568
rect 10307 6537 10319 6540
rect 10261 6531 10319 6537
rect 10537 6537 10549 6540
rect 10583 6537 10595 6571
rect 14858 6568 14864 6580
rect 14819 6540 14864 6568
rect 10537 6531 10595 6537
rect 14858 6528 14864 6540
rect 14916 6528 14922 6580
rect 15060 6568 15088 6599
rect 15134 6596 15140 6648
rect 15192 6636 15198 6648
rect 15321 6639 15379 6645
rect 15192 6608 15237 6636
rect 15192 6596 15198 6608
rect 15321 6605 15333 6639
rect 15367 6636 15379 6639
rect 15686 6636 15692 6648
rect 15367 6608 15692 6636
rect 15367 6605 15379 6608
rect 15321 6599 15379 6605
rect 15686 6596 15692 6608
rect 15744 6596 15750 6648
rect 18004 6645 18032 6676
rect 21298 6664 21304 6716
rect 21356 6704 21362 6716
rect 21485 6707 21543 6713
rect 21485 6704 21497 6707
rect 21356 6676 21497 6704
rect 21356 6664 21362 6676
rect 21485 6673 21497 6676
rect 21531 6673 21543 6707
rect 21485 6667 21543 6673
rect 23506 6664 23512 6716
rect 23564 6704 23570 6716
rect 23564 6676 23874 6704
rect 23564 6664 23570 6676
rect 17713 6639 17771 6645
rect 17713 6605 17725 6639
rect 17759 6636 17771 6639
rect 17989 6639 18047 6645
rect 17989 6636 18001 6639
rect 17759 6608 18001 6636
rect 17759 6605 17771 6608
rect 17713 6599 17771 6605
rect 17989 6605 18001 6608
rect 18035 6605 18047 6639
rect 17989 6599 18047 6605
rect 18081 6639 18139 6645
rect 18081 6605 18093 6639
rect 18127 6605 18139 6639
rect 18081 6599 18139 6605
rect 18265 6639 18323 6645
rect 18265 6605 18277 6639
rect 18311 6636 18323 6639
rect 18538 6636 18544 6648
rect 18311 6608 18544 6636
rect 18311 6605 18323 6608
rect 18265 6599 18323 6605
rect 15226 6568 15232 6580
rect 15060 6540 15232 6568
rect 15226 6528 15232 6540
rect 15284 6568 15290 6580
rect 15778 6568 15784 6580
rect 15284 6540 15784 6568
rect 15284 6528 15290 6540
rect 15778 6528 15784 6540
rect 15836 6528 15842 6580
rect 16146 6528 16152 6580
rect 16204 6568 16210 6580
rect 17161 6571 17219 6577
rect 17161 6568 17173 6571
rect 16204 6540 17173 6568
rect 16204 6528 16210 6540
rect 17161 6537 17173 6540
rect 17207 6568 17219 6571
rect 17897 6571 17955 6577
rect 17207 6540 17664 6568
rect 17207 6537 17219 6540
rect 17161 6531 17219 6537
rect 10350 6500 10356 6512
rect 9724 6472 10356 6500
rect 10350 6460 10356 6472
rect 10408 6460 10414 6512
rect 11362 6500 11368 6512
rect 11323 6472 11368 6500
rect 11362 6460 11368 6472
rect 11420 6500 11426 6512
rect 12742 6500 12748 6512
rect 11420 6472 12748 6500
rect 11420 6460 11426 6472
rect 12742 6460 12748 6472
rect 12800 6460 12806 6512
rect 14214 6460 14220 6512
rect 14272 6500 14278 6512
rect 14272 6472 14317 6500
rect 14272 6460 14278 6472
rect 15134 6460 15140 6512
rect 15192 6500 15198 6512
rect 15873 6503 15931 6509
rect 15873 6500 15885 6503
rect 15192 6472 15885 6500
rect 15192 6460 15198 6472
rect 15873 6469 15885 6472
rect 15919 6500 15931 6503
rect 17434 6500 17440 6512
rect 15919 6472 17440 6500
rect 15919 6469 15931 6472
rect 15873 6463 15931 6469
rect 17434 6460 17440 6472
rect 17492 6460 17498 6512
rect 17636 6500 17664 6540
rect 17897 6537 17909 6571
rect 17943 6568 17955 6571
rect 18096 6568 18124 6599
rect 18538 6596 18544 6608
rect 18596 6636 18602 6648
rect 18817 6639 18875 6645
rect 18817 6636 18829 6639
rect 18596 6608 18829 6636
rect 18596 6596 18602 6608
rect 18817 6605 18829 6608
rect 18863 6605 18875 6639
rect 20930 6636 20936 6648
rect 20891 6608 20936 6636
rect 18817 6599 18875 6605
rect 20930 6596 20936 6608
rect 20988 6596 20994 6648
rect 21209 6639 21267 6645
rect 21209 6605 21221 6639
rect 21255 6605 21267 6639
rect 21666 6636 21672 6648
rect 21627 6608 21672 6636
rect 21209 6599 21267 6605
rect 20102 6568 20108 6580
rect 17943 6540 20108 6568
rect 17943 6537 17955 6540
rect 17897 6531 17955 6537
rect 20102 6528 20108 6540
rect 20160 6568 20166 6580
rect 20289 6571 20347 6577
rect 20289 6568 20301 6571
rect 20160 6540 20301 6568
rect 20160 6528 20166 6540
rect 20289 6537 20301 6540
rect 20335 6568 20347 6571
rect 21224 6568 21252 6599
rect 21666 6596 21672 6608
rect 21724 6636 21730 6648
rect 22221 6639 22279 6645
rect 22221 6636 22233 6639
rect 21724 6608 22233 6636
rect 21724 6596 21730 6608
rect 22221 6605 22233 6608
rect 22267 6605 22279 6639
rect 22221 6599 22279 6605
rect 22310 6568 22316 6580
rect 20335 6540 22316 6568
rect 20335 6537 20347 6540
rect 20289 6531 20347 6537
rect 22310 6528 22316 6540
rect 22368 6528 22374 6580
rect 23846 6568 23874 6676
rect 24886 6664 24892 6716
rect 24944 6704 24950 6716
rect 25349 6707 25407 6713
rect 25349 6704 25361 6707
rect 24944 6676 25361 6704
rect 24944 6664 24950 6676
rect 25349 6673 25361 6676
rect 25395 6704 25407 6707
rect 25901 6707 25959 6713
rect 25901 6704 25913 6707
rect 25395 6676 25913 6704
rect 25395 6673 25407 6676
rect 25349 6667 25407 6673
rect 25901 6673 25913 6676
rect 25947 6673 25959 6707
rect 25901 6667 25959 6673
rect 24245 6639 24303 6645
rect 24245 6605 24257 6639
rect 24291 6636 24303 6639
rect 24291 6608 24656 6636
rect 24291 6605 24303 6608
rect 24245 6599 24303 6605
rect 24337 6571 24395 6577
rect 24337 6568 24349 6571
rect 23846 6540 24349 6568
rect 24337 6537 24349 6540
rect 24383 6568 24395 6571
rect 24429 6571 24487 6577
rect 24429 6568 24441 6571
rect 24383 6540 24441 6568
rect 24383 6537 24395 6540
rect 24337 6531 24395 6537
rect 24429 6537 24441 6540
rect 24475 6537 24487 6571
rect 24429 6531 24487 6537
rect 24628 6512 24656 6608
rect 25070 6596 25076 6648
rect 25128 6636 25134 6648
rect 25165 6639 25223 6645
rect 25165 6636 25177 6639
rect 25128 6608 25177 6636
rect 25128 6596 25134 6608
rect 25165 6605 25177 6608
rect 25211 6636 25223 6639
rect 25717 6639 25775 6645
rect 25717 6636 25729 6639
rect 25211 6608 25729 6636
rect 25211 6605 25223 6608
rect 25165 6599 25223 6605
rect 25717 6605 25729 6608
rect 25763 6605 25775 6639
rect 25717 6599 25775 6605
rect 18449 6503 18507 6509
rect 18449 6500 18461 6503
rect 17636 6472 18461 6500
rect 18449 6469 18461 6472
rect 18495 6469 18507 6503
rect 19642 6500 19648 6512
rect 19603 6472 19648 6500
rect 18449 6463 18507 6469
rect 19642 6460 19648 6472
rect 19700 6460 19706 6512
rect 24610 6500 24616 6512
rect 24571 6472 24616 6500
rect 24610 6460 24616 6472
rect 24668 6460 24674 6512
rect 400 6410 27264 6432
rect 400 6358 18870 6410
rect 18922 6358 18934 6410
rect 18986 6358 18998 6410
rect 19050 6358 19062 6410
rect 19114 6358 19126 6410
rect 19178 6358 27264 6410
rect 400 6336 27264 6358
rect 1150 6296 1156 6308
rect 800 6268 1156 6296
rect 800 6169 828 6268
rect 1150 6256 1156 6268
rect 1208 6296 1214 6308
rect 1702 6296 1708 6308
rect 1208 6268 1708 6296
rect 1208 6256 1214 6268
rect 1702 6256 1708 6268
rect 1760 6256 1766 6308
rect 1981 6299 2039 6305
rect 1981 6265 1993 6299
rect 2027 6296 2039 6299
rect 2070 6296 2076 6308
rect 2027 6268 2076 6296
rect 2027 6265 2039 6268
rect 1981 6259 2039 6265
rect 2070 6256 2076 6268
rect 2128 6256 2134 6308
rect 3358 6296 3364 6308
rect 3319 6268 3364 6296
rect 3358 6256 3364 6268
rect 3416 6256 3422 6308
rect 10350 6296 10356 6308
rect 10311 6268 10356 6296
rect 10350 6256 10356 6268
rect 10408 6256 10414 6308
rect 11178 6256 11184 6308
rect 11236 6296 11242 6308
rect 11917 6299 11975 6305
rect 11917 6296 11929 6299
rect 11236 6268 11929 6296
rect 11236 6256 11242 6268
rect 11917 6265 11929 6268
rect 11963 6296 11975 6299
rect 12834 6296 12840 6308
rect 11963 6268 12840 6296
rect 11963 6265 11975 6268
rect 11917 6259 11975 6265
rect 12834 6256 12840 6268
rect 12892 6256 12898 6308
rect 15042 6256 15048 6308
rect 15100 6296 15106 6308
rect 15413 6299 15471 6305
rect 15413 6296 15425 6299
rect 15100 6268 15425 6296
rect 15100 6256 15106 6268
rect 15413 6265 15425 6268
rect 15459 6265 15471 6299
rect 15413 6259 15471 6265
rect 18541 6299 18599 6305
rect 18541 6265 18553 6299
rect 18587 6296 18599 6299
rect 19642 6296 19648 6308
rect 18587 6268 19648 6296
rect 18587 6265 18599 6268
rect 18541 6259 18599 6265
rect 19642 6256 19648 6268
rect 19700 6256 19706 6308
rect 20930 6296 20936 6308
rect 20891 6268 20936 6296
rect 20930 6256 20936 6268
rect 20988 6256 20994 6308
rect 874 6188 880 6240
rect 932 6228 938 6240
rect 932 6200 1748 6228
rect 932 6188 938 6200
rect 1720 6169 1748 6200
rect 6578 6188 6584 6240
rect 6636 6228 6642 6240
rect 12282 6228 12288 6240
rect 6636 6200 12288 6228
rect 6636 6188 6642 6200
rect 12282 6188 12288 6200
rect 12340 6188 12346 6240
rect 14214 6188 14220 6240
rect 14272 6228 14278 6240
rect 14582 6228 14588 6240
rect 14272 6200 14588 6228
rect 14272 6188 14278 6200
rect 14582 6188 14588 6200
rect 14640 6188 14646 6240
rect 15226 6228 15232 6240
rect 15187 6200 15232 6228
rect 15226 6188 15232 6200
rect 15284 6188 15290 6240
rect 18630 6228 18636 6240
rect 18591 6200 18636 6228
rect 18630 6188 18636 6200
rect 18688 6188 18694 6240
rect 20197 6231 20255 6237
rect 20197 6228 20209 6231
rect 19706 6200 20209 6228
rect 785 6163 843 6169
rect 785 6129 797 6163
rect 831 6129 843 6163
rect 785 6123 843 6129
rect 1613 6163 1671 6169
rect 1613 6129 1625 6163
rect 1659 6129 1671 6163
rect 1613 6123 1671 6129
rect 1705 6163 1763 6169
rect 1705 6129 1717 6163
rect 1751 6129 1763 6163
rect 1705 6123 1763 6129
rect 877 6095 935 6101
rect 877 6061 889 6095
rect 923 6092 935 6095
rect 1242 6092 1248 6104
rect 923 6064 1248 6092
rect 923 6061 935 6064
rect 877 6055 935 6061
rect 1242 6052 1248 6064
rect 1300 6052 1306 6104
rect 1628 6092 1656 6123
rect 2346 6120 2352 6172
rect 2404 6160 2410 6172
rect 3266 6160 3272 6172
rect 2404 6132 3272 6160
rect 2404 6120 2410 6132
rect 3266 6120 3272 6132
rect 3324 6160 3330 6172
rect 3545 6163 3603 6169
rect 3545 6160 3557 6163
rect 3324 6132 3557 6160
rect 3324 6120 3330 6132
rect 3545 6129 3557 6132
rect 3591 6160 3603 6163
rect 5293 6163 5351 6169
rect 5293 6160 5305 6163
rect 3591 6132 5305 6160
rect 3591 6129 3603 6132
rect 3545 6123 3603 6129
rect 5293 6129 5305 6132
rect 5339 6160 5351 6163
rect 5658 6160 5664 6172
rect 5339 6132 5664 6160
rect 5339 6129 5351 6132
rect 5293 6123 5351 6129
rect 5658 6120 5664 6132
rect 5716 6120 5722 6172
rect 6394 6160 6400 6172
rect 6355 6132 6400 6160
rect 6394 6120 6400 6132
rect 6452 6120 6458 6172
rect 7130 6160 7136 6172
rect 7091 6132 7136 6160
rect 7130 6120 7136 6132
rect 7188 6120 7194 6172
rect 7314 6160 7320 6172
rect 7275 6132 7320 6160
rect 7314 6120 7320 6132
rect 7372 6120 7378 6172
rect 8970 6120 8976 6172
rect 9028 6160 9034 6172
rect 9525 6163 9583 6169
rect 9525 6160 9537 6163
rect 9028 6132 9537 6160
rect 9028 6120 9034 6132
rect 9525 6129 9537 6132
rect 9571 6129 9583 6163
rect 9525 6123 9583 6129
rect 10269 6163 10327 6169
rect 10269 6129 10281 6163
rect 10315 6160 10327 6163
rect 10718 6160 10724 6172
rect 10315 6132 10724 6160
rect 10315 6129 10327 6132
rect 10269 6123 10327 6129
rect 10718 6120 10724 6132
rect 10776 6120 10782 6172
rect 14766 6160 14772 6172
rect 14727 6132 14772 6160
rect 14766 6120 14772 6132
rect 14824 6120 14830 6172
rect 16054 6160 16060 6172
rect 16015 6132 16060 6160
rect 16054 6120 16060 6132
rect 16112 6120 16118 6172
rect 17618 6160 17624 6172
rect 17579 6132 17624 6160
rect 17618 6120 17624 6132
rect 17676 6160 17682 6172
rect 19706 6160 19734 6200
rect 20197 6197 20209 6200
rect 20243 6228 20255 6231
rect 20286 6228 20292 6240
rect 20243 6200 20292 6228
rect 20243 6197 20255 6200
rect 20197 6191 20255 6197
rect 20286 6188 20292 6200
rect 20344 6228 20350 6240
rect 21666 6228 21672 6240
rect 20344 6200 21672 6228
rect 20344 6188 20350 6200
rect 21666 6188 21672 6200
rect 21724 6188 21730 6240
rect 20378 6160 20384 6172
rect 17676 6132 19734 6160
rect 20339 6132 20384 6160
rect 17676 6120 17682 6132
rect 20378 6120 20384 6132
rect 20436 6120 20442 6172
rect 22129 6163 22187 6169
rect 22129 6129 22141 6163
rect 22175 6160 22187 6163
rect 22494 6160 22500 6172
rect 22175 6132 22500 6160
rect 22175 6129 22187 6132
rect 22129 6123 22187 6129
rect 22494 6120 22500 6132
rect 22552 6120 22558 6172
rect 24242 6160 24248 6172
rect 24203 6132 24248 6160
rect 24242 6120 24248 6132
rect 24300 6120 24306 6172
rect 24429 6163 24487 6169
rect 24429 6129 24441 6163
rect 24475 6160 24487 6163
rect 24610 6160 24616 6172
rect 24475 6132 24616 6160
rect 24475 6129 24487 6132
rect 24429 6123 24487 6129
rect 1794 6092 1800 6104
rect 1628 6064 1800 6092
rect 1794 6052 1800 6064
rect 1852 6052 1858 6104
rect 4830 6092 4836 6104
rect 4791 6064 4836 6092
rect 4830 6052 4836 6064
rect 4888 6052 4894 6104
rect 5382 6092 5388 6104
rect 5343 6064 5388 6092
rect 5382 6052 5388 6064
rect 5440 6052 5446 6104
rect 9433 6095 9491 6101
rect 9433 6061 9445 6095
rect 9479 6092 9491 6095
rect 9798 6092 9804 6104
rect 9479 6064 9804 6092
rect 9479 6061 9491 6064
rect 9433 6055 9491 6061
rect 9798 6052 9804 6064
rect 9856 6052 9862 6104
rect 15137 6095 15195 6101
rect 15137 6092 15149 6095
rect 14186 6064 15149 6092
rect 11825 6027 11883 6033
rect 11825 5993 11837 6027
rect 11871 6024 11883 6027
rect 12374 6024 12380 6036
rect 11871 5996 12380 6024
rect 11871 5993 11883 5996
rect 11825 5987 11883 5993
rect 12374 5984 12380 5996
rect 12432 6024 12438 6036
rect 14186 6024 14214 6064
rect 15137 6061 15149 6064
rect 15183 6092 15195 6095
rect 15226 6092 15232 6104
rect 15183 6064 15232 6092
rect 15183 6061 15195 6064
rect 15137 6055 15195 6061
rect 15226 6052 15232 6064
rect 15284 6052 15290 6104
rect 15962 6092 15968 6104
rect 15875 6064 15968 6092
rect 15962 6052 15968 6064
rect 16020 6092 16026 6104
rect 16514 6092 16520 6104
rect 16020 6064 16520 6092
rect 16020 6052 16026 6064
rect 16514 6052 16520 6064
rect 16572 6052 16578 6104
rect 17802 6101 17808 6104
rect 17768 6095 17808 6101
rect 17768 6061 17780 6095
rect 17768 6055 17808 6061
rect 17802 6052 17808 6055
rect 17860 6052 17866 6104
rect 17986 6092 17992 6104
rect 17947 6064 17992 6092
rect 17986 6052 17992 6064
rect 18044 6052 18050 6104
rect 18170 6052 18176 6104
rect 18228 6092 18234 6104
rect 22586 6092 22592 6104
rect 18228 6064 22592 6092
rect 18228 6052 18234 6064
rect 22586 6052 22592 6064
rect 22644 6052 22650 6104
rect 23414 6052 23420 6104
rect 23472 6092 23478 6104
rect 24153 6095 24211 6101
rect 24153 6092 24165 6095
rect 23472 6064 24165 6092
rect 23472 6052 23478 6064
rect 24153 6061 24165 6064
rect 24199 6092 24211 6095
rect 24444 6092 24472 6123
rect 24610 6120 24616 6132
rect 24668 6160 24674 6172
rect 25898 6160 25904 6172
rect 24668 6132 25904 6160
rect 24668 6120 24674 6132
rect 25898 6120 25904 6132
rect 25956 6120 25962 6172
rect 24199 6064 24472 6092
rect 24199 6061 24211 6064
rect 24153 6055 24211 6061
rect 12432 5996 14214 6024
rect 12432 5984 12438 5996
rect 17434 5984 17440 6036
rect 17492 6024 17498 6036
rect 18081 6027 18139 6033
rect 18081 6024 18093 6027
rect 17492 5996 18093 6024
rect 17492 5984 17498 5996
rect 18081 5993 18093 5996
rect 18127 5993 18139 6027
rect 18081 5987 18139 5993
rect 23969 6027 24027 6033
rect 23969 5993 23981 6027
rect 24015 6024 24027 6027
rect 24610 6024 24616 6036
rect 24015 5996 24616 6024
rect 24015 5993 24027 5996
rect 23969 5987 24027 5993
rect 24610 5984 24616 5996
rect 24668 5984 24674 6036
rect 4186 5956 4192 5968
rect 4147 5928 4192 5956
rect 4186 5916 4192 5928
rect 4244 5916 4250 5968
rect 8694 5956 8700 5968
rect 8655 5928 8700 5956
rect 8694 5916 8700 5928
rect 8752 5916 8758 5968
rect 16238 5956 16244 5968
rect 16199 5928 16244 5956
rect 16238 5916 16244 5928
rect 16296 5916 16302 5968
rect 17897 5959 17955 5965
rect 17897 5925 17909 5959
rect 17943 5956 17955 5959
rect 18170 5956 18176 5968
rect 17943 5928 18176 5956
rect 17943 5925 17955 5928
rect 17897 5919 17955 5925
rect 18170 5916 18176 5928
rect 18228 5916 18234 5968
rect 20470 5956 20476 5968
rect 20431 5928 20476 5956
rect 20470 5916 20476 5928
rect 20528 5916 20534 5968
rect 22129 5959 22187 5965
rect 22129 5925 22141 5959
rect 22175 5956 22187 5959
rect 22310 5956 22316 5968
rect 22175 5928 22316 5956
rect 22175 5925 22187 5928
rect 22129 5919 22187 5925
rect 22310 5916 22316 5928
rect 22368 5916 22374 5968
rect 23782 5916 23788 5968
rect 23840 5956 23846 5968
rect 24150 5956 24156 5968
rect 23840 5928 24156 5956
rect 23840 5916 23846 5928
rect 24150 5916 24156 5928
rect 24208 5956 24214 5968
rect 24521 5959 24579 5965
rect 24521 5956 24533 5959
rect 24208 5928 24533 5956
rect 24208 5916 24214 5928
rect 24521 5925 24533 5928
rect 24567 5925 24579 5959
rect 24521 5919 24579 5925
rect 400 5866 27264 5888
rect 400 5814 3510 5866
rect 3562 5814 3574 5866
rect 3626 5814 3638 5866
rect 3690 5814 3702 5866
rect 3754 5814 3766 5866
rect 3818 5814 27264 5866
rect 400 5792 27264 5814
rect 874 5752 880 5764
rect 835 5724 880 5752
rect 874 5712 880 5724
rect 932 5712 938 5764
rect 1150 5752 1156 5764
rect 1111 5724 1156 5752
rect 1150 5712 1156 5724
rect 1208 5712 1214 5764
rect 3266 5712 3272 5764
rect 3324 5752 3330 5764
rect 3453 5755 3511 5761
rect 3453 5752 3465 5755
rect 3324 5724 3465 5752
rect 3324 5712 3330 5724
rect 3453 5721 3465 5724
rect 3499 5721 3511 5755
rect 3453 5715 3511 5721
rect 4830 5712 4836 5764
rect 4888 5752 4894 5764
rect 5293 5755 5351 5761
rect 5293 5752 5305 5755
rect 4888 5724 5305 5752
rect 4888 5712 4894 5724
rect 5293 5721 5305 5724
rect 5339 5721 5351 5755
rect 5293 5715 5351 5721
rect 5382 5712 5388 5764
rect 5440 5752 5446 5764
rect 5477 5755 5535 5761
rect 5477 5752 5489 5755
rect 5440 5724 5489 5752
rect 5440 5712 5446 5724
rect 5477 5721 5489 5724
rect 5523 5721 5535 5755
rect 5658 5752 5664 5764
rect 5619 5724 5664 5752
rect 5477 5715 5535 5721
rect 5658 5712 5664 5724
rect 5716 5712 5722 5764
rect 5937 5755 5995 5761
rect 5937 5721 5949 5755
rect 5983 5752 5995 5755
rect 6026 5752 6032 5764
rect 5983 5724 6032 5752
rect 5983 5721 5995 5724
rect 5937 5715 5995 5721
rect 6026 5712 6032 5724
rect 6084 5712 6090 5764
rect 6394 5752 6400 5764
rect 6307 5724 6400 5752
rect 6394 5712 6400 5724
rect 6452 5752 6458 5764
rect 6581 5755 6639 5761
rect 6581 5752 6593 5755
rect 6452 5724 6593 5752
rect 6452 5712 6458 5724
rect 6581 5721 6593 5724
rect 6627 5752 6639 5755
rect 7409 5755 7467 5761
rect 7409 5752 7421 5755
rect 6627 5724 7421 5752
rect 6627 5721 6639 5724
rect 6581 5715 6639 5721
rect 7409 5721 7421 5724
rect 7455 5752 7467 5755
rect 9522 5752 9528 5764
rect 7455 5724 9528 5752
rect 7455 5721 7467 5724
rect 7409 5715 7467 5721
rect 9522 5712 9528 5724
rect 9580 5712 9586 5764
rect 15962 5752 15968 5764
rect 15923 5724 15968 5752
rect 15962 5712 15968 5724
rect 16020 5712 16026 5764
rect 16054 5712 16060 5764
rect 16112 5752 16118 5764
rect 16149 5755 16207 5761
rect 16149 5752 16161 5755
rect 16112 5724 16161 5752
rect 16112 5712 16118 5724
rect 16149 5721 16161 5724
rect 16195 5721 16207 5755
rect 16149 5715 16207 5721
rect 16238 5712 16244 5764
rect 16296 5752 16302 5764
rect 16333 5755 16391 5761
rect 16333 5752 16345 5755
rect 16296 5724 16345 5752
rect 16296 5712 16302 5724
rect 16333 5721 16345 5724
rect 16379 5721 16391 5755
rect 17618 5752 17624 5764
rect 17579 5724 17624 5752
rect 16333 5715 16391 5721
rect 17618 5712 17624 5724
rect 17676 5712 17682 5764
rect 17894 5752 17900 5764
rect 17855 5724 17900 5752
rect 17894 5712 17900 5724
rect 17952 5712 17958 5764
rect 20286 5752 20292 5764
rect 20247 5724 20292 5752
rect 20286 5712 20292 5724
rect 20344 5712 20350 5764
rect 20470 5752 20476 5764
rect 20431 5724 20476 5752
rect 20470 5712 20476 5724
rect 20528 5712 20534 5764
rect 22310 5752 22316 5764
rect 22271 5724 22316 5752
rect 22310 5712 22316 5724
rect 22368 5712 22374 5764
rect 23414 5752 23420 5764
rect 23375 5724 23420 5752
rect 23414 5712 23420 5724
rect 23472 5712 23478 5764
rect 23601 5755 23659 5761
rect 23601 5721 23613 5755
rect 23647 5752 23659 5755
rect 24242 5752 24248 5764
rect 23647 5724 24248 5752
rect 23647 5721 23659 5724
rect 23601 5715 23659 5721
rect 24242 5712 24248 5724
rect 24300 5712 24306 5764
rect 785 5687 843 5693
rect 785 5653 797 5687
rect 831 5684 843 5687
rect 1794 5684 1800 5696
rect 831 5656 1800 5684
rect 831 5653 843 5656
rect 785 5647 843 5653
rect 1794 5644 1800 5656
rect 1852 5684 1858 5696
rect 2070 5684 2076 5696
rect 1852 5656 2076 5684
rect 1852 5644 1858 5656
rect 2070 5644 2076 5656
rect 2128 5684 2134 5696
rect 3913 5687 3971 5693
rect 3913 5684 3925 5687
rect 2128 5656 3925 5684
rect 2128 5644 2134 5656
rect 3913 5653 3925 5656
rect 3959 5684 3971 5687
rect 4738 5684 4744 5696
rect 3959 5656 4744 5684
rect 3959 5653 3971 5656
rect 3913 5647 3971 5653
rect 4738 5644 4744 5656
rect 4796 5644 4802 5696
rect 2349 5619 2407 5625
rect 2349 5585 2361 5619
rect 2395 5616 2407 5619
rect 2990 5616 2996 5628
rect 2395 5588 2996 5616
rect 2395 5585 2407 5588
rect 2349 5579 2407 5585
rect 2990 5576 2996 5588
rect 3048 5576 3054 5628
rect 3821 5619 3879 5625
rect 3821 5585 3833 5619
rect 3867 5616 3879 5619
rect 3867 5588 4416 5616
rect 3867 5585 3879 5588
rect 3821 5579 3879 5585
rect 1058 5508 1064 5560
rect 1116 5548 1122 5560
rect 2441 5551 2499 5557
rect 2441 5548 2453 5551
rect 1116 5520 2453 5548
rect 1116 5508 1122 5520
rect 2441 5517 2453 5520
rect 2487 5517 2499 5551
rect 2441 5511 2499 5517
rect 2901 5551 2959 5557
rect 2901 5517 2913 5551
rect 2947 5548 2959 5551
rect 4186 5548 4192 5560
rect 2947 5520 3404 5548
rect 4147 5520 4192 5548
rect 2947 5517 2959 5520
rect 2901 5511 2959 5517
rect 2456 5480 2484 5511
rect 3085 5483 3143 5489
rect 3085 5480 3097 5483
rect 2456 5452 3097 5480
rect 3085 5449 3097 5452
rect 3131 5480 3143 5483
rect 3266 5480 3272 5492
rect 3131 5452 3272 5480
rect 3131 5449 3143 5452
rect 3085 5443 3143 5449
rect 3266 5440 3272 5452
rect 3324 5440 3330 5492
rect 3376 5489 3404 5520
rect 4186 5508 4192 5520
rect 4244 5508 4250 5560
rect 3361 5483 3419 5489
rect 3361 5449 3373 5483
rect 3407 5480 3419 5483
rect 4002 5480 4008 5492
rect 3407 5452 4008 5480
rect 3407 5449 3419 5452
rect 3361 5443 3419 5449
rect 4002 5440 4008 5452
rect 4060 5440 4066 5492
rect 4281 5483 4339 5489
rect 4281 5449 4293 5483
rect 4327 5449 4339 5483
rect 4388 5480 4416 5588
rect 4462 5576 4468 5628
rect 4520 5616 4526 5628
rect 4848 5616 4876 5712
rect 6305 5687 6363 5693
rect 6305 5653 6317 5687
rect 6351 5684 6363 5687
rect 6486 5684 6492 5696
rect 6351 5656 6492 5684
rect 6351 5653 6363 5656
rect 6305 5647 6363 5653
rect 6486 5644 6492 5656
rect 6544 5684 6550 5696
rect 7130 5684 7136 5696
rect 6544 5656 7136 5684
rect 6544 5644 6550 5656
rect 7130 5644 7136 5656
rect 7188 5644 7194 5696
rect 14214 5644 14220 5696
rect 14272 5684 14278 5696
rect 14766 5684 14772 5696
rect 14272 5656 14772 5684
rect 14272 5644 14278 5656
rect 14766 5644 14772 5656
rect 14824 5684 14830 5696
rect 15594 5684 15600 5696
rect 14824 5656 15600 5684
rect 14824 5644 14830 5656
rect 15594 5644 15600 5656
rect 15652 5644 15658 5696
rect 6118 5616 6124 5628
rect 4520 5588 4876 5616
rect 5032 5588 6124 5616
rect 4520 5576 4526 5588
rect 4738 5508 4744 5560
rect 4796 5548 4802 5560
rect 5032 5557 5060 5588
rect 6118 5576 6124 5588
rect 6176 5576 6182 5628
rect 6581 5619 6639 5625
rect 6581 5585 6593 5619
rect 6627 5616 6639 5619
rect 6673 5619 6731 5625
rect 6673 5616 6685 5619
rect 6627 5588 6685 5616
rect 6627 5585 6639 5588
rect 6581 5579 6639 5585
rect 6673 5585 6685 5588
rect 6719 5585 6731 5619
rect 7222 5616 7228 5628
rect 7183 5588 7228 5616
rect 6673 5579 6731 5585
rect 7222 5576 7228 5588
rect 7280 5616 7286 5628
rect 7501 5619 7559 5625
rect 7501 5616 7513 5619
rect 7280 5588 7513 5616
rect 7280 5576 7286 5588
rect 7501 5585 7513 5588
rect 7547 5585 7559 5619
rect 7501 5579 7559 5585
rect 8605 5619 8663 5625
rect 8605 5585 8617 5619
rect 8651 5616 8663 5619
rect 8970 5616 8976 5628
rect 8651 5588 8976 5616
rect 8651 5585 8663 5588
rect 8605 5579 8663 5585
rect 8970 5576 8976 5588
rect 9028 5576 9034 5628
rect 10718 5616 10724 5628
rect 10679 5588 10724 5616
rect 10718 5576 10724 5588
rect 10776 5576 10782 5628
rect 11181 5619 11239 5625
rect 11181 5585 11193 5619
rect 11227 5616 11239 5619
rect 13849 5619 13907 5625
rect 11227 5588 12788 5616
rect 11227 5585 11239 5588
rect 11181 5579 11239 5585
rect 12760 5560 12788 5588
rect 13849 5585 13861 5619
rect 13895 5616 13907 5619
rect 16256 5616 16284 5712
rect 13895 5588 16284 5616
rect 17912 5616 17940 5712
rect 23782 5684 23788 5696
rect 23743 5656 23788 5684
rect 23782 5644 23788 5656
rect 23840 5644 23846 5696
rect 18265 5619 18323 5625
rect 18265 5616 18277 5619
rect 17912 5588 18277 5616
rect 13895 5585 13907 5588
rect 13849 5579 13907 5585
rect 5017 5551 5075 5557
rect 5017 5548 5029 5551
rect 4796 5520 5029 5548
rect 4796 5508 4802 5520
rect 5017 5517 5029 5520
rect 5063 5517 5075 5551
rect 5017 5511 5075 5517
rect 5109 5551 5167 5557
rect 5109 5517 5121 5551
rect 5155 5548 5167 5551
rect 6302 5548 6308 5560
rect 5155 5520 6308 5548
rect 5155 5517 5167 5520
rect 5109 5511 5167 5517
rect 5124 5480 5152 5511
rect 6302 5508 6308 5520
rect 6360 5508 6366 5560
rect 8694 5548 8700 5560
rect 8655 5520 8700 5548
rect 8694 5508 8700 5520
rect 8752 5508 8758 5560
rect 11362 5548 11368 5560
rect 11275 5520 11368 5548
rect 11362 5508 11368 5520
rect 11420 5548 11426 5560
rect 12193 5551 12251 5557
rect 12193 5548 12205 5551
rect 11420 5520 12205 5548
rect 11420 5508 11426 5520
rect 12193 5517 12205 5520
rect 12239 5517 12251 5551
rect 12374 5548 12380 5560
rect 12335 5520 12380 5548
rect 12193 5511 12251 5517
rect 12374 5508 12380 5520
rect 12432 5508 12438 5560
rect 12742 5548 12748 5560
rect 12655 5520 12748 5548
rect 12742 5508 12748 5520
rect 12800 5508 12806 5560
rect 12834 5508 12840 5560
rect 12892 5548 12898 5560
rect 14033 5551 14091 5557
rect 12892 5520 12937 5548
rect 12892 5508 12898 5520
rect 14033 5517 14045 5551
rect 14079 5548 14091 5551
rect 14214 5548 14220 5560
rect 14079 5520 14220 5548
rect 14079 5517 14091 5520
rect 14033 5511 14091 5517
rect 14214 5508 14220 5520
rect 14272 5508 14278 5560
rect 14950 5548 14956 5560
rect 14911 5520 14956 5548
rect 14950 5508 14956 5520
rect 15008 5508 15014 5560
rect 15134 5548 15140 5560
rect 15095 5520 15140 5548
rect 15134 5508 15140 5520
rect 15192 5508 15198 5560
rect 15520 5557 15548 5588
rect 18265 5585 18277 5588
rect 18311 5585 18323 5619
rect 18265 5579 18323 5585
rect 18354 5576 18360 5628
rect 18412 5616 18418 5628
rect 20013 5619 20071 5625
rect 20013 5616 20025 5619
rect 18412 5588 20025 5616
rect 18412 5576 18418 5588
rect 20013 5585 20025 5588
rect 20059 5616 20071 5619
rect 20378 5616 20384 5628
rect 20059 5588 20384 5616
rect 20059 5585 20071 5588
rect 20013 5579 20071 5585
rect 20378 5576 20384 5588
rect 20436 5616 20442 5628
rect 20565 5619 20623 5625
rect 20565 5616 20577 5619
rect 20436 5588 20577 5616
rect 20436 5576 20442 5588
rect 20565 5585 20577 5588
rect 20611 5585 20623 5619
rect 23874 5616 23880 5628
rect 23835 5588 23880 5616
rect 20565 5579 20623 5585
rect 23874 5576 23880 5588
rect 23932 5576 23938 5628
rect 24150 5616 24156 5628
rect 24111 5588 24156 5616
rect 24150 5576 24156 5588
rect 24208 5576 24214 5628
rect 25898 5616 25904 5628
rect 25859 5588 25904 5616
rect 25898 5576 25904 5588
rect 25956 5576 25962 5628
rect 15505 5551 15563 5557
rect 15505 5517 15517 5551
rect 15551 5517 15563 5551
rect 15505 5511 15563 5517
rect 15594 5508 15600 5560
rect 15652 5548 15658 5560
rect 15652 5520 15697 5548
rect 15652 5508 15658 5520
rect 15870 5508 15876 5560
rect 15928 5548 15934 5560
rect 17434 5548 17440 5560
rect 15928 5520 17440 5548
rect 15928 5508 15934 5520
rect 17434 5508 17440 5520
rect 17492 5508 17498 5560
rect 17986 5548 17992 5560
rect 17947 5520 17992 5548
rect 17986 5508 17992 5520
rect 18044 5508 18050 5560
rect 19366 5508 19372 5560
rect 19424 5508 19430 5560
rect 19826 5508 19832 5560
rect 19884 5548 19890 5560
rect 21577 5551 21635 5557
rect 21577 5548 21589 5551
rect 19884 5520 21589 5548
rect 19884 5508 19890 5520
rect 21577 5517 21589 5520
rect 21623 5548 21635 5551
rect 21623 5520 22264 5548
rect 21623 5517 21635 5520
rect 21577 5511 21635 5517
rect 4388 5452 5152 5480
rect 8421 5483 8479 5489
rect 4281 5443 4339 5449
rect 8421 5449 8433 5483
rect 8467 5480 8479 5483
rect 8467 5452 8924 5480
rect 8467 5449 8479 5452
rect 8421 5443 8479 5449
rect 1242 5412 1248 5424
rect 1203 5384 1248 5412
rect 1242 5372 1248 5384
rect 1300 5372 1306 5424
rect 4296 5412 4324 5443
rect 4462 5412 4468 5424
rect 4296 5384 4468 5412
rect 4462 5372 4468 5384
rect 4520 5372 4526 5424
rect 8896 5412 8924 5452
rect 8970 5440 8976 5492
rect 9028 5480 9034 5492
rect 9028 5452 9073 5480
rect 9028 5440 9034 5452
rect 9430 5440 9436 5492
rect 9488 5440 9494 5492
rect 11178 5440 11184 5492
rect 11236 5480 11242 5492
rect 11549 5483 11607 5489
rect 11549 5480 11561 5483
rect 11236 5452 11561 5480
rect 11236 5440 11242 5452
rect 11549 5449 11561 5452
rect 11595 5480 11607 5483
rect 11733 5483 11791 5489
rect 11733 5480 11745 5483
rect 11595 5452 11745 5480
rect 11595 5449 11607 5452
rect 11549 5443 11607 5449
rect 11733 5449 11745 5452
rect 11779 5449 11791 5483
rect 11733 5443 11791 5449
rect 14401 5483 14459 5489
rect 14401 5449 14413 5483
rect 14447 5480 14459 5483
rect 14490 5480 14496 5492
rect 14447 5452 14496 5480
rect 14447 5449 14459 5452
rect 14401 5443 14459 5449
rect 14490 5440 14496 5452
rect 14548 5440 14554 5492
rect 14968 5480 14996 5508
rect 15781 5483 15839 5489
rect 15781 5480 15793 5483
rect 14968 5452 15793 5480
rect 15781 5449 15793 5452
rect 15827 5480 15839 5483
rect 17066 5480 17072 5492
rect 15827 5452 17072 5480
rect 15827 5449 15839 5452
rect 15781 5443 15839 5449
rect 17066 5440 17072 5452
rect 17124 5480 17130 5492
rect 17894 5480 17900 5492
rect 17124 5452 17900 5480
rect 17124 5440 17130 5452
rect 17894 5440 17900 5452
rect 17952 5440 17958 5492
rect 22236 5489 22264 5520
rect 21853 5483 21911 5489
rect 21853 5480 21865 5483
rect 21776 5452 21865 5480
rect 9448 5412 9476 5440
rect 21776 5424 21804 5452
rect 21853 5449 21865 5452
rect 21899 5449 21911 5483
rect 21853 5443 21911 5449
rect 22221 5483 22279 5489
rect 22221 5449 22233 5483
rect 22267 5480 22279 5483
rect 22267 5452 23874 5480
rect 22267 5449 22279 5452
rect 22221 5443 22279 5449
rect 13662 5412 13668 5424
rect 8896 5384 9476 5412
rect 13623 5384 13668 5412
rect 13662 5372 13668 5384
rect 13720 5372 13726 5424
rect 21298 5372 21304 5424
rect 21356 5412 21362 5424
rect 21393 5415 21451 5421
rect 21393 5412 21405 5415
rect 21356 5384 21405 5412
rect 21356 5372 21362 5384
rect 21393 5381 21405 5384
rect 21439 5412 21451 5415
rect 21758 5412 21764 5424
rect 21439 5384 21764 5412
rect 21439 5381 21451 5384
rect 21393 5375 21451 5381
rect 21758 5372 21764 5384
rect 21816 5372 21822 5424
rect 22494 5412 22500 5424
rect 22455 5384 22500 5412
rect 22494 5372 22500 5384
rect 22552 5372 22558 5424
rect 23846 5412 23874 5452
rect 24610 5440 24616 5492
rect 24668 5440 24674 5492
rect 24426 5412 24432 5424
rect 23846 5384 24432 5412
rect 24426 5372 24432 5384
rect 24484 5412 24490 5424
rect 25070 5412 25076 5424
rect 24484 5384 25076 5412
rect 24484 5372 24490 5384
rect 25070 5372 25076 5384
rect 25128 5372 25134 5424
rect 400 5322 27264 5344
rect 400 5270 18870 5322
rect 18922 5270 18934 5322
rect 18986 5270 18998 5322
rect 19050 5270 19062 5322
rect 19114 5270 19126 5322
rect 19178 5270 27264 5322
rect 400 5248 27264 5270
rect 3358 5208 3364 5220
rect 3319 5180 3364 5208
rect 3358 5168 3364 5180
rect 3416 5168 3422 5220
rect 4189 5211 4247 5217
rect 4189 5177 4201 5211
rect 4235 5208 4247 5211
rect 4462 5208 4468 5220
rect 4235 5180 4468 5208
rect 4235 5177 4247 5180
rect 4189 5171 4247 5177
rect 4388 5081 4416 5180
rect 4462 5168 4468 5180
rect 4520 5168 4526 5220
rect 6486 5208 6492 5220
rect 6447 5180 6492 5208
rect 6486 5168 6492 5180
rect 6544 5208 6550 5220
rect 6765 5211 6823 5217
rect 6765 5208 6777 5211
rect 6544 5180 6777 5208
rect 6544 5168 6550 5180
rect 6765 5177 6777 5180
rect 6811 5177 6823 5211
rect 6765 5171 6823 5177
rect 8602 5168 8608 5220
rect 8660 5208 8666 5220
rect 8697 5211 8755 5217
rect 8697 5208 8709 5211
rect 8660 5180 8709 5208
rect 8660 5168 8666 5180
rect 8697 5177 8709 5180
rect 8743 5177 8755 5211
rect 8697 5171 8755 5177
rect 8970 5168 8976 5220
rect 9028 5208 9034 5220
rect 9617 5211 9675 5217
rect 9617 5208 9629 5211
rect 9028 5180 9629 5208
rect 9028 5168 9034 5180
rect 9617 5177 9629 5180
rect 9663 5177 9675 5211
rect 9617 5171 9675 5177
rect 9798 5168 9804 5220
rect 9856 5208 9862 5220
rect 9985 5211 10043 5217
rect 9985 5208 9997 5211
rect 9856 5180 9997 5208
rect 9856 5168 9862 5180
rect 9985 5177 9997 5180
rect 10031 5177 10043 5211
rect 9985 5171 10043 5177
rect 10261 5211 10319 5217
rect 10261 5177 10273 5211
rect 10307 5208 10319 5211
rect 10718 5208 10724 5220
rect 10307 5180 10724 5208
rect 10307 5177 10319 5180
rect 10261 5171 10319 5177
rect 10718 5168 10724 5180
rect 10776 5168 10782 5220
rect 13662 5168 13668 5220
rect 13720 5208 13726 5220
rect 13720 5180 14214 5208
rect 13720 5168 13726 5180
rect 5382 5100 5388 5152
rect 5440 5140 5446 5152
rect 6857 5143 6915 5149
rect 6857 5140 6869 5143
rect 5440 5112 6869 5140
rect 5440 5100 5446 5112
rect 6857 5109 6869 5112
rect 6903 5140 6915 5143
rect 6946 5140 6952 5152
rect 6903 5112 6952 5140
rect 6903 5109 6915 5112
rect 6857 5103 6915 5109
rect 6946 5100 6952 5112
rect 7004 5100 7010 5152
rect 9341 5143 9399 5149
rect 9341 5109 9353 5143
rect 9387 5140 9399 5143
rect 9430 5140 9436 5152
rect 9387 5112 9436 5140
rect 9387 5109 9399 5112
rect 9341 5103 9399 5109
rect 9430 5100 9436 5112
rect 9488 5100 9494 5152
rect 9893 5143 9951 5149
rect 9893 5109 9905 5143
rect 9939 5140 9951 5143
rect 10350 5140 10356 5152
rect 9939 5112 10356 5140
rect 9939 5109 9951 5112
rect 9893 5103 9951 5109
rect 10350 5100 10356 5112
rect 10408 5100 10414 5152
rect 11178 5140 11184 5152
rect 11139 5112 11184 5140
rect 11178 5100 11184 5112
rect 11236 5100 11242 5152
rect 11914 5100 11920 5152
rect 11972 5100 11978 5152
rect 12834 5100 12840 5152
rect 12892 5140 12898 5152
rect 12929 5143 12987 5149
rect 12929 5140 12941 5143
rect 12892 5112 12941 5140
rect 12892 5100 12898 5112
rect 12929 5109 12941 5112
rect 12975 5109 12987 5143
rect 14186 5140 14214 5180
rect 14582 5168 14588 5220
rect 14640 5208 14646 5220
rect 15045 5211 15103 5217
rect 15045 5208 15057 5211
rect 14640 5180 15057 5208
rect 14640 5168 14646 5180
rect 15045 5177 15057 5180
rect 15091 5177 15103 5211
rect 15226 5208 15232 5220
rect 15187 5180 15232 5208
rect 15045 5171 15103 5177
rect 15226 5168 15232 5180
rect 15284 5168 15290 5220
rect 17802 5168 17808 5220
rect 17860 5208 17866 5220
rect 17897 5211 17955 5217
rect 17897 5208 17909 5211
rect 17860 5180 17909 5208
rect 17860 5168 17866 5180
rect 17897 5177 17909 5180
rect 17943 5208 17955 5211
rect 18354 5208 18360 5220
rect 17943 5180 18360 5208
rect 17943 5177 17955 5180
rect 17897 5171 17955 5177
rect 18354 5168 18360 5180
rect 18412 5208 18418 5220
rect 23874 5208 23880 5220
rect 18412 5180 18768 5208
rect 23835 5180 23880 5208
rect 18412 5168 18418 5180
rect 14953 5143 15011 5149
rect 14953 5140 14965 5143
rect 14186 5112 14965 5140
rect 12929 5103 12987 5109
rect 14953 5109 14965 5112
rect 14999 5140 15011 5143
rect 15134 5140 15140 5152
rect 14999 5112 15140 5140
rect 14999 5109 15011 5112
rect 14953 5103 15011 5109
rect 15134 5100 15140 5112
rect 15192 5100 15198 5152
rect 17713 5143 17771 5149
rect 17713 5109 17725 5143
rect 17759 5140 17771 5143
rect 18078 5140 18084 5152
rect 17759 5112 18084 5140
rect 17759 5109 17771 5112
rect 17713 5103 17771 5109
rect 18078 5100 18084 5112
rect 18136 5100 18142 5152
rect 4373 5075 4431 5081
rect 4373 5041 4385 5075
rect 4419 5041 4431 5075
rect 4373 5035 4431 5041
rect 5845 5075 5903 5081
rect 5845 5041 5857 5075
rect 5891 5072 5903 5075
rect 6026 5072 6032 5084
rect 5891 5044 6032 5072
rect 5891 5041 5903 5044
rect 5845 5035 5903 5041
rect 6026 5032 6032 5044
rect 6084 5032 6090 5084
rect 9062 5072 9068 5084
rect 9023 5044 9068 5072
rect 9062 5032 9068 5044
rect 9120 5032 9126 5084
rect 14861 5075 14919 5081
rect 14861 5041 14873 5075
rect 14907 5072 14919 5075
rect 15042 5072 15048 5084
rect 14907 5044 15048 5072
rect 14907 5041 14919 5044
rect 14861 5035 14919 5041
rect 15042 5032 15048 5044
rect 15100 5032 15106 5084
rect 15870 5072 15876 5084
rect 15831 5044 15876 5072
rect 15870 5032 15876 5044
rect 15928 5032 15934 5084
rect 18740 5081 18768 5180
rect 23874 5168 23880 5180
rect 23932 5168 23938 5220
rect 24150 5168 24156 5220
rect 24208 5208 24214 5220
rect 24245 5211 24303 5217
rect 24245 5208 24257 5211
rect 24208 5180 24257 5208
rect 24208 5168 24214 5180
rect 24245 5177 24257 5180
rect 24291 5177 24303 5211
rect 24245 5171 24303 5177
rect 18814 5100 18820 5152
rect 18872 5140 18878 5152
rect 19093 5143 19151 5149
rect 19093 5140 19105 5143
rect 18872 5112 19105 5140
rect 18872 5100 18878 5112
rect 19093 5109 19105 5112
rect 19139 5140 19151 5143
rect 19274 5140 19280 5152
rect 19139 5112 19280 5140
rect 19139 5109 19151 5112
rect 19093 5103 19151 5109
rect 19274 5100 19280 5112
rect 19332 5100 19338 5152
rect 21206 5100 21212 5152
rect 21264 5140 21270 5152
rect 21301 5143 21359 5149
rect 21301 5140 21313 5143
rect 21264 5112 21313 5140
rect 21264 5100 21270 5112
rect 21301 5109 21313 5112
rect 21347 5109 21359 5143
rect 21301 5103 21359 5109
rect 21758 5100 21764 5152
rect 21816 5100 21822 5152
rect 24610 5100 24616 5152
rect 24668 5140 24674 5152
rect 24705 5143 24763 5149
rect 24705 5140 24717 5143
rect 24668 5112 24717 5140
rect 24668 5100 24674 5112
rect 24705 5109 24717 5112
rect 24751 5109 24763 5143
rect 24705 5103 24763 5109
rect 18725 5075 18783 5081
rect 18725 5041 18737 5075
rect 18771 5072 18783 5075
rect 18906 5072 18912 5084
rect 18771 5044 18912 5072
rect 18771 5041 18783 5044
rect 18725 5035 18783 5041
rect 18906 5032 18912 5044
rect 18964 5032 18970 5084
rect 24426 5072 24432 5084
rect 24387 5044 24432 5072
rect 24426 5032 24432 5044
rect 24484 5032 24490 5084
rect 10902 5004 10908 5016
rect 10863 4976 10908 5004
rect 10902 4964 10908 4976
rect 10960 4964 10966 5016
rect 15781 5007 15839 5013
rect 15781 4973 15793 5007
rect 15827 5004 15839 5007
rect 15962 5004 15968 5016
rect 15827 4976 15968 5004
rect 15827 4973 15839 4976
rect 15781 4967 15839 4973
rect 15962 4964 15968 4976
rect 16020 4964 16026 5016
rect 17986 4964 17992 5016
rect 18044 5004 18050 5016
rect 18265 5007 18323 5013
rect 18265 5004 18277 5007
rect 18044 4976 18277 5004
rect 18044 4964 18050 4976
rect 18265 4973 18277 4976
rect 18311 5004 18323 5007
rect 21022 5004 21028 5016
rect 18311 4976 21028 5004
rect 18311 4973 18323 4976
rect 18265 4967 18323 4973
rect 21022 4964 21028 4976
rect 21080 4964 21086 5016
rect 22494 4964 22500 5016
rect 22552 5004 22558 5016
rect 23049 5007 23107 5013
rect 23049 5004 23061 5007
rect 22552 4976 23061 5004
rect 22552 4964 22558 4976
rect 23049 4973 23061 4976
rect 23095 4973 23107 5007
rect 23049 4967 23107 4973
rect 5658 4936 5664 4948
rect 5619 4908 5664 4936
rect 5658 4896 5664 4908
rect 5716 4896 5722 4948
rect 18081 4939 18139 4945
rect 18081 4905 18093 4939
rect 18127 4936 18139 4939
rect 18814 4936 18820 4948
rect 18127 4908 18820 4936
rect 18127 4905 18139 4908
rect 18081 4899 18139 4905
rect 18814 4896 18820 4908
rect 18872 4896 18878 4948
rect 2438 4868 2444 4880
rect 2399 4840 2444 4868
rect 2438 4828 2444 4840
rect 2496 4828 2502 4880
rect 14582 4828 14588 4880
rect 14640 4868 14646 4880
rect 16057 4871 16115 4877
rect 16057 4868 16069 4871
rect 14640 4840 16069 4868
rect 14640 4828 14646 4840
rect 16057 4837 16069 4840
rect 16103 4868 16115 4871
rect 16146 4868 16152 4880
rect 16103 4840 16152 4868
rect 16103 4837 16115 4840
rect 16057 4831 16115 4837
rect 16146 4828 16152 4840
rect 16204 4828 16210 4880
rect 400 4778 27264 4800
rect 400 4726 3510 4778
rect 3562 4726 3574 4778
rect 3626 4726 3638 4778
rect 3690 4726 3702 4778
rect 3754 4726 3766 4778
rect 3818 4726 27264 4778
rect 400 4704 27264 4726
rect 2165 4667 2223 4673
rect 2165 4633 2177 4667
rect 2211 4664 2223 4667
rect 2346 4664 2352 4676
rect 2211 4636 2352 4664
rect 2211 4633 2223 4636
rect 2165 4627 2223 4633
rect 2346 4624 2352 4636
rect 2404 4624 2410 4676
rect 4462 4664 4468 4676
rect 4423 4636 4468 4664
rect 4462 4624 4468 4636
rect 4520 4624 4526 4676
rect 4833 4667 4891 4673
rect 4833 4633 4845 4667
rect 4879 4664 4891 4667
rect 6026 4664 6032 4676
rect 4879 4636 6032 4664
rect 4879 4633 4891 4636
rect 4833 4627 4891 4633
rect 6026 4624 6032 4636
rect 6084 4624 6090 4676
rect 6486 4624 6492 4676
rect 6544 4664 6550 4676
rect 6765 4667 6823 4673
rect 6765 4664 6777 4667
rect 6544 4636 6777 4664
rect 6544 4624 6550 4636
rect 6765 4633 6777 4636
rect 6811 4633 6823 4667
rect 6946 4664 6952 4676
rect 6907 4636 6952 4664
rect 6765 4627 6823 4633
rect 6946 4624 6952 4636
rect 7004 4624 7010 4676
rect 9341 4667 9399 4673
rect 9341 4633 9353 4667
rect 9387 4664 9399 4667
rect 9430 4664 9436 4676
rect 9387 4636 9436 4664
rect 9387 4633 9399 4636
rect 9341 4627 9399 4633
rect 9430 4624 9436 4636
rect 9488 4624 9494 4676
rect 10997 4667 11055 4673
rect 10997 4633 11009 4667
rect 11043 4664 11055 4667
rect 11178 4664 11184 4676
rect 11043 4636 11184 4664
rect 11043 4633 11055 4636
rect 10997 4627 11055 4633
rect 11178 4624 11184 4636
rect 11236 4624 11242 4676
rect 12742 4624 12748 4676
rect 12800 4664 12806 4676
rect 13205 4667 13263 4673
rect 13205 4664 13217 4667
rect 12800 4636 13217 4664
rect 12800 4624 12806 4636
rect 13205 4633 13217 4636
rect 13251 4664 13263 4667
rect 13757 4667 13815 4673
rect 13757 4664 13769 4667
rect 13251 4636 13769 4664
rect 13251 4633 13263 4636
rect 13205 4627 13263 4633
rect 13757 4633 13769 4636
rect 13803 4633 13815 4667
rect 13757 4627 13815 4633
rect 14861 4667 14919 4673
rect 14861 4633 14873 4667
rect 14907 4664 14919 4667
rect 15134 4664 15140 4676
rect 14907 4636 15140 4664
rect 14907 4633 14919 4636
rect 14861 4627 14919 4633
rect 15134 4624 15140 4636
rect 15192 4624 15198 4676
rect 15870 4624 15876 4676
rect 15928 4664 15934 4676
rect 15965 4667 16023 4673
rect 15965 4664 15977 4667
rect 15928 4636 15977 4664
rect 15928 4624 15934 4636
rect 15965 4633 15977 4636
rect 16011 4633 16023 4667
rect 16146 4664 16152 4676
rect 16107 4636 16152 4664
rect 15965 4627 16023 4633
rect 16146 4624 16152 4636
rect 16204 4624 16210 4676
rect 18722 4664 18728 4676
rect 18683 4636 18728 4664
rect 18722 4624 18728 4636
rect 18780 4624 18786 4676
rect 18814 4624 18820 4676
rect 18872 4664 18878 4676
rect 19366 4664 19372 4676
rect 18872 4636 19372 4664
rect 18872 4624 18878 4636
rect 19366 4624 19372 4636
rect 19424 4664 19430 4676
rect 19921 4667 19979 4673
rect 19921 4664 19933 4667
rect 19424 4636 19933 4664
rect 19424 4624 19430 4636
rect 19921 4633 19933 4636
rect 19967 4633 19979 4667
rect 21298 4664 21304 4676
rect 21259 4636 21304 4664
rect 19921 4627 19979 4633
rect 21298 4624 21304 4636
rect 21356 4624 21362 4676
rect 21669 4667 21727 4673
rect 21669 4633 21681 4667
rect 21715 4664 21727 4667
rect 22494 4664 22500 4676
rect 21715 4636 22500 4664
rect 21715 4633 21727 4636
rect 21669 4627 21727 4633
rect 22494 4624 22500 4636
rect 22552 4624 22558 4676
rect 24426 4664 24432 4676
rect 24387 4636 24432 4664
rect 24426 4624 24432 4636
rect 24484 4624 24490 4676
rect 24610 4664 24616 4676
rect 24571 4636 24616 4664
rect 24610 4624 24616 4636
rect 24668 4624 24674 4676
rect 2364 4528 2392 4624
rect 11549 4599 11607 4605
rect 11549 4565 11561 4599
rect 11595 4596 11607 4599
rect 12834 4596 12840 4608
rect 11595 4568 12840 4596
rect 11595 4565 11607 4568
rect 11549 4559 11607 4565
rect 12834 4556 12840 4568
rect 12892 4556 12898 4608
rect 14677 4599 14735 4605
rect 14677 4565 14689 4599
rect 14723 4596 14735 4599
rect 15042 4596 15048 4608
rect 14723 4568 15048 4596
rect 14723 4565 14735 4568
rect 14677 4559 14735 4565
rect 15042 4556 15048 4568
rect 15100 4556 15106 4608
rect 18906 4596 18912 4608
rect 18867 4568 18912 4596
rect 18906 4556 18912 4568
rect 18964 4556 18970 4608
rect 19826 4596 19832 4608
rect 19706 4568 19832 4596
rect 4557 4531 4615 4537
rect 4557 4528 4569 4531
rect 2364 4500 4569 4528
rect 2438 4460 2444 4472
rect 2399 4432 2444 4460
rect 2438 4420 2444 4432
rect 2496 4420 2502 4472
rect 3928 4469 3956 4500
rect 4557 4497 4569 4500
rect 4603 4497 4615 4531
rect 4557 4491 4615 4497
rect 6118 4488 6124 4540
rect 6176 4528 6182 4540
rect 10166 4528 10172 4540
rect 6176 4500 10172 4528
rect 6176 4488 6182 4500
rect 10166 4488 10172 4500
rect 10224 4488 10230 4540
rect 11181 4531 11239 4537
rect 11181 4497 11193 4531
rect 11227 4528 11239 4531
rect 11914 4528 11920 4540
rect 11227 4500 11920 4528
rect 11227 4497 11239 4500
rect 11181 4491 11239 4497
rect 11914 4488 11920 4500
rect 11972 4528 11978 4540
rect 12009 4531 12067 4537
rect 12009 4528 12021 4531
rect 11972 4500 12021 4528
rect 11972 4488 11978 4500
rect 12009 4497 12021 4500
rect 12055 4528 12067 4531
rect 12561 4531 12619 4537
rect 12561 4528 12573 4531
rect 12055 4500 12573 4528
rect 12055 4497 12067 4500
rect 12009 4491 12067 4497
rect 12561 4497 12573 4500
rect 12607 4497 12619 4531
rect 12561 4491 12619 4497
rect 15873 4531 15931 4537
rect 15873 4497 15885 4531
rect 15919 4528 15931 4531
rect 15962 4528 15968 4540
rect 15919 4500 15968 4528
rect 15919 4497 15931 4500
rect 15873 4491 15931 4497
rect 15962 4488 15968 4500
rect 16020 4488 16026 4540
rect 18722 4488 18728 4540
rect 18780 4528 18786 4540
rect 19369 4531 19427 4537
rect 19369 4528 19381 4531
rect 18780 4500 19381 4528
rect 18780 4488 18786 4500
rect 19369 4497 19381 4500
rect 19415 4497 19427 4531
rect 19369 4491 19427 4497
rect 3913 4463 3971 4469
rect 3913 4429 3925 4463
rect 3959 4429 3971 4463
rect 3913 4423 3971 4429
rect 11733 4463 11791 4469
rect 11733 4429 11745 4463
rect 11779 4460 11791 4463
rect 11825 4463 11883 4469
rect 11825 4460 11837 4463
rect 11779 4432 11837 4460
rect 11779 4429 11791 4432
rect 11733 4423 11791 4429
rect 11825 4429 11837 4432
rect 11871 4429 11883 4463
rect 11825 4423 11883 4429
rect 12374 4420 12380 4472
rect 12432 4460 12438 4472
rect 13113 4463 13171 4469
rect 13113 4460 13125 4463
rect 12432 4432 13125 4460
rect 12432 4420 12438 4432
rect 13113 4429 13125 4432
rect 13159 4460 13171 4463
rect 13573 4463 13631 4469
rect 13573 4460 13585 4463
rect 13159 4432 13585 4460
rect 13159 4429 13171 4432
rect 13113 4423 13171 4429
rect 13573 4429 13585 4432
rect 13619 4429 13631 4463
rect 13573 4423 13631 4429
rect 17894 4420 17900 4472
rect 17952 4460 17958 4472
rect 19185 4463 19243 4469
rect 19185 4460 19197 4463
rect 17952 4432 19197 4460
rect 17952 4420 17958 4432
rect 19185 4429 19197 4432
rect 19231 4460 19243 4463
rect 19706 4460 19734 4568
rect 19826 4556 19832 4568
rect 19884 4556 19890 4608
rect 21022 4556 21028 4608
rect 21080 4596 21086 4608
rect 21485 4599 21543 4605
rect 21485 4596 21497 4599
rect 21080 4568 21497 4596
rect 21080 4556 21086 4568
rect 21485 4565 21497 4568
rect 21531 4596 21543 4599
rect 23874 4596 23880 4608
rect 21531 4568 23880 4596
rect 21531 4565 21543 4568
rect 21485 4559 21543 4565
rect 23874 4556 23880 4568
rect 23932 4556 23938 4608
rect 21117 4531 21175 4537
rect 21117 4497 21129 4531
rect 21163 4528 21175 4531
rect 21298 4528 21304 4540
rect 21163 4500 21304 4528
rect 21163 4497 21175 4500
rect 21117 4491 21175 4497
rect 21298 4488 21304 4500
rect 21356 4488 21362 4540
rect 19231 4432 19734 4460
rect 19231 4429 19243 4432
rect 19185 4423 19243 4429
rect 2349 4395 2407 4401
rect 2349 4361 2361 4395
rect 2395 4392 2407 4395
rect 4002 4392 4008 4404
rect 2395 4364 4008 4392
rect 2395 4361 2407 4364
rect 2349 4355 2407 4361
rect 4002 4352 4008 4364
rect 4060 4352 4066 4404
rect 8694 4352 8700 4404
rect 8752 4392 8758 4404
rect 10902 4392 10908 4404
rect 8752 4364 10908 4392
rect 8752 4352 8758 4364
rect 10902 4352 10908 4364
rect 10960 4392 10966 4404
rect 11365 4395 11423 4401
rect 11365 4392 11377 4395
rect 10960 4364 11377 4392
rect 10960 4352 10966 4364
rect 11365 4361 11377 4364
rect 11411 4392 11423 4395
rect 11411 4364 12512 4392
rect 11411 4361 11423 4364
rect 11365 4355 11423 4361
rect 6210 4284 6216 4336
rect 6268 4324 6274 4336
rect 9062 4324 9068 4336
rect 6268 4296 9068 4324
rect 6268 4284 6274 4296
rect 9062 4284 9068 4296
rect 9120 4324 9126 4336
rect 11733 4327 11791 4333
rect 11733 4324 11745 4327
rect 9120 4296 11745 4324
rect 9120 4284 9126 4296
rect 11733 4293 11745 4296
rect 11779 4324 11791 4327
rect 12374 4324 12380 4336
rect 11779 4296 12380 4324
rect 11779 4293 11791 4296
rect 11733 4287 11791 4293
rect 12374 4284 12380 4296
rect 12432 4284 12438 4336
rect 12484 4324 12512 4364
rect 15502 4324 15508 4336
rect 12484 4296 15508 4324
rect 15502 4284 15508 4296
rect 15560 4284 15566 4336
rect 400 4234 27264 4256
rect 400 4182 18870 4234
rect 18922 4182 18934 4234
rect 18986 4182 18998 4234
rect 19050 4182 19062 4234
rect 19114 4182 19126 4234
rect 19178 4182 27264 4234
rect 400 4160 27264 4182
rect 23598 4080 23604 4132
rect 23656 4120 23662 4132
rect 23693 4123 23751 4129
rect 23693 4120 23705 4123
rect 23656 4092 23705 4120
rect 23656 4080 23662 4092
rect 23693 4089 23705 4092
rect 23739 4120 23751 4123
rect 25346 4120 25352 4132
rect 23739 4092 25352 4120
rect 23739 4089 23751 4092
rect 23693 4083 23751 4089
rect 25346 4080 25352 4092
rect 25404 4080 25410 4132
rect 1334 4012 1340 4064
rect 1392 4052 1398 4064
rect 2257 4055 2315 4061
rect 2257 4052 2269 4055
rect 1392 4024 2269 4052
rect 1392 4012 1398 4024
rect 2257 4021 2269 4024
rect 2303 4052 2315 4055
rect 2714 4052 2720 4064
rect 2303 4024 2720 4052
rect 2303 4021 2315 4024
rect 2257 4015 2315 4021
rect 2714 4012 2720 4024
rect 2772 4012 2778 4064
rect 3266 4012 3272 4064
rect 3324 4052 3330 4064
rect 3361 4055 3419 4061
rect 3361 4052 3373 4055
rect 3324 4024 3373 4052
rect 3324 4012 3330 4024
rect 3361 4021 3373 4024
rect 3407 4021 3419 4055
rect 3361 4015 3419 4021
rect 14490 4012 14496 4064
rect 14548 4052 14554 4064
rect 15226 4052 15232 4064
rect 14548 4024 15232 4052
rect 14548 4012 14554 4024
rect 15226 4012 15232 4024
rect 15284 4052 15290 4064
rect 15505 4055 15563 4061
rect 15505 4052 15517 4055
rect 15284 4024 15517 4052
rect 15284 4012 15290 4024
rect 15505 4021 15517 4024
rect 15551 4021 15563 4055
rect 15505 4015 15563 4021
rect 15962 4012 15968 4064
rect 16020 4012 16026 4064
rect 22589 4055 22647 4061
rect 22589 4021 22601 4055
rect 22635 4052 22647 4055
rect 22678 4052 22684 4064
rect 22635 4024 22684 4052
rect 22635 4021 22647 4024
rect 22589 4015 22647 4021
rect 22678 4012 22684 4024
rect 22736 4012 22742 4064
rect 693 3987 751 3993
rect 693 3953 705 3987
rect 739 3984 751 3987
rect 782 3984 788 3996
rect 739 3956 788 3984
rect 739 3953 751 3956
rect 693 3947 751 3953
rect 782 3944 788 3956
rect 840 3984 846 3996
rect 1242 3984 1248 3996
rect 840 3956 1248 3984
rect 840 3944 846 3956
rect 1242 3944 1248 3956
rect 1300 3944 1306 3996
rect 1518 3944 1524 3996
rect 1576 3984 1582 3996
rect 1613 3987 1671 3993
rect 1613 3984 1625 3987
rect 1576 3956 1625 3984
rect 1576 3944 1582 3956
rect 1613 3953 1625 3956
rect 1659 3953 1671 3987
rect 1613 3947 1671 3953
rect 3545 3987 3603 3993
rect 3545 3953 3557 3987
rect 3591 3953 3603 3987
rect 9154 3984 9160 3996
rect 9115 3956 9160 3984
rect 3545 3947 3603 3953
rect 3358 3876 3364 3928
rect 3416 3916 3422 3928
rect 3560 3916 3588 3947
rect 9154 3944 9160 3956
rect 9212 3944 9218 3996
rect 22770 3984 22776 3996
rect 22731 3956 22776 3984
rect 22770 3944 22776 3956
rect 22828 3944 22834 3996
rect 3416 3888 3588 3916
rect 15229 3919 15287 3925
rect 3416 3876 3422 3888
rect 15229 3885 15241 3919
rect 15275 3916 15287 3919
rect 15502 3916 15508 3928
rect 15275 3888 15508 3916
rect 15275 3885 15287 3888
rect 15229 3879 15287 3885
rect 15502 3876 15508 3888
rect 15560 3876 15566 3928
rect 15870 3876 15876 3928
rect 15928 3916 15934 3928
rect 17066 3916 17072 3928
rect 15928 3888 17072 3916
rect 15928 3876 15934 3888
rect 17066 3876 17072 3888
rect 17124 3916 17130 3928
rect 17253 3919 17311 3925
rect 17253 3916 17265 3919
rect 17124 3888 17265 3916
rect 17124 3876 17130 3888
rect 17253 3885 17265 3888
rect 17299 3885 17311 3919
rect 17253 3879 17311 3885
rect 2438 3808 2444 3860
rect 2496 3848 2502 3860
rect 3729 3851 3787 3857
rect 3729 3848 3741 3851
rect 2496 3820 3741 3848
rect 2496 3808 2502 3820
rect 3729 3817 3741 3820
rect 3775 3848 3787 3851
rect 3910 3848 3916 3860
rect 3775 3820 3916 3848
rect 3775 3817 3787 3820
rect 3729 3811 3787 3817
rect 3910 3808 3916 3820
rect 3968 3808 3974 3860
rect 9154 3780 9160 3792
rect 9115 3752 9160 3780
rect 9154 3740 9160 3752
rect 9212 3740 9218 3792
rect 22494 3740 22500 3792
rect 22552 3780 22558 3792
rect 22865 3783 22923 3789
rect 22865 3780 22877 3783
rect 22552 3752 22877 3780
rect 22552 3740 22558 3752
rect 22865 3749 22877 3752
rect 22911 3749 22923 3783
rect 22865 3743 22923 3749
rect 23874 3740 23880 3792
rect 23932 3780 23938 3792
rect 24061 3783 24119 3789
rect 23932 3752 23977 3780
rect 23932 3740 23938 3752
rect 24061 3749 24073 3783
rect 24107 3780 24119 3783
rect 24334 3780 24340 3792
rect 24107 3752 24340 3780
rect 24107 3749 24119 3752
rect 24061 3743 24119 3749
rect 24334 3740 24340 3752
rect 24392 3740 24398 3792
rect 400 3690 27264 3712
rect 400 3638 3510 3690
rect 3562 3638 3574 3690
rect 3626 3638 3638 3690
rect 3690 3638 3702 3690
rect 3754 3638 3766 3690
rect 3818 3638 27264 3690
rect 400 3616 27264 3638
rect 782 3576 788 3588
rect 743 3548 788 3576
rect 782 3536 788 3548
rect 840 3536 846 3588
rect 3266 3536 3272 3588
rect 3324 3576 3330 3588
rect 3545 3579 3603 3585
rect 3545 3576 3557 3579
rect 3324 3548 3557 3576
rect 3324 3536 3330 3548
rect 3545 3545 3557 3548
rect 3591 3545 3603 3579
rect 3545 3539 3603 3545
rect 3821 3579 3879 3585
rect 3821 3545 3833 3579
rect 3867 3576 3879 3579
rect 3910 3576 3916 3588
rect 3867 3548 3916 3576
rect 3867 3545 3879 3548
rect 3821 3539 3879 3545
rect 3910 3536 3916 3548
rect 3968 3536 3974 3588
rect 4002 3536 4008 3588
rect 4060 3576 4066 3588
rect 4557 3579 4615 3585
rect 4557 3576 4569 3579
rect 4060 3548 4569 3576
rect 4060 3536 4066 3548
rect 4557 3545 4569 3548
rect 4603 3545 4615 3579
rect 4557 3539 4615 3545
rect 8421 3579 8479 3585
rect 8421 3545 8433 3579
rect 8467 3576 8479 3579
rect 8605 3579 8663 3585
rect 8605 3576 8617 3579
rect 8467 3548 8617 3576
rect 8467 3545 8479 3548
rect 8421 3539 8479 3545
rect 8605 3545 8617 3548
rect 8651 3576 8663 3579
rect 8694 3576 8700 3588
rect 8651 3548 8700 3576
rect 8651 3545 8663 3548
rect 8605 3539 8663 3545
rect 800 3440 828 3536
rect 1334 3508 1340 3520
rect 1295 3480 1340 3508
rect 1334 3468 1340 3480
rect 1392 3468 1398 3520
rect 4572 3508 4600 3539
rect 8694 3536 8700 3548
rect 8752 3536 8758 3588
rect 15226 3576 15232 3588
rect 15187 3548 15232 3576
rect 15226 3536 15232 3548
rect 15284 3536 15290 3588
rect 15870 3576 15876 3588
rect 15831 3548 15876 3576
rect 15870 3536 15876 3548
rect 15928 3536 15934 3588
rect 21022 3576 21028 3588
rect 20983 3548 21028 3576
rect 21022 3536 21028 3548
rect 21080 3536 21086 3588
rect 22494 3576 22500 3588
rect 22455 3548 22500 3576
rect 22494 3536 22500 3548
rect 22552 3536 22558 3588
rect 22770 3536 22776 3588
rect 22828 3576 22834 3588
rect 22957 3579 23015 3585
rect 22957 3576 22969 3579
rect 22828 3548 22969 3576
rect 22828 3536 22834 3548
rect 22957 3545 22969 3548
rect 23003 3545 23015 3579
rect 22957 3539 23015 3545
rect 4925 3511 4983 3517
rect 4925 3508 4937 3511
rect 4572 3480 4937 3508
rect 4925 3477 4937 3480
rect 4971 3508 4983 3511
rect 9062 3508 9068 3520
rect 4971 3480 9068 3508
rect 4971 3477 4983 3480
rect 4925 3471 4983 3477
rect 9062 3468 9068 3480
rect 9120 3468 9126 3520
rect 15505 3511 15563 3517
rect 15505 3477 15517 3511
rect 15551 3508 15563 3511
rect 15962 3508 15968 3520
rect 15551 3480 15968 3508
rect 15551 3477 15563 3480
rect 15505 3471 15563 3477
rect 15962 3468 15968 3480
rect 16020 3508 16026 3520
rect 16020 3480 17572 3508
rect 16020 3468 16026 3480
rect 17544 3449 17572 3480
rect 877 3443 935 3449
rect 877 3440 889 3443
rect 800 3412 889 3440
rect 877 3409 889 3412
rect 923 3440 935 3443
rect 1521 3443 1579 3449
rect 1521 3440 1533 3443
rect 923 3412 1533 3440
rect 923 3409 935 3412
rect 877 3403 935 3409
rect 1521 3409 1533 3412
rect 1567 3409 1579 3443
rect 5661 3443 5719 3449
rect 5661 3440 5673 3443
rect 1521 3403 1579 3409
rect 4480 3412 5673 3440
rect 3358 3332 3364 3384
rect 3416 3372 3422 3384
rect 4189 3375 4247 3381
rect 4189 3372 4201 3375
rect 3416 3344 4201 3372
rect 3416 3332 3422 3344
rect 4189 3341 4201 3344
rect 4235 3341 4247 3375
rect 4189 3335 4247 3341
rect 1429 3307 1487 3313
rect 1429 3273 1441 3307
rect 1475 3304 1487 3307
rect 1610 3304 1616 3316
rect 1475 3276 1616 3304
rect 1475 3273 1487 3276
rect 1429 3267 1487 3273
rect 1610 3264 1616 3276
rect 1668 3304 1674 3316
rect 1705 3307 1763 3313
rect 1705 3304 1717 3307
rect 1668 3276 1717 3304
rect 1668 3264 1674 3276
rect 1705 3273 1717 3276
rect 1751 3273 1763 3307
rect 4204 3304 4232 3335
rect 4480 3304 4508 3412
rect 5661 3409 5673 3412
rect 5707 3440 5719 3443
rect 17529 3443 17587 3449
rect 5707 3412 6624 3440
rect 5707 3409 5719 3412
rect 5661 3403 5719 3409
rect 4557 3375 4615 3381
rect 4557 3341 4569 3375
rect 4603 3372 4615 3375
rect 6118 3372 6124 3384
rect 4603 3344 5152 3372
rect 6079 3344 6124 3372
rect 4603 3341 4615 3344
rect 4557 3335 4615 3341
rect 4649 3307 4707 3313
rect 4649 3304 4661 3307
rect 4204 3276 4661 3304
rect 1705 3267 1763 3273
rect 4649 3273 4661 3276
rect 4695 3273 4707 3307
rect 4649 3267 4707 3273
rect 5124 3248 5152 3344
rect 6118 3332 6124 3344
rect 6176 3332 6182 3384
rect 6596 3381 6624 3412
rect 17529 3409 17541 3443
rect 17575 3440 17587 3443
rect 18081 3443 18139 3449
rect 18081 3440 18093 3443
rect 17575 3412 18093 3440
rect 17575 3409 17587 3412
rect 17529 3403 17587 3409
rect 18081 3409 18093 3412
rect 18127 3409 18139 3443
rect 22972 3440 23000 3539
rect 23874 3536 23880 3588
rect 23932 3576 23938 3588
rect 25303 3579 25361 3585
rect 25303 3576 25315 3579
rect 23932 3548 25315 3576
rect 23932 3536 23938 3548
rect 25303 3545 25315 3548
rect 25349 3545 25361 3579
rect 25303 3539 25361 3545
rect 23874 3440 23880 3452
rect 22972 3412 23880 3440
rect 18081 3403 18139 3409
rect 23874 3400 23880 3412
rect 23932 3400 23938 3452
rect 6581 3375 6639 3381
rect 6581 3341 6593 3375
rect 6627 3341 6639 3375
rect 6581 3335 6639 3341
rect 8237 3375 8295 3381
rect 8237 3341 8249 3375
rect 8283 3372 8295 3375
rect 9154 3372 9160 3384
rect 8283 3344 9160 3372
rect 8283 3341 8295 3344
rect 8237 3335 8295 3341
rect 9154 3332 9160 3344
rect 9212 3372 9218 3384
rect 9433 3375 9491 3381
rect 9433 3372 9445 3375
rect 9212 3344 9445 3372
rect 9212 3332 9218 3344
rect 9433 3341 9445 3344
rect 9479 3372 9491 3375
rect 9709 3375 9767 3381
rect 9709 3372 9721 3375
rect 9479 3344 9721 3372
rect 9479 3341 9491 3344
rect 9433 3335 9491 3341
rect 9709 3341 9721 3344
rect 9755 3341 9767 3375
rect 9709 3335 9767 3341
rect 12374 3332 12380 3384
rect 12432 3372 12438 3384
rect 17345 3375 17403 3381
rect 17345 3372 17357 3375
rect 12432 3344 17357 3372
rect 12432 3332 12438 3344
rect 17345 3341 17357 3344
rect 17391 3372 17403 3375
rect 17894 3372 17900 3384
rect 17391 3344 17900 3372
rect 17391 3341 17403 3344
rect 17345 3335 17403 3341
rect 17894 3332 17900 3344
rect 17952 3332 17958 3384
rect 23598 3372 23604 3384
rect 23559 3344 23604 3372
rect 23598 3332 23604 3344
rect 23656 3332 23662 3384
rect 6136 3304 6164 3332
rect 6949 3307 7007 3313
rect 6949 3304 6961 3307
rect 6136 3276 6961 3304
rect 6949 3273 6961 3276
rect 6995 3273 7007 3307
rect 6949 3267 7007 3273
rect 11917 3307 11975 3313
rect 11917 3273 11929 3307
rect 11963 3304 11975 3307
rect 12193 3307 12251 3313
rect 12193 3304 12205 3307
rect 11963 3276 12205 3304
rect 11963 3273 11975 3276
rect 11917 3267 11975 3273
rect 12193 3273 12205 3276
rect 12239 3304 12251 3307
rect 12466 3304 12472 3316
rect 12239 3276 12472 3304
rect 12239 3273 12251 3276
rect 12193 3267 12251 3273
rect 12466 3264 12472 3276
rect 12524 3264 12530 3316
rect 15502 3264 15508 3316
rect 15560 3304 15566 3316
rect 15689 3307 15747 3313
rect 15689 3304 15701 3307
rect 15560 3276 15701 3304
rect 15560 3264 15566 3276
rect 15689 3273 15701 3276
rect 15735 3304 15747 3307
rect 17986 3304 17992 3316
rect 15735 3276 17992 3304
rect 15735 3273 15747 3276
rect 15689 3267 15747 3273
rect 17986 3264 17992 3276
rect 18044 3264 18050 3316
rect 23877 3307 23935 3313
rect 23877 3273 23889 3307
rect 23923 3304 23935 3307
rect 23923 3276 23957 3304
rect 23923 3273 23935 3276
rect 23877 3267 23935 3273
rect 3266 3196 3272 3248
rect 3324 3236 3330 3248
rect 3361 3239 3419 3245
rect 3361 3236 3373 3239
rect 3324 3208 3373 3236
rect 3324 3196 3330 3208
rect 3361 3205 3373 3208
rect 3407 3205 3419 3239
rect 5106 3236 5112 3248
rect 5067 3208 5112 3236
rect 3361 3199 3419 3205
rect 5106 3196 5112 3208
rect 5164 3196 5170 3248
rect 5937 3239 5995 3245
rect 5937 3205 5949 3239
rect 5983 3236 5995 3239
rect 6210 3236 6216 3248
rect 5983 3208 6216 3236
rect 5983 3205 5995 3208
rect 5937 3199 5995 3205
rect 6210 3196 6216 3208
rect 6268 3196 6274 3248
rect 11362 3196 11368 3248
rect 11420 3236 11426 3248
rect 11733 3239 11791 3245
rect 11733 3236 11745 3239
rect 11420 3208 11745 3236
rect 11420 3196 11426 3208
rect 11733 3205 11745 3208
rect 11779 3236 11791 3239
rect 12009 3239 12067 3245
rect 12009 3236 12021 3239
rect 11779 3208 12021 3236
rect 11779 3205 11791 3208
rect 11733 3199 11791 3205
rect 12009 3205 12021 3208
rect 12055 3205 12067 3239
rect 22678 3236 22684 3248
rect 22639 3208 22684 3236
rect 12009 3199 12067 3205
rect 22678 3196 22684 3208
rect 22736 3196 22742 3248
rect 23325 3239 23383 3245
rect 23325 3205 23337 3239
rect 23371 3236 23383 3239
rect 23506 3236 23512 3248
rect 23371 3208 23512 3236
rect 23371 3205 23383 3208
rect 23325 3199 23383 3205
rect 23506 3196 23512 3208
rect 23564 3236 23570 3248
rect 23892 3236 23920 3267
rect 24334 3264 24340 3316
rect 24392 3264 24398 3316
rect 25625 3239 25683 3245
rect 25625 3236 25637 3239
rect 23564 3208 25637 3236
rect 23564 3196 23570 3208
rect 25625 3205 25637 3208
rect 25671 3205 25683 3239
rect 25625 3199 25683 3205
rect 400 3146 27264 3168
rect 400 3094 18870 3146
rect 18922 3094 18934 3146
rect 18986 3094 18998 3146
rect 19050 3094 19062 3146
rect 19114 3094 19126 3146
rect 19178 3094 27264 3146
rect 400 3072 27264 3094
rect 785 3035 843 3041
rect 785 3001 797 3035
rect 831 3032 843 3035
rect 969 3035 1027 3041
rect 969 3032 981 3035
rect 831 3004 981 3032
rect 831 3001 843 3004
rect 785 2995 843 3001
rect 969 3001 981 3004
rect 1015 3032 1027 3035
rect 1334 3032 1340 3044
rect 1015 3004 1340 3032
rect 1015 3001 1027 3004
rect 969 2995 1027 3001
rect 1334 2992 1340 3004
rect 1392 2992 1398 3044
rect 9062 3032 9068 3044
rect 9023 3004 9068 3032
rect 9062 2992 9068 3004
rect 9120 2992 9126 3044
rect 22678 2992 22684 3044
rect 22736 3032 22742 3044
rect 24150 3032 24156 3044
rect 22736 3004 24156 3032
rect 22736 2992 22742 3004
rect 24150 2992 24156 3004
rect 24208 3032 24214 3044
rect 24245 3035 24303 3041
rect 24245 3032 24257 3035
rect 24208 3004 24257 3032
rect 24208 2992 24214 3004
rect 24245 3001 24257 3004
rect 24291 3032 24303 3035
rect 25254 3032 25260 3044
rect 24291 3004 25260 3032
rect 24291 3001 24303 3004
rect 24245 2995 24303 3001
rect 25254 2992 25260 3004
rect 25312 2992 25318 3044
rect 1610 2964 1616 2976
rect 1571 2936 1616 2964
rect 1610 2924 1616 2936
rect 1668 2964 1674 2976
rect 1705 2967 1763 2973
rect 1705 2964 1717 2967
rect 1668 2936 1717 2964
rect 1668 2924 1674 2936
rect 1705 2933 1717 2936
rect 1751 2933 1763 2967
rect 18078 2964 18084 2976
rect 18039 2936 18084 2964
rect 1705 2927 1763 2933
rect 18078 2924 18084 2936
rect 18136 2924 18142 2976
rect 20930 2924 20936 2976
rect 20988 2964 20994 2976
rect 20988 2936 21528 2964
rect 20988 2924 20994 2936
rect 1426 2896 1432 2908
rect 1387 2868 1432 2896
rect 1426 2856 1432 2868
rect 1484 2856 1490 2908
rect 4465 2899 4523 2905
rect 4465 2865 4477 2899
rect 4511 2896 4523 2899
rect 5106 2896 5112 2908
rect 4511 2868 5112 2896
rect 4511 2865 4523 2868
rect 4465 2859 4523 2865
rect 5106 2856 5112 2868
rect 5164 2856 5170 2908
rect 6670 2856 6676 2908
rect 6728 2896 6734 2908
rect 6949 2899 7007 2905
rect 6949 2896 6961 2899
rect 6728 2868 6961 2896
rect 6728 2856 6734 2868
rect 6949 2865 6961 2868
rect 6995 2896 7007 2899
rect 10258 2896 10264 2908
rect 6995 2868 10264 2896
rect 6995 2865 7007 2868
rect 6949 2859 7007 2865
rect 10258 2856 10264 2868
rect 10316 2856 10322 2908
rect 11733 2899 11791 2905
rect 11733 2865 11745 2899
rect 11779 2896 11791 2899
rect 11822 2896 11828 2908
rect 11779 2868 11828 2896
rect 11779 2865 11791 2868
rect 11733 2859 11791 2865
rect 11822 2856 11828 2868
rect 11880 2856 11886 2908
rect 13202 2896 13208 2908
rect 13115 2868 13208 2896
rect 13202 2856 13208 2868
rect 13260 2896 13266 2908
rect 14030 2896 14036 2908
rect 13260 2868 14036 2896
rect 13260 2856 13266 2868
rect 14030 2856 14036 2868
rect 14088 2856 14094 2908
rect 14398 2856 14404 2908
rect 14456 2896 14462 2908
rect 15505 2899 15563 2905
rect 15505 2896 15517 2899
rect 14456 2868 15517 2896
rect 14456 2856 14462 2868
rect 15505 2865 15517 2868
rect 15551 2896 15563 2899
rect 15962 2896 15968 2908
rect 15551 2868 15968 2896
rect 15551 2865 15563 2868
rect 15505 2859 15563 2865
rect 15962 2856 15968 2868
rect 16020 2856 16026 2908
rect 18630 2856 18636 2908
rect 18688 2896 18694 2908
rect 21500 2905 21528 2936
rect 18817 2899 18875 2905
rect 18817 2896 18829 2899
rect 18688 2868 18829 2896
rect 18688 2856 18694 2868
rect 18817 2865 18829 2868
rect 18863 2865 18875 2899
rect 18817 2859 18875 2865
rect 21393 2899 21451 2905
rect 21393 2865 21405 2899
rect 21439 2865 21451 2899
rect 21393 2859 21451 2865
rect 21485 2899 21543 2905
rect 21485 2865 21497 2899
rect 21531 2865 21543 2899
rect 22126 2896 22132 2908
rect 22087 2868 22132 2896
rect 21485 2859 21543 2865
rect 1153 2831 1211 2837
rect 1153 2797 1165 2831
rect 1199 2828 1211 2831
rect 1518 2828 1524 2840
rect 1199 2800 1524 2828
rect 1199 2797 1211 2800
rect 1153 2791 1211 2797
rect 1518 2788 1524 2800
rect 1576 2788 1582 2840
rect 7498 2828 7504 2840
rect 7459 2800 7504 2828
rect 7498 2788 7504 2800
rect 7556 2788 7562 2840
rect 13294 2828 13300 2840
rect 13255 2800 13300 2828
rect 13294 2788 13300 2800
rect 13352 2788 13358 2840
rect 14950 2828 14956 2840
rect 14911 2800 14956 2828
rect 14950 2788 14956 2800
rect 15008 2788 15014 2840
rect 17986 2828 17992 2840
rect 17947 2800 17992 2828
rect 17986 2788 17992 2800
rect 18044 2788 18050 2840
rect 18170 2788 18176 2840
rect 18228 2828 18234 2840
rect 18909 2831 18967 2837
rect 18909 2828 18921 2831
rect 18228 2800 18921 2828
rect 18228 2788 18234 2800
rect 18909 2797 18921 2800
rect 18955 2797 18967 2831
rect 20470 2828 20476 2840
rect 20383 2800 20476 2828
rect 18909 2791 18967 2797
rect 20470 2788 20476 2800
rect 20528 2828 20534 2840
rect 21117 2831 21175 2837
rect 21117 2828 21129 2831
rect 20528 2800 21129 2828
rect 20528 2788 20534 2800
rect 21117 2797 21129 2800
rect 21163 2797 21175 2831
rect 21408 2828 21436 2859
rect 22126 2856 22132 2868
rect 22184 2856 22190 2908
rect 22402 2896 22408 2908
rect 22363 2868 22408 2896
rect 22402 2856 22408 2868
rect 22460 2856 22466 2908
rect 23506 2896 23512 2908
rect 23467 2868 23512 2896
rect 23506 2856 23512 2868
rect 23564 2856 23570 2908
rect 23693 2899 23751 2905
rect 23693 2865 23705 2899
rect 23739 2896 23751 2899
rect 23874 2896 23880 2908
rect 23739 2868 23880 2896
rect 23739 2865 23751 2868
rect 23693 2859 23751 2865
rect 23874 2856 23880 2868
rect 23932 2856 23938 2908
rect 22494 2828 22500 2840
rect 21408 2800 22500 2828
rect 21117 2791 21175 2797
rect 22494 2788 22500 2800
rect 22552 2788 22558 2840
rect 7409 2763 7467 2769
rect 7409 2729 7421 2763
rect 7455 2729 7467 2763
rect 7409 2723 7467 2729
rect 15413 2763 15471 2769
rect 15413 2729 15425 2763
rect 15459 2729 15471 2763
rect 15413 2723 15471 2729
rect 20657 2763 20715 2769
rect 20657 2729 20669 2763
rect 20703 2760 20715 2763
rect 20746 2760 20752 2772
rect 20703 2732 20752 2760
rect 20703 2729 20715 2732
rect 20657 2723 20715 2729
rect 4738 2652 4744 2704
rect 4796 2692 4802 2704
rect 6765 2695 6823 2701
rect 6765 2692 6777 2695
rect 4796 2664 6777 2692
rect 4796 2652 4802 2664
rect 6765 2661 6777 2664
rect 6811 2692 6823 2695
rect 7130 2692 7136 2704
rect 6811 2664 7136 2692
rect 6811 2661 6823 2664
rect 6765 2655 6823 2661
rect 7130 2652 7136 2664
rect 7188 2692 7194 2704
rect 7424 2692 7452 2723
rect 7188 2664 7452 2692
rect 9985 2695 10043 2701
rect 7188 2652 7194 2664
rect 9985 2661 9997 2695
rect 10031 2692 10043 2695
rect 10810 2692 10816 2704
rect 10031 2664 10816 2692
rect 10031 2661 10043 2664
rect 9985 2655 10043 2661
rect 10810 2652 10816 2664
rect 10868 2652 10874 2704
rect 15428 2692 15456 2723
rect 20746 2720 20752 2732
rect 20804 2720 20810 2772
rect 15686 2692 15692 2704
rect 15428 2664 15692 2692
rect 15686 2652 15692 2664
rect 15744 2652 15750 2704
rect 22402 2652 22408 2704
rect 22460 2692 22466 2704
rect 23785 2695 23843 2701
rect 23785 2692 23797 2695
rect 22460 2664 23797 2692
rect 22460 2652 22466 2664
rect 23785 2661 23797 2664
rect 23831 2692 23843 2695
rect 24058 2692 24064 2704
rect 23831 2664 24064 2692
rect 23831 2661 23843 2664
rect 23785 2655 23843 2661
rect 24058 2652 24064 2664
rect 24116 2652 24122 2704
rect 24426 2692 24432 2704
rect 24387 2664 24432 2692
rect 24426 2652 24432 2664
rect 24484 2652 24490 2704
rect 400 2602 27264 2624
rect 400 2550 3510 2602
rect 3562 2550 3574 2602
rect 3626 2550 3638 2602
rect 3690 2550 3702 2602
rect 3754 2550 3766 2602
rect 3818 2550 27264 2602
rect 400 2528 27264 2550
rect 1518 2448 1524 2500
rect 1576 2488 1582 2500
rect 2349 2491 2407 2497
rect 2349 2488 2361 2491
rect 1576 2460 2361 2488
rect 1576 2448 1582 2460
rect 877 2355 935 2361
rect 877 2321 889 2355
rect 923 2352 935 2355
rect 1061 2355 1119 2361
rect 1061 2352 1073 2355
rect 923 2324 1073 2352
rect 923 2321 935 2324
rect 877 2315 935 2321
rect 1061 2321 1073 2324
rect 1107 2352 1119 2355
rect 1426 2352 1432 2364
rect 1107 2324 1432 2352
rect 1107 2321 1119 2324
rect 1061 2315 1119 2321
rect 1426 2312 1432 2324
rect 1484 2352 1490 2364
rect 1484 2324 1656 2352
rect 1484 2312 1490 2324
rect 1337 2287 1395 2293
rect 1337 2253 1349 2287
rect 1383 2253 1395 2287
rect 1337 2247 1395 2253
rect 1352 2160 1380 2247
rect 1628 2228 1656 2324
rect 2272 2293 2300 2460
rect 2349 2457 2361 2460
rect 2395 2457 2407 2491
rect 5106 2488 5112 2500
rect 5067 2460 5112 2488
rect 2349 2451 2407 2457
rect 5106 2448 5112 2460
rect 5164 2448 5170 2500
rect 6489 2491 6547 2497
rect 6489 2457 6501 2491
rect 6535 2488 6547 2491
rect 6670 2488 6676 2500
rect 6535 2460 6676 2488
rect 6535 2457 6547 2460
rect 6489 2451 6547 2457
rect 6670 2448 6676 2460
rect 6728 2448 6734 2500
rect 11822 2488 11828 2500
rect 11783 2460 11828 2488
rect 11822 2448 11828 2460
rect 11880 2488 11886 2500
rect 12561 2491 12619 2497
rect 12561 2488 12573 2491
rect 11880 2460 12573 2488
rect 11880 2448 11886 2460
rect 12561 2457 12573 2460
rect 12607 2457 12619 2491
rect 14398 2488 14404 2500
rect 14359 2460 14404 2488
rect 12561 2451 12619 2457
rect 14398 2448 14404 2460
rect 14456 2448 14462 2500
rect 14585 2491 14643 2497
rect 14585 2457 14597 2491
rect 14631 2488 14643 2491
rect 14769 2491 14827 2497
rect 14769 2488 14781 2491
rect 14631 2460 14781 2488
rect 14631 2457 14643 2460
rect 14585 2451 14643 2457
rect 14769 2457 14781 2460
rect 14815 2488 14827 2491
rect 14950 2488 14956 2500
rect 14815 2460 14956 2488
rect 14815 2457 14827 2460
rect 14769 2451 14827 2457
rect 7130 2380 7136 2432
rect 7188 2420 7194 2432
rect 8053 2423 8111 2429
rect 8053 2420 8065 2423
rect 7188 2392 8065 2420
rect 7188 2380 7194 2392
rect 8053 2389 8065 2392
rect 8099 2389 8111 2423
rect 8053 2383 8111 2389
rect 9617 2355 9675 2361
rect 3560 2324 4692 2352
rect 3560 2293 3588 2324
rect 2257 2287 2315 2293
rect 2257 2253 2269 2287
rect 2303 2284 2315 2287
rect 3269 2287 3327 2293
rect 3269 2284 3281 2287
rect 2303 2256 3281 2284
rect 2303 2253 2315 2256
rect 2257 2247 2315 2253
rect 3269 2253 3281 2256
rect 3315 2284 3327 2287
rect 3545 2287 3603 2293
rect 3545 2284 3557 2287
rect 3315 2256 3557 2284
rect 3315 2253 3327 2256
rect 3269 2247 3327 2253
rect 3545 2253 3557 2256
rect 3591 2253 3603 2287
rect 3545 2247 3603 2253
rect 1610 2176 1616 2228
rect 1668 2216 1674 2228
rect 4664 2225 4692 2324
rect 9617 2321 9629 2355
rect 9663 2352 9675 2355
rect 11840 2352 11868 2448
rect 13754 2380 13760 2432
rect 13812 2420 13818 2432
rect 14600 2420 14628 2451
rect 13812 2392 14628 2420
rect 13812 2380 13818 2392
rect 11917 2355 11975 2361
rect 11917 2352 11929 2355
rect 9663 2324 10672 2352
rect 11840 2324 11929 2352
rect 9663 2321 9675 2324
rect 9617 2315 9675 2321
rect 6670 2244 6676 2296
rect 6728 2284 6734 2296
rect 6765 2287 6823 2293
rect 6765 2284 6777 2287
rect 6728 2256 6777 2284
rect 6728 2244 6734 2256
rect 6765 2253 6777 2256
rect 6811 2253 6823 2287
rect 7774 2284 7780 2296
rect 7735 2256 7780 2284
rect 6765 2247 6823 2253
rect 7774 2244 7780 2256
rect 7832 2244 7838 2296
rect 10644 2293 10672 2324
rect 11917 2321 11929 2324
rect 11963 2321 11975 2355
rect 12466 2352 12472 2364
rect 12427 2324 12472 2352
rect 11917 2315 11975 2321
rect 12466 2312 12472 2324
rect 12524 2352 12530 2364
rect 12745 2355 12803 2361
rect 12745 2352 12757 2355
rect 12524 2324 12757 2352
rect 12524 2312 12530 2324
rect 12745 2321 12757 2324
rect 12791 2321 12803 2355
rect 12745 2315 12803 2321
rect 9893 2287 9951 2293
rect 9893 2253 9905 2287
rect 9939 2253 9951 2287
rect 9893 2247 9951 2253
rect 10629 2287 10687 2293
rect 10629 2253 10641 2287
rect 10675 2284 10687 2287
rect 11270 2284 11276 2296
rect 10675 2256 11276 2284
rect 10675 2253 10687 2256
rect 10629 2247 10687 2253
rect 1981 2219 2039 2225
rect 1981 2216 1993 2219
rect 1668 2188 1993 2216
rect 1668 2176 1674 2188
rect 1981 2185 1993 2188
rect 2027 2185 2039 2219
rect 1981 2179 2039 2185
rect 4465 2219 4523 2225
rect 4465 2185 4477 2219
rect 4511 2216 4523 2219
rect 4649 2219 4707 2225
rect 4511 2188 4600 2216
rect 4511 2185 4523 2188
rect 4465 2179 4523 2185
rect 1245 2151 1303 2157
rect 1245 2117 1257 2151
rect 1291 2148 1303 2151
rect 1334 2148 1340 2160
rect 1291 2120 1340 2148
rect 1291 2117 1303 2120
rect 1245 2111 1303 2117
rect 1334 2108 1340 2120
rect 1392 2108 1398 2160
rect 3082 2148 3088 2160
rect 3043 2120 3088 2148
rect 3082 2108 3088 2120
rect 3140 2148 3146 2160
rect 3361 2151 3419 2157
rect 3361 2148 3373 2151
rect 3140 2120 3373 2148
rect 3140 2108 3146 2120
rect 3361 2117 3373 2120
rect 3407 2117 3419 2151
rect 4572 2148 4600 2188
rect 4649 2185 4661 2219
rect 4695 2216 4707 2219
rect 4925 2219 4983 2225
rect 4925 2216 4937 2219
rect 4695 2188 4937 2216
rect 4695 2185 4707 2188
rect 4649 2179 4707 2185
rect 4925 2185 4937 2188
rect 4971 2185 4983 2219
rect 4925 2179 4983 2185
rect 4738 2148 4744 2160
rect 4572 2120 4744 2148
rect 3361 2111 3419 2117
rect 4738 2108 4744 2120
rect 4796 2108 4802 2160
rect 6210 2148 6216 2160
rect 6171 2120 6216 2148
rect 6210 2108 6216 2120
rect 6268 2108 6274 2160
rect 9798 2148 9804 2160
rect 9711 2120 9804 2148
rect 9798 2108 9804 2120
rect 9856 2148 9862 2160
rect 9908 2148 9936 2247
rect 11270 2244 11276 2256
rect 11328 2244 11334 2296
rect 12377 2287 12435 2293
rect 12377 2253 12389 2287
rect 12423 2284 12435 2287
rect 13294 2284 13300 2296
rect 12423 2256 13300 2284
rect 12423 2253 12435 2256
rect 12377 2247 12435 2253
rect 10810 2216 10816 2228
rect 10771 2188 10816 2216
rect 10810 2176 10816 2188
rect 10868 2176 10874 2228
rect 11365 2219 11423 2225
rect 11365 2185 11377 2219
rect 11411 2216 11423 2219
rect 11549 2219 11607 2225
rect 11549 2216 11561 2219
rect 11411 2188 11561 2216
rect 11411 2185 11423 2188
rect 11365 2179 11423 2185
rect 11549 2185 11561 2188
rect 11595 2216 11607 2219
rect 12392 2216 12420 2247
rect 13294 2244 13300 2256
rect 13352 2284 13358 2296
rect 14876 2293 14904 2460
rect 14950 2448 14956 2460
rect 15008 2448 15014 2500
rect 17434 2488 17440 2500
rect 17395 2460 17440 2488
rect 17434 2448 17440 2460
rect 17492 2488 17498 2500
rect 17621 2491 17679 2497
rect 17621 2488 17633 2491
rect 17492 2460 17633 2488
rect 17492 2448 17498 2460
rect 17621 2457 17633 2460
rect 17667 2457 17679 2491
rect 17621 2451 17679 2457
rect 17897 2491 17955 2497
rect 17897 2457 17909 2491
rect 17943 2488 17955 2491
rect 18078 2488 18084 2500
rect 17943 2460 18084 2488
rect 17943 2457 17955 2460
rect 17897 2451 17955 2457
rect 18078 2448 18084 2460
rect 18136 2448 18142 2500
rect 22126 2488 22132 2500
rect 22087 2460 22132 2488
rect 22126 2448 22132 2460
rect 22184 2448 22190 2500
rect 22313 2491 22371 2497
rect 22313 2457 22325 2491
rect 22359 2488 22371 2491
rect 22494 2488 22500 2500
rect 22359 2460 22500 2488
rect 22359 2457 22371 2460
rect 22313 2451 22371 2457
rect 22494 2448 22500 2460
rect 22552 2448 22558 2500
rect 23598 2448 23604 2500
rect 23656 2488 23662 2500
rect 23785 2491 23843 2497
rect 23785 2488 23797 2491
rect 23656 2460 23797 2488
rect 23656 2448 23662 2460
rect 23785 2457 23797 2460
rect 23831 2488 23843 2491
rect 23969 2491 24027 2497
rect 23969 2488 23981 2491
rect 23831 2460 23981 2488
rect 23831 2457 23843 2460
rect 23785 2451 23843 2457
rect 23969 2457 23981 2460
rect 24015 2488 24027 2491
rect 24015 2460 24288 2488
rect 24015 2457 24027 2460
rect 23969 2451 24027 2457
rect 20289 2423 20347 2429
rect 20289 2389 20301 2423
rect 20335 2420 20347 2423
rect 22402 2420 22408 2432
rect 20335 2392 22408 2420
rect 20335 2389 20347 2392
rect 20289 2383 20347 2389
rect 22402 2380 22408 2392
rect 22460 2380 22466 2432
rect 22589 2423 22647 2429
rect 22589 2389 22601 2423
rect 22635 2420 22647 2423
rect 23049 2423 23107 2429
rect 23049 2420 23061 2423
rect 22635 2392 23061 2420
rect 22635 2389 22647 2392
rect 22589 2383 22647 2389
rect 23049 2389 23061 2392
rect 23095 2389 23107 2423
rect 23049 2383 23107 2389
rect 17161 2355 17219 2361
rect 17161 2321 17173 2355
rect 17207 2352 17219 2355
rect 18630 2352 18636 2364
rect 17207 2324 18636 2352
rect 17207 2321 17219 2324
rect 17161 2315 17219 2321
rect 18630 2312 18636 2324
rect 18688 2312 18694 2364
rect 20746 2312 20752 2364
rect 20804 2352 20810 2364
rect 20933 2355 20991 2361
rect 20933 2352 20945 2355
rect 20804 2324 20945 2352
rect 20804 2312 20810 2324
rect 20933 2321 20945 2324
rect 20979 2321 20991 2355
rect 20933 2315 20991 2321
rect 21114 2312 21120 2364
rect 21172 2352 21178 2364
rect 21172 2324 21804 2352
rect 21172 2312 21178 2324
rect 13849 2287 13907 2293
rect 13849 2284 13861 2287
rect 13352 2256 13861 2284
rect 13352 2244 13358 2256
rect 13849 2253 13861 2256
rect 13895 2284 13907 2287
rect 14125 2287 14183 2293
rect 14125 2284 14137 2287
rect 13895 2256 14137 2284
rect 13895 2253 13907 2256
rect 13849 2247 13907 2253
rect 14125 2253 14137 2256
rect 14171 2253 14183 2287
rect 14125 2247 14183 2253
rect 14861 2287 14919 2293
rect 14861 2253 14873 2287
rect 14907 2253 14919 2287
rect 14861 2247 14919 2253
rect 15781 2287 15839 2293
rect 15781 2253 15793 2287
rect 15827 2284 15839 2287
rect 16514 2284 16520 2296
rect 15827 2256 16520 2284
rect 15827 2253 15839 2256
rect 15781 2247 15839 2253
rect 15502 2216 15508 2228
rect 11595 2188 12420 2216
rect 13956 2188 15508 2216
rect 11595 2185 11607 2188
rect 11549 2179 11607 2185
rect 10902 2148 10908 2160
rect 9856 2120 10908 2148
rect 9856 2108 9862 2120
rect 10902 2108 10908 2120
rect 10960 2108 10966 2160
rect 13956 2157 13984 2188
rect 15502 2176 15508 2188
rect 15560 2216 15566 2228
rect 15796 2216 15824 2247
rect 16514 2244 16520 2256
rect 16572 2244 16578 2296
rect 17894 2244 17900 2296
rect 17952 2284 17958 2296
rect 17989 2287 18047 2293
rect 17989 2284 18001 2287
rect 17952 2256 18001 2284
rect 17952 2244 17958 2256
rect 17989 2253 18001 2256
rect 18035 2253 18047 2287
rect 17989 2247 18047 2253
rect 19550 2244 19556 2296
rect 19608 2284 19614 2296
rect 19691 2287 19749 2293
rect 19691 2284 19703 2287
rect 19608 2256 19703 2284
rect 19608 2244 19614 2256
rect 19691 2253 19703 2256
rect 19737 2253 19749 2287
rect 19691 2247 19749 2253
rect 20473 2287 20531 2293
rect 20473 2253 20485 2287
rect 20519 2284 20531 2287
rect 21022 2284 21028 2296
rect 20519 2256 21028 2284
rect 20519 2253 20531 2256
rect 20473 2247 20531 2253
rect 21022 2244 21028 2256
rect 21080 2284 21086 2296
rect 21776 2293 21804 2324
rect 21485 2287 21543 2293
rect 21485 2284 21497 2287
rect 21080 2256 21497 2284
rect 21080 2244 21086 2256
rect 21485 2253 21497 2256
rect 21531 2253 21543 2287
rect 21485 2247 21543 2253
rect 21761 2287 21819 2293
rect 21761 2253 21773 2287
rect 21807 2253 21819 2287
rect 21761 2247 21819 2253
rect 21945 2287 22003 2293
rect 21945 2253 21957 2287
rect 21991 2253 22003 2287
rect 21945 2247 22003 2253
rect 22957 2287 23015 2293
rect 22957 2253 22969 2287
rect 23003 2253 23015 2287
rect 22957 2247 23015 2253
rect 15560 2188 15824 2216
rect 16425 2219 16483 2225
rect 15560 2176 15566 2188
rect 16425 2185 16437 2219
rect 16471 2216 16483 2219
rect 16698 2216 16704 2228
rect 16471 2188 16704 2216
rect 16471 2185 16483 2188
rect 16425 2179 16483 2185
rect 16698 2176 16704 2188
rect 16756 2176 16762 2228
rect 17434 2176 17440 2228
rect 17492 2216 17498 2228
rect 18170 2216 18176 2228
rect 17492 2188 18176 2216
rect 17492 2176 17498 2188
rect 18170 2176 18176 2188
rect 18228 2216 18234 2228
rect 18265 2219 18323 2225
rect 18265 2216 18277 2219
rect 18228 2188 18277 2216
rect 18228 2176 18234 2188
rect 18265 2185 18277 2188
rect 18311 2185 18323 2219
rect 18265 2179 18323 2185
rect 13665 2151 13723 2157
rect 13665 2117 13677 2151
rect 13711 2148 13723 2151
rect 13941 2151 13999 2157
rect 13941 2148 13953 2151
rect 13711 2120 13953 2148
rect 13711 2117 13723 2120
rect 13665 2111 13723 2117
rect 13941 2117 13953 2120
rect 13987 2117 13999 2151
rect 18280 2148 18308 2179
rect 19274 2176 19280 2228
rect 19332 2176 19338 2228
rect 20657 2219 20715 2225
rect 20657 2185 20669 2219
rect 20703 2216 20715 2219
rect 21960 2216 21988 2247
rect 22681 2219 22739 2225
rect 22681 2216 22693 2219
rect 20703 2188 22693 2216
rect 20703 2185 20715 2188
rect 20657 2179 20715 2185
rect 22681 2185 22693 2188
rect 22727 2216 22739 2219
rect 22972 2216 23000 2247
rect 22727 2188 23000 2216
rect 23064 2216 23092 2383
rect 24150 2352 24156 2364
rect 24111 2324 24156 2352
rect 24150 2312 24156 2324
rect 24208 2312 24214 2364
rect 24260 2352 24288 2460
rect 24426 2448 24432 2500
rect 24484 2488 24490 2500
rect 25855 2491 25913 2497
rect 25855 2488 25867 2491
rect 24484 2460 25867 2488
rect 24484 2448 24490 2460
rect 25855 2457 25867 2460
rect 25901 2457 25913 2491
rect 25855 2451 25913 2457
rect 24429 2355 24487 2361
rect 24429 2352 24441 2355
rect 24260 2324 24441 2352
rect 24429 2321 24441 2324
rect 24475 2352 24487 2355
rect 26177 2355 26235 2361
rect 26177 2352 26189 2355
rect 24475 2324 26189 2352
rect 24475 2321 24487 2324
rect 24429 2315 24487 2321
rect 26177 2321 26189 2324
rect 26223 2321 26235 2355
rect 26177 2315 26235 2321
rect 23874 2216 23880 2228
rect 23064 2188 23880 2216
rect 22727 2185 22739 2188
rect 22681 2179 22739 2185
rect 20013 2151 20071 2157
rect 20013 2148 20025 2151
rect 18280 2120 20025 2148
rect 13941 2111 13999 2117
rect 20013 2117 20025 2120
rect 20059 2117 20071 2151
rect 20013 2111 20071 2117
rect 20841 2151 20899 2157
rect 20841 2117 20853 2151
rect 20887 2148 20899 2151
rect 20930 2148 20936 2160
rect 20887 2120 20936 2148
rect 20887 2117 20899 2120
rect 20841 2111 20899 2117
rect 20930 2108 20936 2120
rect 20988 2108 20994 2160
rect 22972 2148 23000 2188
rect 23874 2176 23880 2188
rect 23932 2176 23938 2228
rect 24334 2176 24340 2228
rect 24392 2216 24398 2228
rect 24886 2216 24892 2228
rect 24392 2188 24892 2216
rect 24392 2176 24398 2188
rect 24886 2176 24892 2188
rect 24944 2176 24950 2228
rect 23414 2148 23420 2160
rect 22972 2120 23420 2148
rect 23414 2108 23420 2120
rect 23472 2108 23478 2160
rect 23506 2108 23512 2160
rect 23564 2148 23570 2160
rect 23564 2120 23609 2148
rect 23564 2108 23570 2120
rect 400 2058 27264 2080
rect 400 2006 18870 2058
rect 18922 2006 18934 2058
rect 18986 2006 18998 2058
rect 19050 2006 19062 2058
rect 19114 2006 19126 2058
rect 19178 2006 27264 2058
rect 400 1984 27264 2006
rect 7041 1947 7099 1953
rect 7041 1913 7053 1947
rect 7087 1944 7099 1947
rect 7498 1944 7504 1956
rect 7087 1916 7504 1944
rect 7087 1913 7099 1916
rect 7041 1907 7099 1913
rect 7498 1904 7504 1916
rect 7556 1904 7562 1956
rect 10810 1904 10816 1956
rect 10868 1944 10874 1956
rect 11825 1947 11883 1953
rect 11825 1944 11837 1947
rect 10868 1916 11837 1944
rect 10868 1904 10874 1916
rect 11825 1913 11837 1916
rect 11871 1944 11883 1947
rect 12190 1944 12196 1956
rect 11871 1916 12196 1944
rect 11871 1913 11883 1916
rect 11825 1907 11883 1913
rect 12190 1904 12196 1916
rect 12248 1944 12254 1956
rect 13202 1944 13208 1956
rect 12248 1916 13208 1944
rect 12248 1904 12254 1916
rect 13202 1904 13208 1916
rect 13260 1904 13266 1956
rect 17986 1904 17992 1956
rect 18044 1944 18050 1956
rect 18357 1947 18415 1953
rect 18357 1944 18369 1947
rect 18044 1916 18369 1944
rect 18044 1904 18050 1916
rect 18357 1913 18369 1916
rect 18403 1913 18415 1947
rect 18357 1907 18415 1913
rect 18633 1947 18691 1953
rect 18633 1913 18645 1947
rect 18679 1944 18691 1947
rect 19550 1944 19556 1956
rect 18679 1916 19556 1944
rect 18679 1913 18691 1916
rect 18633 1907 18691 1913
rect 4186 1836 4192 1888
rect 4244 1876 4250 1888
rect 4244 1848 4600 1876
rect 4244 1836 4250 1848
rect 1334 1768 1340 1820
rect 1392 1808 1398 1820
rect 1521 1811 1579 1817
rect 1521 1808 1533 1811
rect 1392 1780 1533 1808
rect 1392 1768 1398 1780
rect 1521 1777 1533 1780
rect 1567 1777 1579 1811
rect 1521 1771 1579 1777
rect 2070 1768 2076 1820
rect 2128 1808 2134 1820
rect 2257 1811 2315 1817
rect 2257 1808 2269 1811
rect 2128 1780 2269 1808
rect 2128 1768 2134 1780
rect 2257 1777 2269 1780
rect 2303 1777 2315 1811
rect 2257 1771 2315 1777
rect 2530 1768 2536 1820
rect 2588 1808 2594 1820
rect 3358 1808 3364 1820
rect 2588 1780 3364 1808
rect 2588 1768 2594 1780
rect 3358 1768 3364 1780
rect 3416 1808 3422 1820
rect 4572 1817 4600 1848
rect 6210 1836 6216 1888
rect 6268 1876 6274 1888
rect 6765 1879 6823 1885
rect 6765 1876 6777 1879
rect 6268 1848 6777 1876
rect 6268 1836 6274 1848
rect 6765 1845 6777 1848
rect 6811 1845 6823 1879
rect 7130 1876 7136 1888
rect 7091 1848 7136 1876
rect 6765 1839 6823 1845
rect 3729 1811 3787 1817
rect 3729 1808 3741 1811
rect 3416 1780 3741 1808
rect 3416 1768 3422 1780
rect 3729 1777 3741 1780
rect 3775 1777 3787 1811
rect 3729 1771 3787 1777
rect 4557 1811 4615 1817
rect 4557 1777 4569 1811
rect 4603 1777 4615 1811
rect 5842 1808 5848 1820
rect 5803 1780 5848 1808
rect 4557 1771 4615 1777
rect 5842 1768 5848 1780
rect 5900 1768 5906 1820
rect 6578 1808 6584 1820
rect 6539 1780 6584 1808
rect 6578 1768 6584 1780
rect 6636 1768 6642 1820
rect 6780 1808 6808 1839
rect 7130 1836 7136 1848
rect 7188 1836 7194 1888
rect 8878 1836 8884 1888
rect 8936 1876 8942 1888
rect 9157 1879 9215 1885
rect 9157 1876 9169 1879
rect 8936 1848 9169 1876
rect 8936 1836 8942 1848
rect 9157 1845 9169 1848
rect 9203 1876 9215 1879
rect 9798 1876 9804 1888
rect 9203 1848 9804 1876
rect 9203 1845 9215 1848
rect 9157 1839 9215 1845
rect 9798 1836 9804 1848
rect 9856 1836 9862 1888
rect 11362 1876 11368 1888
rect 11323 1848 11368 1876
rect 11362 1836 11368 1848
rect 11420 1836 11426 1888
rect 15502 1876 15508 1888
rect 15463 1848 15508 1876
rect 15502 1836 15508 1848
rect 15560 1836 15566 1888
rect 15686 1876 15692 1888
rect 15599 1848 15692 1876
rect 15686 1836 15692 1848
rect 15744 1876 15750 1888
rect 16698 1876 16704 1888
rect 15744 1848 16704 1876
rect 15744 1836 15750 1848
rect 16698 1836 16704 1848
rect 16756 1836 16762 1888
rect 18081 1879 18139 1885
rect 18081 1845 18093 1879
rect 18127 1876 18139 1879
rect 18170 1876 18176 1888
rect 18127 1848 18176 1876
rect 18127 1845 18139 1848
rect 18081 1839 18139 1845
rect 18170 1836 18176 1848
rect 18228 1836 18234 1888
rect 18372 1876 18400 1907
rect 19550 1904 19556 1916
rect 19608 1904 19614 1956
rect 20657 1947 20715 1953
rect 20657 1913 20669 1947
rect 20703 1944 20715 1947
rect 20746 1944 20752 1956
rect 20703 1916 20752 1944
rect 20703 1913 20715 1916
rect 20657 1907 20715 1913
rect 20746 1904 20752 1916
rect 20804 1904 20810 1956
rect 22126 1904 22132 1956
rect 22184 1944 22190 1956
rect 23046 1944 23052 1956
rect 22184 1916 23052 1944
rect 22184 1904 22190 1916
rect 23046 1904 23052 1916
rect 23104 1944 23110 1956
rect 23509 1947 23567 1953
rect 23509 1944 23521 1947
rect 23104 1916 23521 1944
rect 23104 1904 23110 1916
rect 23509 1913 23521 1916
rect 23555 1913 23567 1947
rect 23509 1907 23567 1913
rect 23874 1904 23880 1956
rect 23932 1944 23938 1956
rect 23932 1916 23977 1944
rect 23932 1904 23938 1916
rect 24058 1904 24064 1956
rect 24116 1944 24122 1956
rect 24245 1947 24303 1953
rect 24245 1944 24257 1947
rect 24116 1916 24257 1944
rect 24116 1904 24122 1916
rect 24245 1913 24257 1916
rect 24291 1913 24303 1947
rect 24245 1907 24303 1913
rect 24334 1904 24340 1956
rect 24392 1944 24398 1956
rect 24429 1947 24487 1953
rect 24429 1944 24441 1947
rect 24392 1916 24441 1944
rect 24392 1904 24398 1916
rect 24429 1913 24441 1916
rect 24475 1913 24487 1947
rect 24429 1907 24487 1913
rect 24702 1904 24708 1956
rect 24760 1944 24766 1956
rect 25901 1947 25959 1953
rect 25901 1944 25913 1947
rect 24760 1916 25913 1944
rect 24760 1904 24766 1916
rect 25901 1913 25913 1916
rect 25947 1944 25959 1947
rect 26358 1944 26364 1956
rect 25947 1916 26364 1944
rect 25947 1913 25959 1916
rect 25901 1907 25959 1913
rect 26358 1904 26364 1916
rect 26416 1904 26422 1956
rect 19277 1879 19335 1885
rect 19277 1876 19289 1879
rect 18372 1848 19289 1876
rect 19277 1845 19289 1848
rect 19323 1876 19335 1879
rect 19458 1876 19464 1888
rect 19323 1848 19464 1876
rect 19323 1845 19335 1848
rect 19277 1839 19335 1845
rect 19458 1836 19464 1848
rect 19516 1836 19522 1888
rect 23230 1876 23236 1888
rect 23143 1848 23236 1876
rect 23230 1836 23236 1848
rect 23288 1876 23294 1888
rect 23598 1876 23604 1888
rect 23288 1848 23604 1876
rect 23288 1836 23294 1848
rect 23598 1836 23604 1848
rect 23656 1836 23662 1888
rect 24150 1876 24156 1888
rect 24111 1848 24156 1876
rect 24150 1836 24156 1848
rect 24208 1836 24214 1888
rect 7774 1808 7780 1820
rect 6780 1780 7780 1808
rect 7774 1768 7780 1780
rect 7832 1768 7838 1820
rect 8142 1768 8148 1820
rect 8200 1808 8206 1820
rect 9065 1811 9123 1817
rect 9065 1808 9077 1811
rect 8200 1780 9077 1808
rect 8200 1768 8206 1780
rect 9065 1777 9077 1780
rect 9111 1808 9123 1811
rect 9706 1808 9712 1820
rect 9111 1780 9712 1808
rect 9111 1777 9123 1780
rect 9065 1771 9123 1777
rect 9706 1768 9712 1780
rect 9764 1768 9770 1820
rect 9890 1808 9896 1820
rect 9803 1780 9896 1808
rect 9890 1768 9896 1780
rect 9948 1808 9954 1820
rect 10166 1808 10172 1820
rect 9948 1780 10172 1808
rect 9948 1768 9954 1780
rect 10166 1768 10172 1780
rect 10224 1768 10230 1820
rect 12282 1768 12288 1820
rect 12340 1808 12346 1820
rect 12561 1811 12619 1817
rect 12561 1808 12573 1811
rect 12340 1780 12573 1808
rect 12340 1768 12346 1780
rect 12561 1777 12573 1780
rect 12607 1777 12619 1811
rect 13386 1808 13392 1820
rect 13347 1780 13392 1808
rect 12561 1771 12619 1777
rect 13386 1768 13392 1780
rect 13444 1768 13450 1820
rect 14582 1808 14588 1820
rect 14543 1780 14588 1808
rect 14582 1768 14588 1780
rect 14640 1768 14646 1820
rect 15226 1808 15232 1820
rect 15187 1780 15232 1808
rect 15226 1768 15232 1780
rect 15284 1768 15290 1820
rect 16514 1808 16520 1820
rect 16475 1780 16520 1808
rect 16514 1768 16520 1780
rect 16572 1768 16578 1820
rect 18725 1811 18783 1817
rect 18725 1777 18737 1811
rect 18771 1777 18783 1811
rect 18906 1808 18912 1820
rect 18867 1780 18912 1808
rect 18725 1771 18783 1777
rect 1242 1700 1248 1752
rect 1300 1740 1306 1752
rect 1429 1743 1487 1749
rect 1429 1740 1441 1743
rect 1300 1712 1441 1740
rect 1300 1700 1306 1712
rect 1429 1709 1441 1712
rect 1475 1740 1487 1743
rect 2162 1740 2168 1752
rect 1475 1712 2168 1740
rect 1475 1709 1487 1712
rect 1429 1703 1487 1709
rect 2162 1700 2168 1712
rect 2220 1700 2226 1752
rect 2346 1740 2352 1752
rect 2307 1712 2352 1740
rect 2346 1700 2352 1712
rect 2404 1700 2410 1752
rect 3821 1743 3879 1749
rect 3821 1709 3833 1743
rect 3867 1740 3879 1743
rect 3910 1740 3916 1752
rect 3867 1712 3916 1740
rect 3867 1709 3879 1712
rect 3821 1703 3879 1709
rect 3910 1700 3916 1712
rect 3968 1700 3974 1752
rect 4278 1700 4284 1752
rect 4336 1740 4342 1752
rect 4649 1743 4707 1749
rect 4649 1740 4661 1743
rect 4336 1712 4661 1740
rect 4336 1700 4342 1712
rect 4649 1709 4661 1712
rect 4695 1709 4707 1743
rect 9982 1740 9988 1752
rect 9943 1712 9988 1740
rect 4649 1703 4707 1709
rect 9982 1700 9988 1712
rect 10040 1700 10046 1752
rect 10902 1740 10908 1752
rect 10863 1712 10908 1740
rect 10902 1700 10908 1712
rect 10960 1700 10966 1752
rect 11454 1740 11460 1752
rect 11415 1712 11460 1740
rect 11454 1700 11460 1712
rect 11512 1700 11518 1752
rect 12653 1743 12711 1749
rect 12653 1709 12665 1743
rect 12699 1740 12711 1743
rect 13018 1740 13024 1752
rect 12699 1712 13024 1740
rect 12699 1709 12711 1712
rect 12653 1703 12711 1709
rect 13018 1700 13024 1712
rect 13076 1700 13082 1752
rect 13478 1740 13484 1752
rect 13439 1712 13484 1740
rect 13478 1700 13484 1712
rect 13536 1740 13542 1752
rect 14398 1740 14404 1752
rect 13536 1712 14404 1740
rect 13536 1700 13542 1712
rect 14398 1700 14404 1712
rect 14456 1700 14462 1752
rect 18078 1700 18084 1752
rect 18136 1740 18142 1752
rect 18173 1743 18231 1749
rect 18173 1740 18185 1743
rect 18136 1712 18185 1740
rect 18136 1700 18142 1712
rect 18173 1709 18185 1712
rect 18219 1709 18231 1743
rect 18740 1740 18768 1771
rect 18906 1768 18912 1780
rect 18964 1768 18970 1820
rect 20838 1808 20844 1820
rect 20799 1780 20844 1808
rect 20838 1768 20844 1780
rect 20896 1768 20902 1820
rect 23414 1808 23420 1820
rect 23375 1780 23420 1808
rect 23414 1768 23420 1780
rect 23472 1768 23478 1820
rect 26085 1811 26143 1817
rect 26085 1777 26097 1811
rect 26131 1808 26143 1811
rect 26266 1808 26272 1820
rect 26131 1780 26272 1808
rect 26131 1777 26143 1780
rect 26085 1771 26143 1777
rect 26266 1768 26272 1780
rect 26324 1768 26330 1820
rect 18998 1740 19004 1752
rect 18740 1712 19004 1740
rect 18173 1703 18231 1709
rect 18998 1700 19004 1712
rect 19056 1740 19062 1752
rect 20470 1740 20476 1752
rect 19056 1712 20476 1740
rect 19056 1700 19062 1712
rect 20470 1700 20476 1712
rect 20528 1700 20534 1752
rect 21758 1740 21764 1752
rect 21719 1712 21764 1740
rect 21758 1700 21764 1712
rect 21816 1700 21822 1752
rect 7590 1604 7596 1616
rect 7551 1576 7596 1604
rect 7590 1564 7596 1576
rect 7648 1564 7654 1616
rect 11822 1564 11828 1616
rect 11880 1604 11886 1616
rect 15686 1604 15692 1616
rect 11880 1576 15692 1604
rect 11880 1564 11886 1576
rect 15686 1564 15692 1576
rect 15744 1564 15750 1616
rect 16330 1604 16336 1616
rect 16291 1576 16336 1604
rect 16330 1564 16336 1576
rect 16388 1564 16394 1616
rect 17894 1604 17900 1616
rect 17855 1576 17900 1604
rect 17894 1564 17900 1576
rect 17952 1564 17958 1616
rect 400 1514 27264 1536
rect 400 1462 3510 1514
rect 3562 1462 3574 1514
rect 3626 1462 3638 1514
rect 3690 1462 3702 1514
rect 3754 1462 3766 1514
rect 3818 1462 27264 1514
rect 400 1440 27264 1462
rect 1242 1400 1248 1412
rect 1203 1372 1248 1400
rect 1242 1360 1248 1372
rect 1300 1360 1306 1412
rect 2070 1400 2076 1412
rect 2031 1372 2076 1400
rect 2070 1360 2076 1372
rect 2128 1360 2134 1412
rect 2257 1403 2315 1409
rect 2257 1369 2269 1403
rect 2303 1400 2315 1403
rect 2346 1400 2352 1412
rect 2303 1372 2352 1400
rect 2303 1369 2315 1372
rect 2257 1363 2315 1369
rect 2346 1360 2352 1372
rect 2404 1360 2410 1412
rect 3085 1403 3143 1409
rect 3085 1369 3097 1403
rect 3131 1400 3143 1403
rect 3266 1400 3272 1412
rect 3131 1372 3272 1400
rect 3131 1369 3143 1372
rect 3085 1363 3143 1369
rect 3266 1360 3272 1372
rect 3324 1400 3330 1412
rect 3453 1403 3511 1409
rect 3453 1400 3465 1403
rect 3324 1372 3465 1400
rect 3324 1360 3330 1372
rect 3453 1369 3465 1372
rect 3499 1369 3511 1403
rect 7041 1403 7099 1409
rect 7041 1400 7053 1403
rect 3453 1363 3511 1369
rect 6688 1372 7053 1400
rect 2088 1332 2116 1360
rect 4186 1332 4192 1344
rect 2088 1304 4192 1332
rect 4186 1292 4192 1304
rect 4244 1292 4250 1344
rect 414 1224 420 1276
rect 472 1264 478 1276
rect 6688 1273 6716 1372
rect 7041 1369 7053 1372
rect 7087 1400 7099 1403
rect 7590 1400 7596 1412
rect 7087 1372 7596 1400
rect 7087 1369 7099 1372
rect 7041 1363 7099 1369
rect 7590 1360 7596 1372
rect 7648 1400 7654 1412
rect 7777 1403 7835 1409
rect 7777 1400 7789 1403
rect 7648 1372 7789 1400
rect 7648 1360 7654 1372
rect 7777 1369 7789 1372
rect 7823 1369 7835 1403
rect 7777 1363 7835 1369
rect 7866 1360 7872 1412
rect 7924 1400 7930 1412
rect 8329 1403 8387 1409
rect 8329 1400 8341 1403
rect 7924 1372 8341 1400
rect 7924 1360 7930 1372
rect 8329 1369 8341 1372
rect 8375 1369 8387 1403
rect 8878 1400 8884 1412
rect 8839 1372 8884 1400
rect 8329 1363 8387 1369
rect 8344 1332 8372 1363
rect 8878 1360 8884 1372
rect 8936 1360 8942 1412
rect 9706 1400 9712 1412
rect 9667 1372 9712 1400
rect 9706 1360 9712 1372
rect 9764 1360 9770 1412
rect 10077 1403 10135 1409
rect 10077 1400 10089 1403
rect 9816 1372 10089 1400
rect 9617 1335 9675 1341
rect 9617 1332 9629 1335
rect 8344 1304 9629 1332
rect 9617 1301 9629 1304
rect 9663 1332 9675 1335
rect 9816 1332 9844 1372
rect 10077 1369 10089 1372
rect 10123 1369 10135 1403
rect 10902 1400 10908 1412
rect 10863 1372 10908 1400
rect 10077 1363 10135 1369
rect 10902 1360 10908 1372
rect 10960 1360 10966 1412
rect 11181 1403 11239 1409
rect 11181 1369 11193 1403
rect 11227 1400 11239 1403
rect 11454 1400 11460 1412
rect 11227 1372 11460 1400
rect 11227 1369 11239 1372
rect 11181 1363 11239 1369
rect 11454 1360 11460 1372
rect 11512 1400 11518 1412
rect 11733 1403 11791 1409
rect 11733 1400 11745 1403
rect 11512 1372 11745 1400
rect 11512 1360 11518 1372
rect 11733 1369 11745 1372
rect 11779 1400 11791 1403
rect 12009 1403 12067 1409
rect 12009 1400 12021 1403
rect 11779 1372 12021 1400
rect 11779 1369 11791 1372
rect 11733 1363 11791 1369
rect 12009 1369 12021 1372
rect 12055 1369 12067 1403
rect 12190 1400 12196 1412
rect 12151 1372 12196 1400
rect 12009 1363 12067 1369
rect 12190 1360 12196 1372
rect 12248 1360 12254 1412
rect 12745 1403 12803 1409
rect 12745 1369 12757 1403
rect 12791 1400 12803 1403
rect 13478 1400 13484 1412
rect 12791 1372 13484 1400
rect 12791 1369 12803 1372
rect 12745 1363 12803 1369
rect 13478 1360 13484 1372
rect 13536 1360 13542 1412
rect 16330 1400 16336 1412
rect 15060 1372 16336 1400
rect 9663 1304 9844 1332
rect 9985 1335 10043 1341
rect 9663 1301 9675 1304
rect 9617 1295 9675 1301
rect 9985 1301 9997 1335
rect 10031 1332 10043 1335
rect 11822 1332 11828 1344
rect 10031 1304 11828 1332
rect 10031 1301 10043 1304
rect 9985 1295 10043 1301
rect 4005 1267 4063 1273
rect 4005 1264 4017 1267
rect 472 1236 4017 1264
rect 472 1224 478 1236
rect 1061 1199 1119 1205
rect 1061 1165 1073 1199
rect 1107 1196 1119 1199
rect 1334 1196 1340 1208
rect 1107 1168 1340 1196
rect 1107 1165 1119 1168
rect 1061 1159 1119 1165
rect 1334 1156 1340 1168
rect 1392 1156 1398 1208
rect 3376 1205 3404 1236
rect 4005 1233 4017 1236
rect 4051 1233 4063 1267
rect 4005 1227 4063 1233
rect 6673 1267 6731 1273
rect 6673 1233 6685 1267
rect 6719 1233 6731 1267
rect 6673 1227 6731 1233
rect 7498 1224 7504 1276
rect 7556 1264 7562 1276
rect 7593 1267 7651 1273
rect 7593 1264 7605 1267
rect 7556 1236 7605 1264
rect 7556 1224 7562 1236
rect 7593 1233 7605 1236
rect 7639 1264 7651 1267
rect 8145 1267 8203 1273
rect 8145 1264 8157 1267
rect 7639 1236 8157 1264
rect 7639 1233 7651 1236
rect 7593 1227 7651 1233
rect 8145 1233 8157 1236
rect 8191 1233 8203 1267
rect 8145 1227 8203 1233
rect 8326 1224 8332 1276
rect 8384 1264 8390 1276
rect 9065 1267 9123 1273
rect 9065 1264 9077 1267
rect 8384 1236 9077 1264
rect 8384 1224 8390 1236
rect 9065 1233 9077 1236
rect 9111 1264 9123 1267
rect 9890 1264 9896 1276
rect 9111 1236 9896 1264
rect 9111 1233 9123 1236
rect 9065 1227 9123 1233
rect 9890 1224 9896 1236
rect 9948 1224 9954 1276
rect 3361 1199 3419 1205
rect 3361 1165 3373 1199
rect 3407 1165 3419 1199
rect 3361 1159 3419 1165
rect 3910 1156 3916 1208
rect 3968 1196 3974 1208
rect 5842 1196 5848 1208
rect 3968 1168 5848 1196
rect 3968 1156 3974 1168
rect 5842 1156 5848 1168
rect 5900 1196 5906 1208
rect 6121 1199 6179 1205
rect 6121 1196 6133 1199
rect 5900 1168 6133 1196
rect 5900 1156 5906 1168
rect 6121 1165 6133 1168
rect 6167 1196 6179 1199
rect 6765 1199 6823 1205
rect 6765 1196 6777 1199
rect 6167 1168 6777 1196
rect 6167 1165 6179 1168
rect 6121 1159 6179 1165
rect 6765 1165 6777 1168
rect 6811 1165 6823 1199
rect 6765 1159 6823 1165
rect 9249 1199 9307 1205
rect 9249 1165 9261 1199
rect 9295 1196 9307 1199
rect 9982 1196 9988 1208
rect 9295 1168 9988 1196
rect 9295 1165 9307 1168
rect 9249 1159 9307 1165
rect 9982 1156 9988 1168
rect 10040 1156 10046 1208
rect 877 1131 935 1137
rect 877 1097 889 1131
rect 923 1128 935 1131
rect 923 1100 1380 1128
rect 923 1097 935 1100
rect 877 1091 935 1097
rect 1352 1060 1380 1100
rect 1610 1088 1616 1140
rect 1668 1128 1674 1140
rect 1797 1131 1855 1137
rect 1797 1128 1809 1131
rect 1668 1100 1809 1128
rect 1668 1088 1674 1100
rect 1797 1097 1809 1100
rect 1843 1097 1855 1131
rect 1797 1091 1855 1097
rect 1889 1131 1947 1137
rect 1889 1097 1901 1131
rect 1935 1128 1947 1131
rect 3082 1128 3088 1140
rect 1935 1100 3088 1128
rect 1935 1097 1947 1100
rect 1889 1091 1947 1097
rect 1904 1060 1932 1091
rect 3082 1088 3088 1100
rect 3140 1088 3146 1140
rect 3177 1131 3235 1137
rect 3177 1097 3189 1131
rect 3223 1128 3235 1131
rect 5569 1131 5627 1137
rect 3223 1100 3956 1128
rect 3223 1097 3235 1100
rect 3177 1091 3235 1097
rect 3928 1072 3956 1100
rect 5569 1097 5581 1131
rect 5615 1128 5627 1131
rect 5753 1131 5811 1137
rect 5753 1128 5765 1131
rect 5615 1100 5765 1128
rect 5615 1097 5627 1100
rect 5569 1091 5627 1097
rect 5753 1097 5765 1100
rect 5799 1128 5811 1131
rect 6578 1128 6584 1140
rect 5799 1100 6584 1128
rect 5799 1097 5811 1100
rect 5753 1091 5811 1097
rect 6578 1088 6584 1100
rect 6636 1128 6642 1140
rect 7501 1131 7559 1137
rect 7501 1128 7513 1131
rect 6636 1100 7513 1128
rect 6636 1088 6642 1100
rect 7501 1097 7513 1100
rect 7547 1128 7559 1131
rect 7961 1131 8019 1137
rect 7961 1128 7973 1131
rect 7547 1100 7973 1128
rect 7547 1097 7559 1100
rect 7501 1091 7559 1097
rect 7961 1097 7973 1100
rect 8007 1097 8019 1131
rect 7961 1091 8019 1097
rect 9433 1131 9491 1137
rect 9433 1097 9445 1131
rect 9479 1128 9491 1131
rect 10092 1128 10120 1304
rect 11822 1292 11828 1304
rect 11880 1292 11886 1344
rect 12282 1292 12288 1344
rect 12340 1332 12346 1344
rect 12837 1335 12895 1341
rect 12837 1332 12849 1335
rect 12340 1304 12849 1332
rect 12340 1292 12346 1304
rect 12837 1301 12849 1304
rect 12883 1301 12895 1335
rect 13018 1332 13024 1344
rect 12979 1304 13024 1332
rect 12837 1295 12895 1301
rect 13018 1292 13024 1304
rect 13076 1332 13082 1344
rect 13076 1304 14214 1332
rect 13076 1292 13082 1304
rect 11362 1264 11368 1276
rect 11323 1236 11368 1264
rect 11362 1224 11368 1236
rect 11420 1224 11426 1276
rect 11917 1199 11975 1205
rect 11917 1165 11929 1199
rect 11963 1196 11975 1199
rect 12190 1196 12196 1208
rect 11963 1168 12196 1196
rect 11963 1165 11975 1168
rect 11917 1159 11975 1165
rect 12190 1156 12196 1168
rect 12248 1156 12254 1208
rect 14186 1196 14214 1304
rect 15060 1273 15088 1372
rect 16330 1360 16336 1372
rect 16388 1360 16394 1412
rect 16606 1360 16612 1412
rect 16664 1400 16670 1412
rect 16701 1403 16759 1409
rect 16701 1400 16713 1403
rect 16664 1372 16713 1400
rect 16664 1360 16670 1372
rect 16701 1369 16713 1372
rect 16747 1369 16759 1403
rect 18998 1400 19004 1412
rect 18959 1372 19004 1400
rect 16701 1363 16759 1369
rect 18998 1360 19004 1372
rect 19056 1360 19062 1412
rect 19277 1403 19335 1409
rect 19277 1369 19289 1403
rect 19323 1400 19335 1403
rect 19737 1403 19795 1409
rect 19737 1400 19749 1403
rect 19323 1372 19749 1400
rect 19323 1369 19335 1372
rect 19277 1363 19335 1369
rect 19737 1369 19749 1372
rect 19783 1400 19795 1403
rect 20565 1403 20623 1409
rect 20565 1400 20577 1403
rect 19783 1372 20577 1400
rect 19783 1369 19795 1372
rect 19737 1363 19795 1369
rect 20565 1369 20577 1372
rect 20611 1400 20623 1403
rect 20838 1400 20844 1412
rect 20611 1372 20844 1400
rect 20611 1369 20623 1372
rect 20565 1363 20623 1369
rect 20838 1360 20844 1372
rect 20896 1360 20902 1412
rect 20933 1403 20991 1409
rect 20933 1369 20945 1403
rect 20979 1400 20991 1403
rect 21022 1400 21028 1412
rect 20979 1372 21028 1400
rect 20979 1369 20991 1372
rect 20933 1363 20991 1369
rect 21022 1360 21028 1372
rect 21080 1400 21086 1412
rect 21485 1403 21543 1409
rect 21485 1400 21497 1403
rect 21080 1372 21497 1400
rect 21080 1360 21086 1372
rect 21485 1369 21497 1372
rect 21531 1369 21543 1403
rect 23046 1400 23052 1412
rect 23007 1372 23052 1400
rect 21485 1363 21543 1369
rect 23046 1360 23052 1372
rect 23104 1360 23110 1412
rect 23230 1400 23236 1412
rect 23191 1372 23236 1400
rect 23230 1360 23236 1372
rect 23288 1360 23294 1412
rect 23414 1400 23420 1412
rect 23375 1372 23420 1400
rect 23414 1360 23420 1372
rect 23472 1360 23478 1412
rect 23785 1403 23843 1409
rect 23785 1369 23797 1403
rect 23831 1400 23843 1403
rect 24150 1400 24156 1412
rect 23831 1372 24156 1400
rect 23831 1369 23843 1372
rect 23785 1363 23843 1369
rect 24150 1360 24156 1372
rect 24208 1360 24214 1412
rect 26358 1400 26364 1412
rect 26319 1372 26364 1400
rect 26358 1360 26364 1372
rect 26416 1360 26422 1412
rect 15962 1332 15968 1344
rect 15923 1304 15968 1332
rect 15962 1292 15968 1304
rect 16020 1332 16026 1344
rect 16517 1335 16575 1341
rect 16517 1332 16529 1335
rect 16020 1304 16529 1332
rect 16020 1292 16026 1304
rect 16517 1301 16529 1304
rect 16563 1301 16575 1335
rect 19458 1332 19464 1344
rect 19419 1304 19464 1332
rect 16517 1295 16575 1301
rect 19458 1292 19464 1304
rect 19516 1292 19522 1344
rect 21209 1335 21267 1341
rect 21209 1301 21221 1335
rect 21255 1332 21267 1335
rect 21758 1332 21764 1344
rect 21255 1304 21764 1332
rect 21255 1301 21267 1304
rect 21209 1295 21267 1301
rect 21758 1292 21764 1304
rect 21816 1332 21822 1344
rect 21816 1304 23874 1332
rect 21816 1292 21822 1304
rect 14401 1267 14459 1273
rect 14401 1233 14413 1267
rect 14447 1264 14459 1267
rect 15045 1267 15103 1273
rect 15045 1264 15057 1267
rect 14447 1236 15057 1264
rect 14447 1233 14459 1236
rect 14401 1227 14459 1233
rect 15045 1233 15057 1236
rect 15091 1233 15103 1267
rect 15045 1227 15103 1233
rect 15229 1267 15287 1273
rect 15229 1233 15241 1267
rect 15275 1264 15287 1267
rect 15321 1267 15379 1273
rect 15321 1264 15333 1267
rect 15275 1236 15333 1264
rect 15275 1233 15287 1236
rect 15229 1227 15287 1233
rect 15321 1233 15333 1236
rect 15367 1233 15379 1267
rect 15321 1227 15379 1233
rect 14493 1199 14551 1205
rect 14493 1196 14505 1199
rect 14186 1168 14505 1196
rect 14493 1165 14505 1168
rect 14539 1196 14551 1199
rect 14582 1196 14588 1208
rect 14539 1168 14588 1196
rect 14539 1165 14551 1168
rect 14493 1159 14551 1165
rect 14582 1156 14588 1168
rect 14640 1196 14646 1208
rect 15244 1196 15272 1227
rect 18446 1224 18452 1276
rect 18504 1264 18510 1276
rect 20930 1264 20936 1276
rect 18504 1236 20936 1264
rect 18504 1224 18510 1236
rect 14640 1168 15272 1196
rect 15873 1199 15931 1205
rect 14640 1156 14646 1168
rect 15873 1165 15885 1199
rect 15919 1196 15931 1199
rect 16149 1199 16207 1205
rect 16149 1196 16161 1199
rect 15919 1168 16161 1196
rect 15919 1165 15931 1168
rect 15873 1159 15931 1165
rect 16149 1165 16161 1168
rect 16195 1165 16207 1199
rect 16149 1159 16207 1165
rect 9479 1100 10120 1128
rect 14033 1131 14091 1137
rect 9479 1097 9491 1100
rect 9433 1091 9491 1097
rect 14033 1097 14045 1131
rect 14079 1128 14091 1131
rect 14217 1131 14275 1137
rect 14217 1128 14229 1131
rect 14079 1100 14229 1128
rect 14079 1097 14091 1100
rect 14033 1091 14091 1097
rect 14217 1097 14229 1100
rect 14263 1128 14275 1131
rect 14953 1131 15011 1137
rect 14953 1128 14965 1131
rect 14263 1100 14965 1128
rect 14263 1097 14275 1100
rect 14217 1091 14275 1097
rect 14953 1097 14965 1100
rect 14999 1128 15011 1131
rect 15226 1128 15232 1140
rect 14999 1100 15232 1128
rect 14999 1097 15011 1100
rect 14953 1091 15011 1097
rect 15226 1088 15232 1100
rect 15284 1128 15290 1140
rect 15888 1128 15916 1159
rect 16422 1156 16428 1208
rect 16480 1196 16486 1208
rect 20672 1205 20700 1236
rect 20930 1224 20936 1236
rect 20988 1264 20994 1276
rect 21301 1267 21359 1273
rect 21301 1264 21313 1267
rect 20988 1236 21313 1264
rect 20988 1224 20994 1236
rect 21301 1233 21313 1236
rect 21347 1233 21359 1267
rect 21301 1227 21359 1233
rect 17897 1199 17955 1205
rect 17897 1196 17909 1199
rect 16480 1168 17909 1196
rect 16480 1156 16486 1168
rect 17897 1165 17909 1168
rect 17943 1196 17955 1199
rect 18357 1199 18415 1205
rect 18357 1196 18369 1199
rect 17943 1168 18369 1196
rect 17943 1165 17955 1168
rect 17897 1159 17955 1165
rect 18357 1165 18369 1168
rect 18403 1165 18415 1199
rect 19277 1199 19335 1205
rect 19277 1196 19289 1199
rect 18357 1159 18415 1165
rect 18464 1168 19289 1196
rect 15284 1100 15916 1128
rect 15284 1088 15290 1100
rect 16698 1088 16704 1140
rect 16756 1128 16762 1140
rect 18464 1128 18492 1168
rect 19277 1165 19289 1168
rect 19323 1196 19335 1199
rect 19829 1199 19887 1205
rect 19829 1196 19841 1199
rect 19323 1168 19841 1196
rect 19323 1165 19335 1168
rect 19277 1159 19335 1165
rect 19829 1165 19841 1168
rect 19875 1165 19887 1199
rect 19829 1159 19887 1165
rect 20657 1199 20715 1205
rect 20657 1165 20669 1199
rect 20703 1165 20715 1199
rect 23846 1196 23874 1304
rect 24168 1264 24196 1360
rect 24337 1267 24395 1273
rect 24337 1264 24349 1267
rect 24168 1236 24349 1264
rect 24337 1233 24349 1236
rect 24383 1264 24395 1267
rect 26085 1267 26143 1273
rect 26085 1264 26097 1267
rect 24383 1236 26097 1264
rect 24383 1233 24395 1236
rect 24337 1227 24395 1233
rect 26085 1233 26097 1236
rect 26131 1233 26143 1267
rect 26085 1227 26143 1233
rect 24061 1199 24119 1205
rect 24061 1196 24073 1199
rect 23846 1168 24073 1196
rect 20657 1159 20715 1165
rect 24061 1165 24073 1168
rect 24107 1165 24119 1199
rect 24061 1159 24119 1165
rect 16756 1100 18492 1128
rect 18817 1131 18875 1137
rect 16756 1088 16762 1100
rect 18817 1097 18829 1131
rect 18863 1128 18875 1131
rect 18906 1128 18912 1140
rect 18863 1100 18912 1128
rect 18863 1097 18875 1100
rect 18817 1091 18875 1097
rect 18906 1088 18912 1100
rect 18964 1128 18970 1140
rect 20470 1128 20476 1140
rect 18964 1100 20476 1128
rect 18964 1088 18970 1100
rect 20470 1088 20476 1100
rect 20528 1088 20534 1140
rect 3910 1060 3916 1072
rect 1352 1032 1932 1060
rect 3871 1032 3916 1060
rect 3910 1020 3916 1032
rect 3968 1020 3974 1072
rect 4278 1020 4284 1072
rect 4336 1060 4342 1072
rect 4373 1063 4431 1069
rect 4373 1060 4385 1063
rect 4336 1032 4385 1060
rect 4336 1020 4342 1032
rect 4373 1029 4385 1032
rect 4419 1029 4431 1063
rect 4373 1023 4431 1029
rect 9890 1020 9896 1072
rect 9948 1060 9954 1072
rect 12469 1063 12527 1069
rect 12469 1060 12481 1063
rect 9948 1032 12481 1060
rect 9948 1020 9954 1032
rect 12469 1029 12481 1032
rect 12515 1060 12527 1063
rect 13386 1060 13392 1072
rect 12515 1032 13392 1060
rect 12515 1029 12527 1032
rect 12469 1023 12527 1029
rect 13386 1020 13392 1032
rect 13444 1020 13450 1072
rect 17894 1020 17900 1072
rect 17952 1060 17958 1072
rect 18173 1063 18231 1069
rect 18173 1060 18185 1063
rect 17952 1032 18185 1060
rect 17952 1020 17958 1032
rect 18173 1029 18185 1032
rect 18219 1060 18231 1063
rect 18630 1060 18636 1072
rect 18219 1032 18636 1060
rect 18219 1029 18231 1032
rect 18173 1023 18231 1029
rect 18630 1020 18636 1032
rect 18688 1020 18694 1072
rect 23969 1063 24027 1069
rect 23969 1029 23981 1063
rect 24015 1060 24027 1063
rect 24076 1060 24104 1159
rect 25622 1156 25628 1208
rect 25680 1196 25686 1208
rect 25763 1199 25821 1205
rect 25763 1196 25775 1199
rect 25680 1168 25775 1196
rect 25680 1156 25686 1168
rect 25763 1165 25775 1168
rect 25809 1165 25821 1199
rect 25763 1159 25821 1165
rect 24886 1088 24892 1140
rect 24944 1088 24950 1140
rect 24518 1060 24524 1072
rect 24015 1032 24524 1060
rect 24015 1029 24027 1032
rect 23969 1023 24027 1029
rect 24518 1020 24524 1032
rect 24576 1020 24582 1072
rect 26266 1060 26272 1072
rect 26227 1032 26272 1060
rect 26266 1020 26272 1032
rect 26324 1020 26330 1072
rect 400 970 27264 992
rect 400 918 18870 970
rect 18922 918 18934 970
rect 18986 918 18998 970
rect 19050 918 19062 970
rect 19114 918 19126 970
rect 19178 918 27264 970
rect 400 896 27264 918
rect 1334 856 1340 868
rect 1295 828 1340 856
rect 1334 816 1340 828
rect 1392 816 1398 868
rect 1610 856 1616 868
rect 1571 828 1616 856
rect 1610 816 1616 828
rect 1668 816 1674 868
rect 3358 816 3364 868
rect 3416 856 3422 868
rect 3637 859 3695 865
rect 3637 856 3649 859
rect 3416 828 3649 856
rect 3416 816 3422 828
rect 3637 825 3649 828
rect 3683 825 3695 859
rect 3818 856 3824 868
rect 3779 828 3824 856
rect 3637 819 3695 825
rect 3818 816 3824 828
rect 3876 816 3882 868
rect 3910 816 3916 868
rect 3968 856 3974 868
rect 5937 859 5995 865
rect 3968 828 4554 856
rect 3968 816 3974 828
rect 4526 788 4554 828
rect 5937 825 5949 859
rect 5983 856 5995 859
rect 6210 856 6216 868
rect 5983 828 6216 856
rect 5983 825 5995 828
rect 5937 819 5995 825
rect 6210 816 6216 828
rect 6268 816 6274 868
rect 14861 859 14919 865
rect 14861 825 14873 859
rect 14907 856 14919 859
rect 15502 856 15508 868
rect 14907 828 15508 856
rect 14907 825 14919 828
rect 14861 819 14919 825
rect 15502 816 15508 828
rect 15560 816 15566 868
rect 24153 859 24211 865
rect 24153 825 24165 859
rect 24199 856 24211 859
rect 25622 856 25628 868
rect 24199 828 25628 856
rect 24199 825 24211 828
rect 24153 819 24211 825
rect 25622 816 25628 828
rect 25680 816 25686 868
rect 16422 788 16428 800
rect 4526 760 16428 788
rect 16422 748 16428 760
rect 16480 748 16486 800
rect 24337 791 24395 797
rect 24337 757 24349 791
rect 24383 788 24395 791
rect 24886 788 24892 800
rect 24383 760 24892 788
rect 24383 757 24395 760
rect 24337 751 24395 757
rect 24886 748 24892 760
rect 24944 748 24950 800
rect 11638 544 11644 596
rect 11696 584 11702 596
rect 12374 584 12380 596
rect 11696 556 12380 584
rect 11696 544 11702 556
rect 12374 544 12380 556
rect 12432 544 12438 596
rect 400 426 27264 448
rect 400 374 3510 426
rect 3562 374 3574 426
rect 3626 374 3638 426
rect 3690 374 3702 426
rect 3754 374 3766 426
rect 3818 374 27264 426
rect 400 352 27264 374
<< via1 >>
rect 25444 27268 25496 27320
rect 26364 27268 26416 27320
rect 18870 27030 18922 27082
rect 18934 27030 18986 27082
rect 18998 27030 19050 27082
rect 19062 27030 19114 27082
rect 19126 27030 19178 27082
rect 6216 26767 6268 26776
rect 6216 26733 6225 26767
rect 6225 26733 6259 26767
rect 6259 26733 6268 26767
rect 6216 26724 6268 26733
rect 6492 26724 6544 26776
rect 6676 26699 6728 26708
rect 6676 26665 6685 26699
rect 6685 26665 6719 26699
rect 6719 26665 6728 26699
rect 6676 26656 6728 26665
rect 7688 26588 7740 26640
rect 24064 26588 24116 26640
rect 3510 26486 3562 26538
rect 3574 26486 3626 26538
rect 3638 26486 3690 26538
rect 3702 26486 3754 26538
rect 3766 26486 3818 26538
rect 6676 26427 6728 26436
rect 6676 26393 6685 26427
rect 6685 26393 6719 26427
rect 6719 26393 6728 26427
rect 6676 26384 6728 26393
rect 23604 26384 23656 26436
rect 2168 26223 2220 26232
rect 2168 26189 2177 26223
rect 2177 26189 2211 26223
rect 2211 26189 2220 26223
rect 3916 26316 3968 26368
rect 4284 26316 4336 26368
rect 2996 26291 3048 26300
rect 2996 26257 3005 26291
rect 3005 26257 3039 26291
rect 3039 26257 3048 26291
rect 2996 26248 3048 26257
rect 12196 26248 12248 26300
rect 2168 26180 2220 26189
rect 3364 26180 3416 26232
rect 6400 26180 6452 26232
rect 7320 26180 7372 26232
rect 7688 26180 7740 26232
rect 11736 26223 11788 26232
rect 1708 26044 1760 26096
rect 7412 26112 7464 26164
rect 4192 26044 4244 26096
rect 6216 26087 6268 26096
rect 6216 26053 6225 26087
rect 6225 26053 6259 26087
rect 6259 26053 6268 26087
rect 6216 26044 6268 26053
rect 6492 26087 6544 26096
rect 6492 26053 6501 26087
rect 6501 26053 6535 26087
rect 6535 26053 6544 26087
rect 6492 26044 6544 26053
rect 7320 26044 7372 26096
rect 11736 26189 11745 26223
rect 11745 26189 11779 26223
rect 11779 26189 11788 26223
rect 17716 26316 17768 26368
rect 19280 26248 19332 26300
rect 11736 26180 11788 26189
rect 12196 26155 12248 26164
rect 12196 26121 12205 26155
rect 12205 26121 12239 26155
rect 12239 26121 12248 26155
rect 12196 26112 12248 26121
rect 12472 26112 12524 26164
rect 14864 26112 14916 26164
rect 9068 26044 9120 26096
rect 16520 26180 16572 26232
rect 17716 26223 17768 26232
rect 17716 26189 17725 26223
rect 17725 26189 17759 26223
rect 17759 26189 17768 26223
rect 17716 26180 17768 26189
rect 23696 26248 23748 26300
rect 24064 26291 24116 26300
rect 24064 26257 24073 26291
rect 24073 26257 24107 26291
rect 24107 26257 24116 26291
rect 24064 26248 24116 26257
rect 17900 26044 17952 26096
rect 18360 26044 18412 26096
rect 20476 26112 20528 26164
rect 21856 26155 21908 26164
rect 21856 26121 21865 26155
rect 21865 26121 21899 26155
rect 21899 26121 21908 26155
rect 21856 26112 21908 26121
rect 20568 26044 20620 26096
rect 23512 26087 23564 26096
rect 23512 26053 23521 26087
rect 23521 26053 23555 26087
rect 23555 26053 23564 26087
rect 23512 26044 23564 26053
rect 23696 26087 23748 26096
rect 23696 26053 23705 26087
rect 23705 26053 23739 26087
rect 23739 26053 23748 26087
rect 23696 26044 23748 26053
rect 24432 26044 24484 26096
rect 18870 25942 18922 25994
rect 18934 25942 18986 25994
rect 18998 25942 19050 25994
rect 19062 25942 19114 25994
rect 19126 25942 19178 25994
rect 7412 25883 7464 25892
rect 7412 25849 7421 25883
rect 7421 25849 7455 25883
rect 7455 25849 7464 25883
rect 7412 25840 7464 25849
rect 2168 25772 2220 25824
rect 8332 25772 8384 25824
rect 9252 25772 9304 25824
rect 11736 25815 11788 25824
rect 11736 25781 11745 25815
rect 11745 25781 11779 25815
rect 11779 25781 11788 25815
rect 11736 25772 11788 25781
rect 14864 25815 14916 25824
rect 14864 25781 14873 25815
rect 14873 25781 14907 25815
rect 14907 25781 14916 25815
rect 14864 25772 14916 25781
rect 15876 25772 15928 25824
rect 21856 25772 21908 25824
rect 972 25704 1024 25756
rect 1892 25747 1944 25756
rect 1892 25713 1901 25747
rect 1901 25713 1935 25747
rect 1935 25713 1944 25747
rect 1892 25704 1944 25713
rect 3364 25747 3416 25756
rect 3364 25713 3373 25747
rect 3373 25713 3407 25747
rect 3407 25713 3416 25747
rect 3364 25704 3416 25713
rect 4284 25747 4336 25756
rect 4284 25713 4293 25747
rect 4293 25713 4327 25747
rect 4327 25713 4336 25747
rect 4284 25704 4336 25713
rect 6400 25704 6452 25756
rect 6768 25747 6820 25756
rect 6768 25713 6777 25747
rect 6777 25713 6811 25747
rect 6811 25713 6820 25747
rect 6768 25704 6820 25713
rect 10080 25747 10132 25756
rect 5388 25636 5440 25688
rect 6216 25636 6268 25688
rect 4192 25568 4244 25620
rect 6492 25500 6544 25552
rect 7780 25500 7832 25552
rect 10080 25713 10089 25747
rect 10089 25713 10123 25747
rect 10123 25713 10132 25747
rect 10080 25704 10132 25713
rect 10264 25704 10316 25756
rect 12380 25704 12432 25756
rect 18360 25704 18412 25756
rect 19648 25704 19700 25756
rect 9160 25636 9212 25688
rect 11092 25636 11144 25688
rect 12564 25679 12616 25688
rect 12564 25645 12573 25679
rect 12573 25645 12607 25679
rect 12607 25645 12616 25679
rect 12564 25636 12616 25645
rect 14220 25636 14272 25688
rect 14404 25636 14456 25688
rect 15232 25636 15284 25688
rect 16152 25636 16204 25688
rect 17624 25636 17676 25688
rect 19004 25679 19056 25688
rect 17716 25568 17768 25620
rect 19004 25645 19013 25679
rect 19013 25645 19047 25679
rect 19047 25645 19056 25679
rect 19004 25636 19056 25645
rect 20844 25679 20896 25688
rect 20844 25645 20853 25679
rect 20853 25645 20887 25679
rect 20887 25645 20896 25679
rect 20844 25636 20896 25645
rect 21120 25679 21172 25688
rect 21120 25645 21129 25679
rect 21129 25645 21163 25679
rect 21163 25645 21172 25679
rect 21120 25636 21172 25645
rect 22868 25679 22920 25688
rect 22868 25645 22877 25679
rect 22877 25645 22911 25679
rect 22911 25645 22920 25679
rect 22868 25636 22920 25645
rect 19464 25568 19516 25620
rect 20660 25611 20712 25620
rect 20660 25577 20669 25611
rect 20669 25577 20703 25611
rect 20703 25577 20712 25611
rect 20660 25568 20712 25577
rect 8424 25500 8476 25552
rect 16796 25500 16848 25552
rect 19004 25500 19056 25552
rect 20476 25543 20528 25552
rect 20476 25509 20485 25543
rect 20485 25509 20519 25543
rect 20519 25509 20528 25543
rect 20476 25500 20528 25509
rect 24248 25500 24300 25552
rect 3510 25398 3562 25450
rect 3574 25398 3626 25450
rect 3638 25398 3690 25450
rect 3702 25398 3754 25450
rect 3766 25398 3818 25450
rect 2996 25339 3048 25348
rect 2996 25305 3005 25339
rect 3005 25305 3039 25339
rect 3039 25305 3048 25339
rect 2996 25296 3048 25305
rect 3364 25339 3416 25348
rect 3364 25305 3373 25339
rect 3373 25305 3407 25339
rect 3407 25305 3416 25339
rect 3364 25296 3416 25305
rect 3916 25296 3968 25348
rect 4284 25296 4336 25348
rect 6768 25296 6820 25348
rect 7780 25339 7832 25348
rect 7780 25305 7789 25339
rect 7789 25305 7823 25339
rect 7823 25305 7832 25339
rect 7780 25296 7832 25305
rect 10080 25296 10132 25348
rect 12564 25296 12616 25348
rect 14864 25296 14916 25348
rect 15876 25339 15928 25348
rect 1708 25203 1760 25212
rect 1708 25169 1717 25203
rect 1717 25169 1751 25203
rect 1751 25169 1760 25203
rect 1708 25160 1760 25169
rect 972 25092 1024 25144
rect 6216 25135 6268 25144
rect 6216 25101 6225 25135
rect 6225 25101 6259 25135
rect 6259 25101 6268 25135
rect 6216 25092 6268 25101
rect 6676 25092 6728 25144
rect 7412 25092 7464 25144
rect 1892 25024 1944 25076
rect 4192 25024 4244 25076
rect 10448 25228 10500 25280
rect 15232 25228 15284 25280
rect 9068 25203 9120 25212
rect 9068 25169 9077 25203
rect 9077 25169 9111 25203
rect 9111 25169 9120 25203
rect 9068 25160 9120 25169
rect 10264 25160 10316 25212
rect 15876 25305 15885 25339
rect 15885 25305 15919 25339
rect 15919 25305 15928 25339
rect 15876 25296 15928 25305
rect 16796 25339 16848 25348
rect 16796 25305 16805 25339
rect 16805 25305 16839 25339
rect 16839 25305 16848 25339
rect 16796 25296 16848 25305
rect 19464 25339 19516 25348
rect 19464 25305 19473 25339
rect 19473 25305 19507 25339
rect 19507 25305 19516 25339
rect 19464 25296 19516 25305
rect 21948 25339 22000 25348
rect 21948 25305 21957 25339
rect 21957 25305 21991 25339
rect 21991 25305 22000 25339
rect 21948 25296 22000 25305
rect 22868 25296 22920 25348
rect 9252 25135 9304 25144
rect 9252 25101 9261 25135
rect 9261 25101 9295 25135
rect 9295 25101 9304 25135
rect 9252 25092 9304 25101
rect 9804 25092 9856 25144
rect 11736 25135 11788 25144
rect 5388 24999 5440 25008
rect 5388 24965 5397 24999
rect 5397 24965 5431 24999
rect 5431 24965 5440 24999
rect 5388 24956 5440 24965
rect 5480 24956 5532 25008
rect 6952 24956 7004 25008
rect 9160 25024 9212 25076
rect 11736 25101 11745 25135
rect 11745 25101 11779 25135
rect 11779 25101 11788 25135
rect 11736 25092 11788 25101
rect 12196 25092 12248 25144
rect 14956 25092 15008 25144
rect 16520 25228 16572 25280
rect 21120 25271 21172 25280
rect 21120 25237 21129 25271
rect 21129 25237 21163 25271
rect 21163 25237 21172 25271
rect 21120 25228 21172 25237
rect 17624 25203 17676 25212
rect 17624 25169 17633 25203
rect 17633 25169 17667 25203
rect 17667 25169 17676 25203
rect 17624 25160 17676 25169
rect 17992 25160 18044 25212
rect 17348 25135 17400 25144
rect 17348 25101 17357 25135
rect 17357 25101 17391 25135
rect 17391 25101 17400 25135
rect 17348 25092 17400 25101
rect 20476 25135 20528 25144
rect 20476 25101 20485 25135
rect 20485 25101 20519 25135
rect 20519 25101 20528 25135
rect 20476 25092 20528 25101
rect 20660 25092 20712 25144
rect 22408 25160 22460 25212
rect 24156 25160 24208 25212
rect 23420 25092 23472 25144
rect 12564 25024 12616 25076
rect 14404 25024 14456 25076
rect 18360 25024 18412 25076
rect 19004 25024 19056 25076
rect 20568 25024 20620 25076
rect 24248 25024 24300 25076
rect 24708 25024 24760 25076
rect 8424 24956 8476 25008
rect 11092 24999 11144 25008
rect 11092 24965 11101 24999
rect 11101 24965 11135 24999
rect 11135 24965 11144 24999
rect 11092 24956 11144 24965
rect 12380 24956 12432 25008
rect 19648 24999 19700 25008
rect 19648 24965 19657 24999
rect 19657 24965 19691 24999
rect 19691 24965 19700 24999
rect 19648 24956 19700 24965
rect 23512 24999 23564 25008
rect 23512 24965 23521 24999
rect 23521 24965 23555 24999
rect 23555 24965 23564 24999
rect 23512 24956 23564 24965
rect 18870 24854 18922 24906
rect 18934 24854 18986 24906
rect 18998 24854 19050 24906
rect 19062 24854 19114 24906
rect 19126 24854 19178 24906
rect 880 24795 932 24804
rect 880 24761 889 24795
rect 889 24761 923 24795
rect 923 24761 932 24795
rect 880 24752 932 24761
rect 1892 24752 1944 24804
rect 6216 24752 6268 24804
rect 6952 24795 7004 24804
rect 6952 24761 6961 24795
rect 6961 24761 6995 24795
rect 6995 24761 7004 24795
rect 6952 24752 7004 24761
rect 7412 24795 7464 24804
rect 7412 24761 7421 24795
rect 7421 24761 7455 24795
rect 7455 24761 7464 24795
rect 7412 24752 7464 24761
rect 11736 24795 11788 24804
rect 11736 24761 11745 24795
rect 11745 24761 11779 24795
rect 11779 24761 11788 24795
rect 11736 24752 11788 24761
rect 2168 24684 2220 24736
rect 10448 24727 10500 24736
rect 10448 24693 10457 24727
rect 10457 24693 10491 24727
rect 10491 24693 10500 24727
rect 10448 24684 10500 24693
rect 11368 24727 11420 24736
rect 11368 24693 11377 24727
rect 11377 24693 11411 24727
rect 11411 24693 11420 24727
rect 12196 24752 12248 24804
rect 12472 24752 12524 24804
rect 20844 24752 20896 24804
rect 23236 24752 23288 24804
rect 23512 24752 23564 24804
rect 24064 24752 24116 24804
rect 11368 24684 11420 24693
rect 4192 24659 4244 24668
rect 4192 24625 4201 24659
rect 4201 24625 4235 24659
rect 4235 24625 4244 24659
rect 4192 24616 4244 24625
rect 5480 24616 5532 24668
rect 6400 24659 6452 24668
rect 6400 24625 6409 24659
rect 6409 24625 6443 24659
rect 6443 24625 6452 24659
rect 6400 24616 6452 24625
rect 12564 24659 12616 24668
rect 12564 24625 12573 24659
rect 12573 24625 12607 24659
rect 12607 24625 12616 24659
rect 12564 24616 12616 24625
rect 14956 24616 15008 24668
rect 18452 24659 18504 24668
rect 18452 24625 18461 24659
rect 18461 24625 18495 24659
rect 18495 24625 18504 24659
rect 18452 24616 18504 24625
rect 18820 24659 18872 24668
rect 18820 24625 18829 24659
rect 18829 24625 18863 24659
rect 18863 24625 18872 24659
rect 18820 24616 18872 24625
rect 5572 24591 5624 24600
rect 5572 24557 5581 24591
rect 5581 24557 5615 24591
rect 5615 24557 5624 24591
rect 5572 24548 5624 24557
rect 5664 24591 5716 24600
rect 5664 24557 5673 24591
rect 5673 24557 5707 24591
rect 5707 24557 5716 24591
rect 6492 24591 6544 24600
rect 5664 24548 5716 24557
rect 6492 24557 6501 24591
rect 6501 24557 6535 24591
rect 6535 24557 6544 24591
rect 6492 24548 6544 24557
rect 9252 24591 9304 24600
rect 9252 24557 9261 24591
rect 9261 24557 9295 24591
rect 9295 24557 9304 24591
rect 9252 24548 9304 24557
rect 9988 24591 10040 24600
rect 9988 24557 9997 24591
rect 9997 24557 10031 24591
rect 10031 24557 10040 24591
rect 9988 24548 10040 24557
rect 15140 24591 15192 24600
rect 1064 24455 1116 24464
rect 1064 24421 1073 24455
rect 1073 24421 1107 24455
rect 1107 24421 1116 24455
rect 1064 24412 1116 24421
rect 4284 24455 4336 24464
rect 4284 24421 4293 24455
rect 4293 24421 4327 24455
rect 4327 24421 4336 24455
rect 4284 24412 4336 24421
rect 7504 24455 7556 24464
rect 7504 24421 7513 24455
rect 7513 24421 7547 24455
rect 7547 24421 7556 24455
rect 7504 24412 7556 24421
rect 7964 24412 8016 24464
rect 9804 24412 9856 24464
rect 15140 24557 15149 24591
rect 15149 24557 15183 24591
rect 15183 24557 15192 24591
rect 15140 24548 15192 24557
rect 17992 24548 18044 24600
rect 18728 24548 18780 24600
rect 19648 24616 19700 24668
rect 21488 24616 21540 24668
rect 22868 24616 22920 24668
rect 24432 24659 24484 24668
rect 24432 24625 24441 24659
rect 24441 24625 24475 24659
rect 24475 24625 24484 24659
rect 24432 24616 24484 24625
rect 20568 24548 20620 24600
rect 24708 24591 24760 24600
rect 24708 24557 24717 24591
rect 24717 24557 24751 24591
rect 24751 24557 24760 24591
rect 24708 24548 24760 24557
rect 20752 24480 20804 24532
rect 11460 24455 11512 24464
rect 11460 24421 11469 24455
rect 11469 24421 11503 24455
rect 11503 24421 11512 24455
rect 11460 24412 11512 24421
rect 16428 24412 16480 24464
rect 17348 24455 17400 24464
rect 17348 24421 17357 24455
rect 17357 24421 17391 24455
rect 17391 24421 17400 24455
rect 17348 24412 17400 24421
rect 17900 24455 17952 24464
rect 17900 24421 17909 24455
rect 17909 24421 17943 24455
rect 17943 24421 17952 24455
rect 17900 24412 17952 24421
rect 18544 24412 18596 24464
rect 20660 24455 20712 24464
rect 20660 24421 20669 24455
rect 20669 24421 20703 24455
rect 20703 24421 20712 24455
rect 20660 24412 20712 24421
rect 21028 24412 21080 24464
rect 21396 24412 21448 24464
rect 22408 24455 22460 24464
rect 22408 24421 22417 24455
rect 22417 24421 22451 24455
rect 22451 24421 22460 24455
rect 22408 24412 22460 24421
rect 3510 24310 3562 24362
rect 3574 24310 3626 24362
rect 3638 24310 3690 24362
rect 3702 24310 3754 24362
rect 3766 24310 3818 24362
rect 3916 24208 3968 24260
rect 4284 24251 4336 24260
rect 4284 24217 4293 24251
rect 4293 24217 4327 24251
rect 4327 24217 4336 24251
rect 4284 24208 4336 24217
rect 5664 24208 5716 24260
rect 6952 24208 7004 24260
rect 7504 24208 7556 24260
rect 9988 24251 10040 24260
rect 9988 24217 9997 24251
rect 9997 24217 10031 24251
rect 10031 24217 10040 24251
rect 9988 24208 10040 24217
rect 11460 24208 11512 24260
rect 12472 24251 12524 24260
rect 12472 24217 12481 24251
rect 12481 24217 12515 24251
rect 12515 24217 12524 24251
rect 12472 24208 12524 24217
rect 12564 24251 12616 24260
rect 12564 24217 12573 24251
rect 12573 24217 12607 24251
rect 12607 24217 12616 24251
rect 18452 24251 18504 24260
rect 12564 24208 12616 24217
rect 18452 24217 18461 24251
rect 18461 24217 18495 24251
rect 18495 24217 18504 24251
rect 18452 24208 18504 24217
rect 18544 24251 18596 24260
rect 18544 24217 18553 24251
rect 18553 24217 18587 24251
rect 18587 24217 18596 24251
rect 18544 24208 18596 24217
rect 21488 24208 21540 24260
rect 22868 24208 22920 24260
rect 23604 24251 23656 24260
rect 23604 24217 23613 24251
rect 23613 24217 23647 24251
rect 23647 24217 23656 24251
rect 23604 24208 23656 24217
rect 880 24140 932 24192
rect 4192 24183 4244 24192
rect 1064 24115 1116 24124
rect 1064 24081 1073 24115
rect 1073 24081 1107 24115
rect 1107 24081 1116 24115
rect 1064 24072 1116 24081
rect 4192 24149 4201 24183
rect 4201 24149 4235 24183
rect 4235 24149 4244 24183
rect 4192 24140 4244 24149
rect 5572 24140 5624 24192
rect 7412 24140 7464 24192
rect 10448 24183 10500 24192
rect 10448 24149 10457 24183
rect 10457 24149 10491 24183
rect 10491 24149 10500 24183
rect 10448 24140 10500 24149
rect 11368 24183 11420 24192
rect 11368 24149 11377 24183
rect 11377 24149 11411 24183
rect 11411 24149 11420 24183
rect 11368 24140 11420 24149
rect 18728 24140 18780 24192
rect 20476 24140 20528 24192
rect 20660 24183 20712 24192
rect 20660 24149 20669 24183
rect 20669 24149 20703 24183
rect 20703 24149 20712 24183
rect 20660 24140 20712 24149
rect 22408 24183 22460 24192
rect 22408 24149 22417 24183
rect 22417 24149 22451 24183
rect 22451 24149 22460 24183
rect 22408 24140 22460 24149
rect 6492 24072 6544 24124
rect 15140 24072 15192 24124
rect 16428 24115 16480 24124
rect 16428 24081 16437 24115
rect 16437 24081 16471 24115
rect 16471 24081 16480 24115
rect 16428 24072 16480 24081
rect 18820 24072 18872 24124
rect 20752 24072 20804 24124
rect 788 24004 840 24056
rect 1524 24004 1576 24056
rect 5480 24047 5532 24056
rect 5480 24013 5489 24047
rect 5489 24013 5523 24047
rect 5523 24013 5532 24047
rect 5480 24004 5532 24013
rect 7412 24047 7464 24056
rect 7412 24013 7421 24047
rect 7421 24013 7455 24047
rect 7455 24013 7464 24047
rect 7412 24004 7464 24013
rect 8424 24047 8476 24056
rect 8424 24013 8433 24047
rect 8433 24013 8467 24047
rect 8467 24013 8476 24047
rect 8424 24004 8476 24013
rect 14404 24047 14456 24056
rect 14404 24013 14413 24047
rect 14413 24013 14447 24047
rect 14447 24013 14456 24047
rect 14404 24004 14456 24013
rect 21028 24004 21080 24056
rect 2168 23936 2220 23988
rect 9068 23979 9120 23988
rect 9068 23945 9077 23979
rect 9077 23945 9111 23979
rect 9111 23945 9120 23979
rect 9068 23936 9120 23945
rect 15140 23936 15192 23988
rect 20476 23936 20528 23988
rect 24064 24004 24116 24056
rect 23420 23936 23472 23988
rect 16520 23868 16572 23920
rect 16888 23868 16940 23920
rect 17992 23911 18044 23920
rect 17992 23877 18001 23911
rect 18001 23877 18035 23911
rect 18035 23877 18044 23911
rect 17992 23868 18044 23877
rect 21396 23868 21448 23920
rect 24432 23868 24484 23920
rect 18870 23766 18922 23818
rect 18934 23766 18986 23818
rect 18998 23766 19050 23818
rect 19062 23766 19114 23818
rect 19126 23766 19178 23818
rect 14956 23707 15008 23716
rect 14956 23673 14965 23707
rect 14965 23673 14999 23707
rect 14999 23673 15008 23707
rect 14956 23664 15008 23673
rect 15140 23707 15192 23716
rect 15140 23673 15149 23707
rect 15149 23673 15183 23707
rect 15183 23673 15192 23707
rect 15140 23664 15192 23673
rect 18360 23707 18412 23716
rect 18360 23673 18369 23707
rect 18369 23673 18403 23707
rect 18403 23673 18412 23707
rect 18360 23664 18412 23673
rect 21488 23707 21540 23716
rect 21488 23673 21497 23707
rect 21497 23673 21531 23707
rect 21531 23673 21540 23707
rect 21488 23664 21540 23673
rect 24708 23664 24760 23716
rect 7504 23596 7556 23648
rect 12472 23596 12524 23648
rect 1064 23528 1116 23580
rect 1892 23528 1944 23580
rect 4192 23571 4244 23580
rect 4192 23537 4201 23571
rect 4201 23537 4235 23571
rect 4235 23537 4244 23571
rect 4192 23528 4244 23537
rect 4284 23528 4336 23580
rect 13392 23571 13444 23580
rect 13392 23537 13401 23571
rect 13401 23537 13435 23571
rect 13435 23537 13444 23571
rect 16244 23596 16296 23648
rect 13392 23528 13444 23537
rect 15968 23528 16020 23580
rect 16428 23528 16480 23580
rect 18084 23571 18136 23580
rect 18084 23537 18093 23571
rect 18093 23537 18127 23571
rect 18127 23537 18136 23571
rect 18084 23528 18136 23537
rect 18636 23571 18688 23580
rect 18636 23537 18645 23571
rect 18645 23537 18679 23571
rect 18679 23537 18688 23571
rect 18636 23528 18688 23537
rect 20568 23571 20620 23580
rect 20568 23537 20577 23571
rect 20577 23537 20611 23571
rect 20611 23537 20620 23571
rect 20568 23528 20620 23537
rect 20660 23571 20712 23580
rect 20660 23537 20669 23571
rect 20669 23537 20703 23571
rect 20703 23537 20712 23571
rect 20660 23528 20712 23537
rect 1800 23503 1852 23512
rect 1800 23469 1809 23503
rect 1809 23469 1843 23503
rect 1843 23469 1852 23503
rect 1800 23460 1852 23469
rect 5756 23503 5808 23512
rect 5756 23469 5765 23503
rect 5765 23469 5799 23503
rect 5799 23469 5808 23503
rect 5756 23460 5808 23469
rect 7412 23460 7464 23512
rect 12288 23460 12340 23512
rect 12564 23503 12616 23512
rect 12564 23469 12573 23503
rect 12573 23469 12607 23503
rect 12607 23469 12616 23503
rect 12564 23460 12616 23469
rect 20936 23460 20988 23512
rect 7964 23435 8016 23444
rect 7964 23401 7973 23435
rect 7973 23401 8007 23435
rect 8007 23401 8016 23435
rect 7964 23392 8016 23401
rect 788 23324 840 23376
rect 1156 23324 1208 23376
rect 1984 23367 2036 23376
rect 1984 23333 1993 23367
rect 1993 23333 2027 23367
rect 2027 23333 2036 23367
rect 1984 23324 2036 23333
rect 16704 23324 16756 23376
rect 20844 23367 20896 23376
rect 20844 23333 20853 23367
rect 20853 23333 20887 23367
rect 20887 23333 20896 23367
rect 20844 23324 20896 23333
rect 24156 23367 24208 23376
rect 24156 23333 24165 23367
rect 24165 23333 24199 23367
rect 24199 23333 24208 23367
rect 24156 23324 24208 23333
rect 3510 23222 3562 23274
rect 3574 23222 3626 23274
rect 3638 23222 3690 23274
rect 3702 23222 3754 23274
rect 3766 23222 3818 23274
rect 1064 23163 1116 23172
rect 1064 23129 1073 23163
rect 1073 23129 1107 23163
rect 1107 23129 1116 23163
rect 1064 23120 1116 23129
rect 4192 23163 4244 23172
rect 4192 23129 4201 23163
rect 4201 23129 4235 23163
rect 4235 23129 4244 23163
rect 4192 23120 4244 23129
rect 1800 23052 1852 23104
rect 4284 23052 4336 23104
rect 5664 23120 5716 23172
rect 7504 23120 7556 23172
rect 13392 23120 13444 23172
rect 16704 23163 16756 23172
rect 16704 23129 16713 23163
rect 16713 23129 16747 23163
rect 16747 23129 16756 23163
rect 16704 23120 16756 23129
rect 18360 23163 18412 23172
rect 18360 23129 18369 23163
rect 18369 23129 18403 23163
rect 18403 23129 18412 23163
rect 18360 23120 18412 23129
rect 18728 23120 18780 23172
rect 20660 23120 20712 23172
rect 20936 23163 20988 23172
rect 20936 23129 20945 23163
rect 20945 23129 20979 23163
rect 20979 23129 20988 23163
rect 20936 23120 20988 23129
rect 9804 23095 9856 23104
rect 9804 23061 9813 23095
rect 9813 23061 9847 23095
rect 9847 23061 9856 23095
rect 9804 23052 9856 23061
rect 7412 22984 7464 23036
rect 11828 22984 11880 23036
rect 24156 23027 24208 23036
rect 1064 22916 1116 22968
rect 1984 22916 2036 22968
rect 5756 22916 5808 22968
rect 7964 22959 8016 22968
rect 7964 22925 7973 22959
rect 7973 22925 8007 22959
rect 8007 22925 8016 22959
rect 7964 22916 8016 22925
rect 9068 22916 9120 22968
rect 12012 22916 12064 22968
rect 12564 22959 12616 22968
rect 12564 22925 12573 22959
rect 12573 22925 12607 22959
rect 12607 22925 12616 22959
rect 12564 22916 12616 22925
rect 13484 22916 13536 22968
rect 15876 22916 15928 22968
rect 16152 22916 16204 22968
rect 18084 22916 18136 22968
rect 18544 22959 18596 22968
rect 18544 22925 18553 22959
rect 18553 22925 18587 22959
rect 18587 22925 18596 22959
rect 18544 22916 18596 22925
rect 18636 22959 18688 22968
rect 18636 22925 18645 22959
rect 18645 22925 18679 22959
rect 18679 22925 18688 22959
rect 18636 22916 18688 22925
rect 23236 22916 23288 22968
rect 24156 22993 24165 23027
rect 24165 22993 24199 23027
rect 24199 22993 24208 23027
rect 24156 22984 24208 22993
rect 24432 22984 24484 23036
rect 1892 22891 1944 22900
rect 1892 22857 1901 22891
rect 1901 22857 1935 22891
rect 1935 22857 1944 22891
rect 1892 22848 1944 22857
rect 5204 22891 5256 22900
rect 5204 22857 5213 22891
rect 5213 22857 5247 22891
rect 5247 22857 5256 22891
rect 5204 22848 5256 22857
rect 8884 22848 8936 22900
rect 11000 22848 11052 22900
rect 13116 22891 13168 22900
rect 13116 22857 13125 22891
rect 13125 22857 13159 22891
rect 13159 22857 13168 22891
rect 13116 22848 13168 22857
rect 16428 22891 16480 22900
rect 16428 22857 16437 22891
rect 16437 22857 16471 22891
rect 16471 22857 16480 22891
rect 16428 22848 16480 22857
rect 21672 22848 21724 22900
rect 24432 22891 24484 22900
rect 24432 22857 24441 22891
rect 24441 22857 24475 22891
rect 24475 22857 24484 22891
rect 24432 22848 24484 22857
rect 24708 22848 24760 22900
rect 12012 22823 12064 22832
rect 12012 22789 12021 22823
rect 12021 22789 12055 22823
rect 12055 22789 12064 22823
rect 12012 22780 12064 22789
rect 12288 22823 12340 22832
rect 12288 22789 12297 22823
rect 12297 22789 12331 22823
rect 12331 22789 12340 22823
rect 12288 22780 12340 22789
rect 15968 22823 16020 22832
rect 15968 22789 15977 22823
rect 15977 22789 16011 22823
rect 16011 22789 16020 22823
rect 15968 22780 16020 22789
rect 20844 22823 20896 22832
rect 20844 22789 20853 22823
rect 20853 22789 20887 22823
rect 20887 22789 20896 22823
rect 20844 22780 20896 22789
rect 18870 22678 18922 22730
rect 18934 22678 18986 22730
rect 18998 22678 19050 22730
rect 19062 22678 19114 22730
rect 19126 22678 19178 22730
rect 1800 22576 1852 22628
rect 2168 22619 2220 22628
rect 2168 22585 2177 22619
rect 2177 22585 2211 22619
rect 2211 22585 2220 22619
rect 2168 22576 2220 22585
rect 18544 22619 18596 22628
rect 18544 22585 18553 22619
rect 18553 22585 18587 22619
rect 18587 22585 18596 22619
rect 18544 22576 18596 22585
rect 24248 22619 24300 22628
rect 24248 22585 24257 22619
rect 24257 22585 24291 22619
rect 24291 22585 24300 22619
rect 24248 22576 24300 22585
rect 5204 22551 5256 22560
rect 5204 22517 5213 22551
rect 5213 22517 5247 22551
rect 5247 22517 5256 22551
rect 5204 22508 5256 22517
rect 17716 22508 17768 22560
rect 24708 22551 24760 22560
rect 24708 22517 24717 22551
rect 24717 22517 24751 22551
rect 24751 22517 24760 22551
rect 24708 22508 24760 22517
rect 4284 22440 4336 22492
rect 4928 22440 4980 22492
rect 11000 22483 11052 22492
rect 11000 22449 11009 22483
rect 11009 22449 11043 22483
rect 11043 22449 11052 22483
rect 11000 22440 11052 22449
rect 11368 22440 11420 22492
rect 12012 22440 12064 22492
rect 12748 22483 12800 22492
rect 12748 22449 12757 22483
rect 12757 22449 12791 22483
rect 12791 22449 12800 22483
rect 12748 22440 12800 22449
rect 16336 22483 16388 22492
rect 16336 22449 16345 22483
rect 16345 22449 16379 22483
rect 16379 22449 16388 22483
rect 16336 22440 16388 22449
rect 16888 22483 16940 22492
rect 16888 22449 16897 22483
rect 16897 22449 16931 22483
rect 16931 22449 16940 22483
rect 16888 22440 16940 22449
rect 20200 22483 20252 22492
rect 20200 22449 20209 22483
rect 20209 22449 20243 22483
rect 20243 22449 20252 22483
rect 20200 22440 20252 22449
rect 20844 22440 20896 22492
rect 22776 22483 22828 22492
rect 22776 22449 22785 22483
rect 22785 22449 22819 22483
rect 22819 22449 22828 22483
rect 22776 22440 22828 22449
rect 24432 22483 24484 22492
rect 24432 22449 24441 22483
rect 24441 22449 24475 22483
rect 24475 22449 24484 22483
rect 24432 22440 24484 22449
rect 1248 22372 1300 22424
rect 1984 22415 2036 22424
rect 1984 22381 1993 22415
rect 1993 22381 2027 22415
rect 2027 22381 2036 22415
rect 1984 22372 2036 22381
rect 13484 22372 13536 22424
rect 16428 22415 16480 22424
rect 16428 22381 16437 22415
rect 16437 22381 16471 22415
rect 16471 22381 16480 22415
rect 16428 22372 16480 22381
rect 16704 22372 16756 22424
rect 20476 22415 20528 22424
rect 20476 22381 20485 22415
rect 20485 22381 20519 22415
rect 20519 22381 20528 22415
rect 20476 22372 20528 22381
rect 22408 22372 22460 22424
rect 16520 22347 16572 22356
rect 16520 22313 16529 22347
rect 16529 22313 16563 22347
rect 16563 22313 16572 22347
rect 16520 22304 16572 22313
rect 23880 22304 23932 22356
rect 4008 22279 4060 22288
rect 4008 22245 4017 22279
rect 4017 22245 4051 22279
rect 4051 22245 4060 22279
rect 4008 22236 4060 22245
rect 7780 22279 7832 22288
rect 7780 22245 7789 22279
rect 7789 22245 7823 22279
rect 7823 22245 7832 22279
rect 7780 22236 7832 22245
rect 10816 22279 10868 22288
rect 10816 22245 10825 22279
rect 10825 22245 10859 22279
rect 10859 22245 10868 22279
rect 10816 22236 10868 22245
rect 15416 22279 15468 22288
rect 15416 22245 15425 22279
rect 15425 22245 15459 22279
rect 15459 22245 15468 22279
rect 15416 22236 15468 22245
rect 19096 22279 19148 22288
rect 19096 22245 19105 22279
rect 19105 22245 19139 22279
rect 19139 22245 19148 22279
rect 19096 22236 19148 22245
rect 21764 22279 21816 22288
rect 21764 22245 21773 22279
rect 21773 22245 21807 22279
rect 21807 22245 21816 22279
rect 21764 22236 21816 22245
rect 22592 22236 22644 22288
rect 23236 22236 23288 22288
rect 24248 22372 24300 22424
rect 3510 22134 3562 22186
rect 3574 22134 3626 22186
rect 3638 22134 3690 22186
rect 3702 22134 3754 22186
rect 3766 22134 3818 22186
rect 4008 22075 4060 22084
rect 4008 22041 4017 22075
rect 4017 22041 4051 22075
rect 4051 22041 4060 22075
rect 4008 22032 4060 22041
rect 5204 22032 5256 22084
rect 6400 22032 6452 22084
rect 8332 22032 8384 22084
rect 11368 22075 11420 22084
rect 11368 22041 11377 22075
rect 11377 22041 11411 22075
rect 11411 22041 11420 22075
rect 11368 22032 11420 22041
rect 13116 22032 13168 22084
rect 16336 22032 16388 22084
rect 16520 22075 16572 22084
rect 16520 22041 16529 22075
rect 16529 22041 16563 22075
rect 16563 22041 16572 22075
rect 16520 22032 16572 22041
rect 19096 22032 19148 22084
rect 2168 21964 2220 22016
rect 4284 21964 4336 22016
rect 2076 21871 2128 21880
rect 2076 21837 2085 21871
rect 2085 21837 2119 21871
rect 2119 21837 2128 21871
rect 2076 21828 2128 21837
rect 11000 21964 11052 22016
rect 7412 21896 7464 21948
rect 8700 21939 8752 21948
rect 8700 21905 8709 21939
rect 8709 21905 8743 21939
rect 8743 21905 8752 21939
rect 8700 21896 8752 21905
rect 10816 21939 10868 21948
rect 10816 21905 10825 21939
rect 10825 21905 10859 21939
rect 10859 21905 10868 21939
rect 10816 21896 10868 21905
rect 1248 21692 1300 21744
rect 5756 21828 5808 21880
rect 7780 21871 7832 21880
rect 7780 21837 7789 21871
rect 7789 21837 7823 21871
rect 7823 21837 7832 21871
rect 7780 21828 7832 21837
rect 8332 21828 8384 21880
rect 11736 21871 11788 21880
rect 11736 21837 11745 21871
rect 11745 21837 11779 21871
rect 11779 21837 11788 21871
rect 11736 21828 11788 21837
rect 12748 21964 12800 22016
rect 15416 22007 15468 22016
rect 15416 21973 15425 22007
rect 15425 21973 15459 22007
rect 15459 21973 15468 22007
rect 15416 21964 15468 21973
rect 16428 21964 16480 22016
rect 13484 21896 13536 21948
rect 15968 21896 16020 21948
rect 22776 22075 22828 22084
rect 22776 22041 22785 22075
rect 22785 22041 22819 22075
rect 22819 22041 22828 22075
rect 22776 22032 22828 22041
rect 22408 22007 22460 22016
rect 22408 21973 22417 22007
rect 22417 21973 22451 22007
rect 22451 21973 22460 22007
rect 22408 21964 22460 21973
rect 23236 21939 23288 21948
rect 23236 21905 23245 21939
rect 23245 21905 23279 21939
rect 23279 21905 23288 21939
rect 23236 21896 23288 21905
rect 24248 21896 24300 21948
rect 15876 21871 15928 21880
rect 4928 21803 4980 21812
rect 4928 21769 4937 21803
rect 4937 21769 4971 21803
rect 4971 21769 4980 21803
rect 4928 21760 4980 21769
rect 4560 21692 4612 21744
rect 6032 21692 6084 21744
rect 15876 21837 15885 21871
rect 15885 21837 15919 21871
rect 15919 21837 15928 21871
rect 15876 21828 15928 21837
rect 16704 21828 16756 21880
rect 19096 21871 19148 21880
rect 17164 21760 17216 21812
rect 15968 21692 16020 21744
rect 17348 21692 17400 21744
rect 19096 21837 19105 21871
rect 19105 21837 19139 21871
rect 19139 21837 19148 21871
rect 19096 21828 19148 21837
rect 20476 21828 20528 21880
rect 19372 21803 19424 21812
rect 19372 21769 19381 21803
rect 19381 21769 19415 21803
rect 19415 21769 19424 21803
rect 19372 21760 19424 21769
rect 23144 21803 23196 21812
rect 20108 21692 20160 21744
rect 23144 21769 23153 21803
rect 23153 21769 23187 21803
rect 23187 21769 23196 21803
rect 23144 21760 23196 21769
rect 24524 21760 24576 21812
rect 21764 21735 21816 21744
rect 21764 21701 21773 21735
rect 21773 21701 21807 21735
rect 21807 21701 21816 21735
rect 21764 21692 21816 21701
rect 22592 21735 22644 21744
rect 22592 21701 22601 21735
rect 22601 21701 22635 21735
rect 22635 21701 22644 21735
rect 22592 21692 22644 21701
rect 23880 21692 23932 21744
rect 18870 21590 18922 21642
rect 18934 21590 18986 21642
rect 18998 21590 19050 21642
rect 19062 21590 19114 21642
rect 19126 21590 19178 21642
rect 1984 21531 2036 21540
rect 1984 21497 1993 21531
rect 1993 21497 2027 21531
rect 2027 21497 2036 21531
rect 1984 21488 2036 21497
rect 4284 21531 4336 21540
rect 4284 21497 4293 21531
rect 4293 21497 4327 21531
rect 4327 21497 4336 21531
rect 4284 21488 4336 21497
rect 7412 21488 7464 21540
rect 11000 21488 11052 21540
rect 15876 21488 15928 21540
rect 16888 21488 16940 21540
rect 20476 21531 20528 21540
rect 20476 21497 20485 21531
rect 20485 21497 20519 21531
rect 20519 21497 20528 21531
rect 20476 21488 20528 21497
rect 2076 21420 2128 21472
rect 4928 21420 4980 21472
rect 11920 21420 11972 21472
rect 20200 21420 20252 21472
rect 24432 21488 24484 21540
rect 24708 21531 24760 21540
rect 24708 21497 24717 21531
rect 24717 21497 24751 21531
rect 24751 21497 24760 21531
rect 24708 21488 24760 21497
rect 22776 21420 22828 21472
rect 23144 21420 23196 21472
rect 1892 21395 1944 21404
rect 1892 21361 1901 21395
rect 1901 21361 1935 21395
rect 1935 21361 1944 21395
rect 1892 21352 1944 21361
rect 4008 21352 4060 21404
rect 4744 21352 4796 21404
rect 7688 21352 7740 21404
rect 9252 21395 9304 21404
rect 9252 21361 9261 21395
rect 9261 21361 9295 21395
rect 9295 21361 9304 21395
rect 9252 21352 9304 21361
rect 9436 21395 9488 21404
rect 9436 21361 9445 21395
rect 9445 21361 9479 21395
rect 9479 21361 9488 21395
rect 9436 21352 9488 21361
rect 11828 21352 11880 21404
rect 13300 21352 13352 21404
rect 16428 21395 16480 21404
rect 16428 21361 16437 21395
rect 16437 21361 16471 21395
rect 16471 21361 16480 21395
rect 16428 21352 16480 21361
rect 16704 21395 16756 21404
rect 16704 21361 16713 21395
rect 16713 21361 16747 21395
rect 16747 21361 16756 21395
rect 16704 21352 16756 21361
rect 17164 21395 17216 21404
rect 17164 21361 17173 21395
rect 17173 21361 17207 21395
rect 17207 21361 17216 21395
rect 17164 21352 17216 21361
rect 21304 21395 21356 21404
rect 4560 21327 4612 21336
rect 4560 21293 4569 21327
rect 4569 21293 4603 21327
rect 4603 21293 4612 21327
rect 4560 21284 4612 21293
rect 12104 21284 12156 21336
rect 12196 21216 12248 21268
rect 1248 21148 1300 21200
rect 9528 21191 9580 21200
rect 9528 21157 9537 21191
rect 9537 21157 9571 21191
rect 9571 21157 9580 21191
rect 9528 21148 9580 21157
rect 13576 21191 13628 21200
rect 13576 21157 13585 21191
rect 13585 21157 13619 21191
rect 13619 21157 13628 21191
rect 13576 21148 13628 21157
rect 16796 21284 16848 21336
rect 21304 21361 21313 21395
rect 21313 21361 21347 21395
rect 21347 21361 21356 21395
rect 21304 21352 21356 21361
rect 21672 21395 21724 21404
rect 21672 21361 21681 21395
rect 21681 21361 21715 21395
rect 21715 21361 21724 21395
rect 21672 21352 21724 21361
rect 22592 21352 22644 21404
rect 23512 21352 23564 21404
rect 23696 21395 23748 21404
rect 23696 21361 23705 21395
rect 23705 21361 23739 21395
rect 23739 21361 23748 21395
rect 23696 21352 23748 21361
rect 21212 21327 21264 21336
rect 21212 21293 21221 21327
rect 21221 21293 21255 21327
rect 21255 21293 21264 21327
rect 21212 21284 21264 21293
rect 21764 21327 21816 21336
rect 21764 21293 21773 21327
rect 21773 21293 21807 21327
rect 21807 21293 21816 21327
rect 21764 21284 21816 21293
rect 23144 21284 23196 21336
rect 23420 21284 23472 21336
rect 16980 21216 17032 21268
rect 23328 21216 23380 21268
rect 18268 21148 18320 21200
rect 20108 21148 20160 21200
rect 20752 21191 20804 21200
rect 20752 21157 20761 21191
rect 20761 21157 20795 21191
rect 20795 21157 20804 21191
rect 20752 21148 20804 21157
rect 24616 21148 24668 21200
rect 3510 21046 3562 21098
rect 3574 21046 3626 21098
rect 3638 21046 3690 21098
rect 3702 21046 3754 21098
rect 3766 21046 3818 21098
rect 1892 20987 1944 20996
rect 1892 20953 1901 20987
rect 1901 20953 1935 20987
rect 1935 20953 1944 20987
rect 1892 20944 1944 20953
rect 1984 20944 2036 20996
rect 4744 20987 4796 20996
rect 4744 20953 4753 20987
rect 4753 20953 4787 20987
rect 4787 20953 4796 20987
rect 4744 20944 4796 20953
rect 4928 20987 4980 20996
rect 4928 20953 4937 20987
rect 4937 20953 4971 20987
rect 4971 20953 4980 20987
rect 4928 20944 4980 20953
rect 9252 20944 9304 20996
rect 9528 20944 9580 20996
rect 12196 20987 12248 20996
rect 12196 20953 12205 20987
rect 12205 20953 12239 20987
rect 12239 20953 12248 20987
rect 12196 20944 12248 20953
rect 13300 20987 13352 20996
rect 13300 20953 13309 20987
rect 13309 20953 13343 20987
rect 13343 20953 13352 20987
rect 13300 20944 13352 20953
rect 16428 20944 16480 20996
rect 17164 20944 17216 20996
rect 19372 20944 19424 20996
rect 21764 20944 21816 20996
rect 22776 20987 22828 20996
rect 22776 20953 22785 20987
rect 22785 20953 22819 20987
rect 22819 20953 22828 20987
rect 22776 20944 22828 20953
rect 23512 20987 23564 20996
rect 23512 20953 23521 20987
rect 23521 20953 23555 20987
rect 23555 20953 23564 20987
rect 23512 20944 23564 20953
rect 12104 20919 12156 20928
rect 12104 20885 12113 20919
rect 12113 20885 12147 20919
rect 12147 20885 12156 20919
rect 12104 20876 12156 20885
rect 16980 20919 17032 20928
rect 16980 20885 16989 20919
rect 16989 20885 17023 20919
rect 17023 20885 17032 20919
rect 16980 20876 17032 20885
rect 4560 20808 4612 20860
rect 10172 20808 10224 20860
rect 13576 20783 13628 20792
rect 7044 20672 7096 20724
rect 6216 20604 6268 20656
rect 13576 20749 13585 20783
rect 13585 20749 13619 20783
rect 13619 20749 13628 20783
rect 13576 20740 13628 20749
rect 16704 20808 16756 20860
rect 24524 20808 24576 20860
rect 9528 20672 9580 20724
rect 11920 20672 11972 20724
rect 13760 20672 13812 20724
rect 11828 20647 11880 20656
rect 11828 20613 11837 20647
rect 11837 20613 11871 20647
rect 11871 20613 11880 20647
rect 11828 20604 11880 20613
rect 13300 20604 13352 20656
rect 20752 20740 20804 20792
rect 24616 20783 24668 20792
rect 24616 20749 24625 20783
rect 24625 20749 24659 20783
rect 24659 20749 24668 20783
rect 24616 20740 24668 20749
rect 20292 20672 20344 20724
rect 21672 20672 21724 20724
rect 22040 20672 22092 20724
rect 23696 20672 23748 20724
rect 24156 20672 24208 20724
rect 16796 20647 16848 20656
rect 16796 20613 16805 20647
rect 16805 20613 16839 20647
rect 16839 20613 16848 20647
rect 16796 20604 16848 20613
rect 18360 20604 18412 20656
rect 21212 20604 21264 20656
rect 21396 20604 21448 20656
rect 23144 20647 23196 20656
rect 23144 20613 23153 20647
rect 23153 20613 23187 20647
rect 23187 20613 23196 20647
rect 23144 20604 23196 20613
rect 23328 20647 23380 20656
rect 23328 20613 23337 20647
rect 23337 20613 23371 20647
rect 23371 20613 23380 20647
rect 23328 20604 23380 20613
rect 25168 20647 25220 20656
rect 25168 20613 25177 20647
rect 25177 20613 25211 20647
rect 25211 20613 25220 20647
rect 25168 20604 25220 20613
rect 18870 20502 18922 20554
rect 18934 20502 18986 20554
rect 18998 20502 19050 20554
rect 19062 20502 19114 20554
rect 19126 20502 19178 20554
rect 6400 20400 6452 20452
rect 7780 20400 7832 20452
rect 8148 20443 8200 20452
rect 8148 20409 8157 20443
rect 8157 20409 8191 20443
rect 8191 20409 8200 20443
rect 8148 20400 8200 20409
rect 11092 20400 11144 20452
rect 23236 20400 23288 20452
rect 1248 20264 1300 20316
rect 1524 20264 1576 20316
rect 788 20239 840 20248
rect 788 20205 797 20239
rect 797 20205 831 20239
rect 831 20205 840 20239
rect 788 20196 840 20205
rect 972 20196 1024 20248
rect 4560 20264 4612 20316
rect 5480 20307 5532 20316
rect 5480 20273 5489 20307
rect 5489 20273 5523 20307
rect 5523 20273 5532 20307
rect 5480 20264 5532 20273
rect 7044 20307 7096 20316
rect 7044 20273 7053 20307
rect 7053 20273 7087 20307
rect 7087 20273 7096 20307
rect 7044 20264 7096 20273
rect 4376 20103 4428 20112
rect 4376 20069 4385 20103
rect 4385 20069 4419 20103
rect 4419 20069 4428 20103
rect 4376 20060 4428 20069
rect 5756 20196 5808 20248
rect 5940 20196 5992 20248
rect 10264 20332 10316 20384
rect 13576 20332 13628 20384
rect 15416 20332 15468 20384
rect 9436 20307 9488 20316
rect 9436 20273 9445 20307
rect 9445 20273 9479 20307
rect 9479 20273 9488 20307
rect 9436 20264 9488 20273
rect 13484 20307 13536 20316
rect 7688 20239 7740 20248
rect 7688 20205 7697 20239
rect 7697 20205 7731 20239
rect 7731 20205 7740 20239
rect 7688 20196 7740 20205
rect 9344 20196 9396 20248
rect 13484 20273 13493 20307
rect 13493 20273 13527 20307
rect 13527 20273 13536 20307
rect 13484 20264 13536 20273
rect 16428 20332 16480 20384
rect 21764 20375 21816 20384
rect 21764 20341 21773 20375
rect 21773 20341 21807 20375
rect 21807 20341 21816 20375
rect 21764 20332 21816 20341
rect 22408 20332 22460 20384
rect 16796 20307 16848 20316
rect 16796 20273 16805 20307
rect 16805 20273 16839 20307
rect 16839 20273 16848 20307
rect 16796 20264 16848 20273
rect 17992 20264 18044 20316
rect 20108 20264 20160 20316
rect 22132 20264 22184 20316
rect 7320 20171 7372 20180
rect 7320 20137 7329 20171
rect 7329 20137 7363 20171
rect 7363 20137 7372 20171
rect 7320 20128 7372 20137
rect 13668 20171 13720 20180
rect 13668 20137 13677 20171
rect 13677 20137 13711 20171
rect 13711 20137 13720 20171
rect 13668 20128 13720 20137
rect 4652 20060 4704 20112
rect 5572 20060 5624 20112
rect 6216 20060 6268 20112
rect 6860 20060 6912 20112
rect 7872 20103 7924 20112
rect 7872 20069 7881 20103
rect 7881 20069 7915 20103
rect 7915 20069 7924 20103
rect 7872 20060 7924 20069
rect 20936 20060 20988 20112
rect 21672 20060 21724 20112
rect 22040 20103 22092 20112
rect 22040 20069 22049 20103
rect 22049 20069 22083 20103
rect 22083 20069 22092 20103
rect 22040 20060 22092 20069
rect 3510 19958 3562 20010
rect 3574 19958 3626 20010
rect 3638 19958 3690 20010
rect 3702 19958 3754 20010
rect 3766 19958 3818 20010
rect 880 19899 932 19908
rect 880 19865 889 19899
rect 889 19865 923 19899
rect 923 19865 932 19899
rect 880 19856 932 19865
rect 1248 19899 1300 19908
rect 1248 19865 1257 19899
rect 1257 19865 1291 19899
rect 1291 19865 1300 19899
rect 1248 19856 1300 19865
rect 2076 19899 2128 19908
rect 2076 19865 2085 19899
rect 2085 19865 2119 19899
rect 2119 19865 2128 19899
rect 2076 19856 2128 19865
rect 5480 19899 5532 19908
rect 788 19788 840 19840
rect 4376 19720 4428 19772
rect 5480 19865 5489 19899
rect 5489 19865 5523 19899
rect 5523 19865 5532 19899
rect 5480 19856 5532 19865
rect 6216 19899 6268 19908
rect 6216 19865 6225 19899
rect 6225 19865 6259 19899
rect 6259 19865 6268 19899
rect 6216 19856 6268 19865
rect 6400 19899 6452 19908
rect 6400 19865 6409 19899
rect 6409 19865 6443 19899
rect 6443 19865 6452 19899
rect 6400 19856 6452 19865
rect 7044 19856 7096 19908
rect 7320 19899 7372 19908
rect 7320 19865 7329 19899
rect 7329 19865 7363 19899
rect 7363 19865 7372 19899
rect 7320 19856 7372 19865
rect 9436 19856 9488 19908
rect 10264 19899 10316 19908
rect 10264 19865 10273 19899
rect 10273 19865 10307 19899
rect 10307 19865 10316 19899
rect 10264 19856 10316 19865
rect 13484 19899 13536 19908
rect 13484 19865 13493 19899
rect 13493 19865 13527 19899
rect 13527 19865 13536 19899
rect 13484 19856 13536 19865
rect 15416 19856 15468 19908
rect 16428 19856 16480 19908
rect 20660 19856 20712 19908
rect 20844 19856 20896 19908
rect 21764 19899 21816 19908
rect 21764 19865 21773 19899
rect 21773 19865 21807 19899
rect 21807 19865 21816 19899
rect 21764 19856 21816 19865
rect 22132 19899 22184 19908
rect 22132 19865 22141 19899
rect 22141 19865 22175 19899
rect 22175 19865 22184 19899
rect 22132 19856 22184 19865
rect 5020 19788 5072 19840
rect 5204 19720 5256 19772
rect 7872 19720 7924 19772
rect 8148 19763 8200 19772
rect 8148 19729 8157 19763
rect 8157 19729 8191 19763
rect 8191 19729 8200 19763
rect 8148 19720 8200 19729
rect 512 19516 564 19568
rect 1524 19516 1576 19568
rect 1708 19584 1760 19636
rect 5940 19652 5992 19704
rect 6860 19695 6912 19704
rect 6860 19661 6869 19695
rect 6869 19661 6903 19695
rect 6903 19661 6912 19695
rect 6860 19652 6912 19661
rect 8056 19652 8108 19704
rect 16796 19788 16848 19840
rect 16980 19788 17032 19840
rect 18084 19720 18136 19772
rect 5756 19627 5808 19636
rect 5756 19593 5765 19627
rect 5765 19593 5799 19627
rect 5799 19593 5808 19627
rect 5756 19584 5808 19593
rect 6584 19584 6636 19636
rect 18728 19652 18780 19704
rect 9344 19584 9396 19636
rect 20476 19720 20528 19772
rect 22040 19788 22092 19840
rect 23236 19720 23288 19772
rect 20292 19695 20344 19704
rect 20292 19661 20301 19695
rect 20301 19661 20335 19695
rect 20335 19661 20344 19695
rect 20292 19652 20344 19661
rect 20936 19695 20988 19704
rect 20936 19661 20945 19695
rect 20945 19661 20979 19695
rect 20979 19661 20988 19695
rect 20936 19652 20988 19661
rect 21856 19652 21908 19704
rect 19372 19584 19424 19636
rect 21672 19584 21724 19636
rect 2260 19516 2312 19568
rect 4192 19559 4244 19568
rect 4192 19525 4201 19559
rect 4201 19525 4235 19559
rect 4235 19525 4244 19559
rect 4192 19516 4244 19525
rect 4468 19516 4520 19568
rect 4652 19516 4704 19568
rect 5940 19559 5992 19568
rect 5940 19525 5949 19559
rect 5949 19525 5983 19559
rect 5983 19525 5992 19559
rect 5940 19516 5992 19525
rect 7136 19559 7188 19568
rect 7136 19525 7145 19559
rect 7145 19525 7179 19559
rect 7179 19525 7188 19559
rect 7136 19516 7188 19525
rect 13668 19559 13720 19568
rect 13668 19525 13677 19559
rect 13677 19525 13711 19559
rect 13711 19525 13720 19559
rect 13668 19516 13720 19525
rect 14128 19516 14180 19568
rect 18176 19559 18228 19568
rect 18176 19525 18185 19559
rect 18185 19525 18219 19559
rect 18219 19525 18228 19559
rect 18176 19516 18228 19525
rect 23236 19559 23288 19568
rect 23236 19525 23245 19559
rect 23245 19525 23279 19559
rect 23279 19525 23288 19559
rect 23236 19516 23288 19525
rect 23788 19516 23840 19568
rect 23972 19584 24024 19636
rect 25812 19627 25864 19636
rect 25812 19593 25821 19627
rect 25821 19593 25855 19627
rect 25855 19593 25864 19627
rect 25812 19584 25864 19593
rect 24984 19516 25036 19568
rect 18870 19414 18922 19466
rect 18934 19414 18986 19466
rect 18998 19414 19050 19466
rect 19062 19414 19114 19466
rect 19126 19414 19178 19466
rect 1340 19355 1392 19364
rect 1340 19321 1349 19355
rect 1349 19321 1383 19355
rect 1383 19321 1392 19355
rect 1340 19312 1392 19321
rect 1708 19312 1760 19364
rect 7688 19312 7740 19364
rect 20108 19312 20160 19364
rect 23144 19312 23196 19364
rect 23512 19312 23564 19364
rect 4560 19244 4612 19296
rect 6216 19244 6268 19296
rect 7044 19244 7096 19296
rect 22408 19244 22460 19296
rect 24064 19244 24116 19296
rect 4744 19176 4796 19228
rect 7596 19219 7648 19228
rect 7596 19185 7605 19219
rect 7605 19185 7639 19219
rect 7639 19185 7648 19219
rect 7596 19176 7648 19185
rect 9988 19176 10040 19228
rect 11092 19219 11144 19228
rect 11092 19185 11101 19219
rect 11101 19185 11135 19219
rect 11135 19185 11144 19219
rect 11092 19176 11144 19185
rect 11828 19176 11880 19228
rect 12932 19176 12984 19228
rect 13484 19219 13536 19228
rect 13484 19185 13493 19219
rect 13493 19185 13527 19219
rect 13527 19185 13536 19219
rect 13484 19176 13536 19185
rect 18544 19176 18596 19228
rect 18728 19219 18780 19228
rect 18728 19185 18737 19219
rect 18737 19185 18771 19219
rect 18771 19185 18780 19219
rect 18728 19176 18780 19185
rect 19372 19176 19424 19228
rect 22224 19219 22276 19228
rect 22224 19185 22233 19219
rect 22233 19185 22267 19219
rect 22267 19185 22276 19219
rect 22224 19176 22276 19185
rect 23328 19176 23380 19228
rect 26180 19244 26232 19296
rect 7504 19151 7556 19160
rect 7504 19117 7513 19151
rect 7513 19117 7547 19151
rect 7547 19117 7556 19151
rect 7504 19108 7556 19117
rect 8976 19108 9028 19160
rect 10172 19040 10224 19092
rect 10816 19108 10868 19160
rect 11000 19151 11052 19160
rect 11000 19117 11009 19151
rect 11009 19117 11043 19151
rect 11043 19117 11052 19151
rect 11000 19108 11052 19117
rect 12748 19151 12800 19160
rect 12748 19117 12757 19151
rect 12757 19117 12791 19151
rect 12791 19117 12800 19151
rect 13576 19151 13628 19160
rect 12748 19108 12800 19117
rect 13576 19117 13585 19151
rect 13585 19117 13619 19151
rect 13619 19117 13628 19151
rect 13576 19108 13628 19117
rect 18176 19151 18228 19160
rect 18176 19117 18185 19151
rect 18185 19117 18219 19151
rect 18219 19117 18228 19151
rect 18176 19108 18228 19117
rect 21396 19151 21448 19160
rect 21396 19117 21405 19151
rect 21405 19117 21439 19151
rect 21439 19117 21448 19151
rect 21396 19108 21448 19117
rect 21856 19108 21908 19160
rect 22408 19151 22460 19160
rect 22408 19117 22417 19151
rect 22417 19117 22451 19151
rect 22451 19117 22460 19151
rect 22408 19108 22460 19117
rect 16336 19040 16388 19092
rect 17900 19040 17952 19092
rect 19280 19040 19332 19092
rect 19924 19040 19976 19092
rect 5020 18972 5072 19024
rect 13852 19015 13904 19024
rect 13852 18981 13861 19015
rect 13861 18981 13895 19015
rect 13895 18981 13904 19015
rect 13852 18972 13904 18981
rect 17992 19015 18044 19024
rect 17992 18981 18001 19015
rect 18001 18981 18035 19015
rect 18035 18981 18044 19015
rect 17992 18972 18044 18981
rect 23236 19015 23288 19024
rect 23236 18981 23245 19015
rect 23245 18981 23279 19015
rect 23279 18981 23288 19015
rect 23236 18972 23288 18981
rect 23604 18972 23656 19024
rect 26088 19015 26140 19024
rect 26088 18981 26097 19015
rect 26097 18981 26131 19015
rect 26131 18981 26140 19015
rect 26088 18972 26140 18981
rect 3510 18870 3562 18922
rect 3574 18870 3626 18922
rect 3638 18870 3690 18922
rect 3702 18870 3754 18922
rect 3766 18870 3818 18922
rect 788 18768 840 18820
rect 1708 18768 1760 18820
rect 4560 18811 4612 18820
rect 4560 18777 4569 18811
rect 4569 18777 4603 18811
rect 4603 18777 4612 18811
rect 4560 18768 4612 18777
rect 7044 18768 7096 18820
rect 880 18632 932 18684
rect 4744 18700 4796 18752
rect 7504 18700 7556 18752
rect 8056 18743 8108 18752
rect 8056 18709 8065 18743
rect 8065 18709 8099 18743
rect 8099 18709 8108 18743
rect 8056 18700 8108 18709
rect 8332 18743 8384 18752
rect 8332 18709 8341 18743
rect 8341 18709 8375 18743
rect 8375 18709 8384 18743
rect 8332 18700 8384 18709
rect 1340 18607 1392 18616
rect 1340 18573 1349 18607
rect 1349 18573 1383 18607
rect 1383 18573 1392 18607
rect 1340 18564 1392 18573
rect 3364 18607 3416 18616
rect 512 18496 564 18548
rect 880 18471 932 18480
rect 880 18437 889 18471
rect 889 18437 923 18471
rect 923 18437 932 18471
rect 880 18428 932 18437
rect 1248 18496 1300 18548
rect 3364 18573 3373 18607
rect 3373 18573 3407 18607
rect 3407 18573 3416 18607
rect 3364 18564 3416 18573
rect 6308 18632 6360 18684
rect 7044 18632 7096 18684
rect 4468 18428 4520 18480
rect 4928 18471 4980 18480
rect 4928 18437 4937 18471
rect 4937 18437 4971 18471
rect 4971 18437 4980 18471
rect 4928 18428 4980 18437
rect 7504 18564 7556 18616
rect 5572 18496 5624 18548
rect 9160 18768 9212 18820
rect 11000 18768 11052 18820
rect 13576 18768 13628 18820
rect 18176 18768 18228 18820
rect 15784 18700 15836 18752
rect 17992 18700 18044 18752
rect 19280 18743 19332 18752
rect 19280 18709 19289 18743
rect 19289 18709 19323 18743
rect 19323 18709 19332 18743
rect 19280 18700 19332 18709
rect 9528 18632 9580 18684
rect 9068 18564 9120 18616
rect 12012 18564 12064 18616
rect 12748 18564 12800 18616
rect 13116 18564 13168 18616
rect 13852 18607 13904 18616
rect 13852 18573 13861 18607
rect 13861 18573 13895 18607
rect 13895 18573 13904 18607
rect 13852 18564 13904 18573
rect 15508 18564 15560 18616
rect 17900 18607 17952 18616
rect 17900 18573 17909 18607
rect 17909 18573 17943 18607
rect 17943 18573 17952 18607
rect 17900 18564 17952 18573
rect 18728 18632 18780 18684
rect 18084 18564 18136 18616
rect 18360 18607 18412 18616
rect 18360 18573 18369 18607
rect 18369 18573 18403 18607
rect 18403 18573 18412 18607
rect 18360 18564 18412 18573
rect 21396 18768 21448 18820
rect 22224 18768 22276 18820
rect 24156 18768 24208 18820
rect 24984 18811 25036 18820
rect 24984 18777 24993 18811
rect 24993 18777 25027 18811
rect 25027 18777 25036 18811
rect 24984 18768 25036 18777
rect 22408 18700 22460 18752
rect 21856 18675 21908 18684
rect 21856 18641 21865 18675
rect 21865 18641 21899 18675
rect 21899 18641 21908 18675
rect 21856 18632 21908 18641
rect 23420 18632 23472 18684
rect 23512 18675 23564 18684
rect 23512 18641 23521 18675
rect 23521 18641 23555 18675
rect 23555 18641 23564 18675
rect 23512 18632 23564 18641
rect 20108 18607 20160 18616
rect 20108 18573 20117 18607
rect 20117 18573 20151 18607
rect 20151 18573 20160 18607
rect 20108 18564 20160 18573
rect 20384 18607 20436 18616
rect 20384 18573 20393 18607
rect 20393 18573 20427 18607
rect 20427 18573 20436 18607
rect 20384 18564 20436 18573
rect 23604 18607 23656 18616
rect 11000 18496 11052 18548
rect 6308 18428 6360 18480
rect 9160 18428 9212 18480
rect 9988 18471 10040 18480
rect 9988 18437 9997 18471
rect 9997 18437 10031 18471
rect 10031 18437 10040 18471
rect 9988 18428 10040 18437
rect 10816 18428 10868 18480
rect 12196 18428 12248 18480
rect 13484 18496 13536 18548
rect 14128 18539 14180 18548
rect 14128 18505 14137 18539
rect 14137 18505 14171 18539
rect 14171 18505 14180 18539
rect 14128 18496 14180 18505
rect 15876 18539 15928 18548
rect 15876 18505 15885 18539
rect 15885 18505 15919 18539
rect 15919 18505 15928 18539
rect 15876 18496 15928 18505
rect 16244 18496 16296 18548
rect 22224 18496 22276 18548
rect 23604 18573 23613 18607
rect 23613 18573 23647 18607
rect 23647 18573 23656 18607
rect 23604 18564 23656 18573
rect 26180 18768 26232 18820
rect 23972 18607 24024 18616
rect 23972 18573 23981 18607
rect 23981 18573 24015 18607
rect 24015 18573 24024 18607
rect 23972 18564 24024 18573
rect 24156 18607 24208 18616
rect 24156 18573 24165 18607
rect 24165 18573 24199 18607
rect 24199 18573 24208 18607
rect 24156 18564 24208 18573
rect 25168 18607 25220 18616
rect 25168 18573 25177 18607
rect 25177 18573 25211 18607
rect 25211 18573 25220 18607
rect 25168 18564 25220 18573
rect 12932 18471 12984 18480
rect 12932 18437 12941 18471
rect 12941 18437 12975 18471
rect 12975 18437 12984 18471
rect 12932 18428 12984 18437
rect 18544 18428 18596 18480
rect 22408 18471 22460 18480
rect 22408 18437 22417 18471
rect 22417 18437 22451 18471
rect 22451 18437 22460 18471
rect 22408 18428 22460 18437
rect 24064 18428 24116 18480
rect 25996 18471 26048 18480
rect 25996 18437 26005 18471
rect 26005 18437 26039 18471
rect 26039 18437 26048 18471
rect 25996 18428 26048 18437
rect 26180 18471 26232 18480
rect 26180 18437 26189 18471
rect 26189 18437 26223 18471
rect 26223 18437 26232 18471
rect 26180 18428 26232 18437
rect 18870 18326 18922 18378
rect 18934 18326 18986 18378
rect 18998 18326 19050 18378
rect 19062 18326 19114 18378
rect 19126 18326 19178 18378
rect 3916 18224 3968 18276
rect 4928 18267 4980 18276
rect 4928 18233 4937 18267
rect 4937 18233 4971 18267
rect 4971 18233 4980 18267
rect 4928 18224 4980 18233
rect 6584 18267 6636 18276
rect 6584 18233 6593 18267
rect 6593 18233 6627 18267
rect 6627 18233 6636 18267
rect 6584 18224 6636 18233
rect 8056 18224 8108 18276
rect 10172 18267 10224 18276
rect 10172 18233 10181 18267
rect 10181 18233 10215 18267
rect 10215 18233 10224 18267
rect 10172 18224 10224 18233
rect 18176 18267 18228 18276
rect 18176 18233 18185 18267
rect 18185 18233 18219 18267
rect 18219 18233 18228 18267
rect 18176 18224 18228 18233
rect 13852 18156 13904 18208
rect 15784 18199 15836 18208
rect 15784 18165 15793 18199
rect 15793 18165 15827 18199
rect 15827 18165 15836 18199
rect 15784 18156 15836 18165
rect 16244 18156 16296 18208
rect 18728 18199 18780 18208
rect 18728 18165 18737 18199
rect 18737 18165 18771 18199
rect 18771 18165 18780 18199
rect 18728 18156 18780 18165
rect 4100 18131 4152 18140
rect 4100 18097 4109 18131
rect 4109 18097 4143 18131
rect 4143 18097 4152 18131
rect 4100 18088 4152 18097
rect 6308 18131 6360 18140
rect 6308 18097 6317 18131
rect 6317 18097 6351 18131
rect 6351 18097 6360 18131
rect 6308 18088 6360 18097
rect 4192 18020 4244 18072
rect 4928 18020 4980 18072
rect 6216 18020 6268 18072
rect 7412 18088 7464 18140
rect 9160 18088 9212 18140
rect 9436 18131 9488 18140
rect 9436 18097 9445 18131
rect 9445 18097 9479 18131
rect 9479 18097 9488 18131
rect 9436 18088 9488 18097
rect 11000 18131 11052 18140
rect 11000 18097 11009 18131
rect 11009 18097 11043 18131
rect 11043 18097 11052 18131
rect 11000 18088 11052 18097
rect 13116 18131 13168 18140
rect 13116 18097 13125 18131
rect 13125 18097 13159 18131
rect 13159 18097 13168 18131
rect 13116 18088 13168 18097
rect 18636 18131 18688 18140
rect 18636 18097 18645 18131
rect 18645 18097 18679 18131
rect 18679 18097 18688 18131
rect 20384 18224 20436 18276
rect 22408 18224 22460 18276
rect 23328 18267 23380 18276
rect 23328 18233 23337 18267
rect 23337 18233 23371 18267
rect 23371 18233 23380 18267
rect 23328 18224 23380 18233
rect 20292 18156 20344 18208
rect 23788 18199 23840 18208
rect 23788 18165 23797 18199
rect 23797 18165 23831 18199
rect 23831 18165 23840 18199
rect 23788 18156 23840 18165
rect 18636 18088 18688 18097
rect 20476 18088 20528 18140
rect 23420 18131 23472 18140
rect 23420 18097 23429 18131
rect 23429 18097 23463 18131
rect 23463 18097 23472 18131
rect 23420 18088 23472 18097
rect 6860 18020 6912 18072
rect 7504 18063 7556 18072
rect 7504 18029 7513 18063
rect 7513 18029 7547 18063
rect 7547 18029 7556 18063
rect 7504 18020 7556 18029
rect 8792 18020 8844 18072
rect 13668 18063 13720 18072
rect 13668 18029 13677 18063
rect 13677 18029 13711 18063
rect 13711 18029 13720 18063
rect 13668 18020 13720 18029
rect 12932 17952 12984 18004
rect 512 17884 564 17936
rect 788 17884 840 17936
rect 1064 17884 1116 17936
rect 1248 17927 1300 17936
rect 1248 17893 1257 17927
rect 1257 17893 1291 17927
rect 1291 17893 1300 17927
rect 1248 17884 1300 17893
rect 4192 17884 4244 17936
rect 4468 17884 4520 17936
rect 4560 17927 4612 17936
rect 4560 17893 4569 17927
rect 4569 17893 4603 17927
rect 4603 17893 4612 17927
rect 4560 17884 4612 17893
rect 5020 17884 5072 17936
rect 7596 17927 7648 17936
rect 7596 17893 7605 17927
rect 7605 17893 7639 17927
rect 7639 17893 7648 17927
rect 7596 17884 7648 17893
rect 9344 17884 9396 17936
rect 10816 17927 10868 17936
rect 10816 17893 10825 17927
rect 10825 17893 10859 17927
rect 10859 17893 10868 17927
rect 10816 17884 10868 17893
rect 14128 17884 14180 17936
rect 18084 18020 18136 18072
rect 20752 18063 20804 18072
rect 20752 18029 20761 18063
rect 20761 18029 20795 18063
rect 20795 18029 20804 18063
rect 20752 18020 20804 18029
rect 23236 18020 23288 18072
rect 15968 17884 16020 17936
rect 24432 17884 24484 17936
rect 3510 17782 3562 17834
rect 3574 17782 3626 17834
rect 3638 17782 3690 17834
rect 3702 17782 3754 17834
rect 3766 17782 3818 17834
rect 4928 17680 4980 17732
rect 5572 17723 5624 17732
rect 5572 17689 5581 17723
rect 5581 17689 5615 17723
rect 5615 17689 5624 17723
rect 5572 17680 5624 17689
rect 788 17587 840 17596
rect 788 17553 797 17587
rect 797 17553 831 17587
rect 831 17553 840 17587
rect 788 17544 840 17553
rect 972 17544 1024 17596
rect 3272 17544 3324 17596
rect 4468 17544 4520 17596
rect 512 17476 564 17528
rect 696 17408 748 17460
rect 4008 17476 4060 17528
rect 4744 17476 4796 17528
rect 6584 17680 6636 17732
rect 6860 17723 6912 17732
rect 6860 17689 6869 17723
rect 6869 17689 6903 17723
rect 6903 17689 6912 17723
rect 6860 17680 6912 17689
rect 7320 17680 7372 17732
rect 9804 17723 9856 17732
rect 9804 17689 9813 17723
rect 9813 17689 9847 17723
rect 9847 17689 9856 17723
rect 9804 17680 9856 17689
rect 13116 17723 13168 17732
rect 13116 17689 13125 17723
rect 13125 17689 13159 17723
rect 13159 17689 13168 17723
rect 13116 17680 13168 17689
rect 13852 17680 13904 17732
rect 15876 17680 15928 17732
rect 18728 17680 18780 17732
rect 20476 17680 20528 17732
rect 23420 17680 23472 17732
rect 23972 17680 24024 17732
rect 6400 17612 6452 17664
rect 13668 17612 13720 17664
rect 18636 17655 18688 17664
rect 18636 17621 18645 17655
rect 18645 17621 18679 17655
rect 18679 17621 18688 17655
rect 18636 17612 18688 17621
rect 4928 17476 4980 17528
rect 6400 17476 6452 17528
rect 7136 17476 7188 17528
rect 8056 17476 8108 17528
rect 5572 17408 5624 17460
rect 6124 17451 6176 17460
rect 6124 17417 6133 17451
rect 6133 17417 6167 17451
rect 6167 17417 6176 17451
rect 6124 17408 6176 17417
rect 6860 17408 6912 17460
rect 2628 17340 2680 17392
rect 4008 17383 4060 17392
rect 4008 17349 4017 17383
rect 4017 17349 4051 17383
rect 4051 17349 4060 17383
rect 4008 17340 4060 17349
rect 4376 17340 4428 17392
rect 7412 17340 7464 17392
rect 7964 17383 8016 17392
rect 7964 17349 7973 17383
rect 7973 17349 8007 17383
rect 8007 17349 8016 17383
rect 9252 17476 9304 17528
rect 15784 17544 15836 17596
rect 20292 17544 20344 17596
rect 9896 17476 9948 17528
rect 10816 17476 10868 17528
rect 14128 17519 14180 17528
rect 14128 17485 14137 17519
rect 14137 17485 14171 17519
rect 14171 17485 14180 17519
rect 14128 17476 14180 17485
rect 20752 17519 20804 17528
rect 20752 17485 20761 17519
rect 20761 17485 20795 17519
rect 20795 17485 20804 17519
rect 21120 17519 21172 17528
rect 20752 17476 20804 17485
rect 21120 17485 21129 17519
rect 21129 17485 21163 17519
rect 21163 17485 21172 17519
rect 21120 17476 21172 17485
rect 23512 17476 23564 17528
rect 9160 17451 9212 17460
rect 9160 17417 9169 17451
rect 9169 17417 9203 17451
rect 9203 17417 9212 17451
rect 9160 17408 9212 17417
rect 9988 17408 10040 17460
rect 13852 17408 13904 17460
rect 14588 17408 14640 17460
rect 21028 17451 21080 17460
rect 21028 17417 21037 17451
rect 21037 17417 21071 17451
rect 21071 17417 21080 17451
rect 24156 17612 24208 17664
rect 23696 17476 23748 17528
rect 24064 17476 24116 17528
rect 24432 17519 24484 17528
rect 24432 17485 24441 17519
rect 24441 17485 24475 17519
rect 24475 17485 24484 17519
rect 25812 17680 25864 17732
rect 24432 17476 24484 17485
rect 21028 17408 21080 17417
rect 7964 17340 8016 17349
rect 9436 17340 9488 17392
rect 11000 17340 11052 17392
rect 12196 17340 12248 17392
rect 15968 17383 16020 17392
rect 15968 17349 15977 17383
rect 15977 17349 16011 17383
rect 16011 17349 16020 17383
rect 15968 17340 16020 17349
rect 23788 17340 23840 17392
rect 18870 17238 18922 17290
rect 18934 17238 18986 17290
rect 18998 17238 19050 17290
rect 19062 17238 19114 17290
rect 19126 17238 19178 17290
rect 972 17179 1024 17188
rect 972 17145 981 17179
rect 981 17145 1015 17179
rect 1015 17145 1024 17179
rect 972 17136 1024 17145
rect 2628 17179 2680 17188
rect 2628 17145 2637 17179
rect 2637 17145 2671 17179
rect 2671 17145 2680 17179
rect 2628 17136 2680 17145
rect 4100 17136 4152 17188
rect 4560 17179 4612 17188
rect 4560 17145 4569 17179
rect 4569 17145 4603 17179
rect 4603 17145 4612 17179
rect 9344 17179 9396 17188
rect 4560 17136 4612 17145
rect 9344 17145 9353 17179
rect 9353 17145 9387 17179
rect 9387 17145 9396 17179
rect 9344 17136 9396 17145
rect 14588 17179 14640 17188
rect 14588 17145 14597 17179
rect 14597 17145 14631 17179
rect 14631 17145 14640 17179
rect 14588 17136 14640 17145
rect 1708 17111 1760 17120
rect 1708 17077 1717 17111
rect 1717 17077 1751 17111
rect 1751 17077 1760 17111
rect 1708 17068 1760 17077
rect 5756 17068 5808 17120
rect 5572 17000 5624 17052
rect 6124 17000 6176 17052
rect 6952 17000 7004 17052
rect 20476 17068 20528 17120
rect 10264 17000 10316 17052
rect 12196 17000 12248 17052
rect 15140 17000 15192 17052
rect 16428 17000 16480 17052
rect 20660 17000 20712 17052
rect 21488 17068 21540 17120
rect 21212 17043 21264 17052
rect 21212 17009 21221 17043
rect 21221 17009 21255 17043
rect 21255 17009 21264 17043
rect 21212 17000 21264 17009
rect 24340 17000 24392 17052
rect 26456 17000 26508 17052
rect 1248 16932 1300 16984
rect 4192 16932 4244 16984
rect 7964 16932 8016 16984
rect 9804 16932 9856 16984
rect 10908 16932 10960 16984
rect 12380 16975 12432 16984
rect 12380 16941 12389 16975
rect 12389 16941 12423 16975
rect 12423 16941 12432 16975
rect 12380 16932 12432 16941
rect 16704 16932 16756 16984
rect 21120 16932 21172 16984
rect 788 16864 840 16916
rect 2536 16864 2588 16916
rect 6216 16864 6268 16916
rect 6308 16864 6360 16916
rect 11552 16864 11604 16916
rect 23236 16864 23288 16916
rect 696 16839 748 16848
rect 696 16805 705 16839
rect 705 16805 739 16839
rect 739 16805 748 16839
rect 696 16796 748 16805
rect 1708 16796 1760 16848
rect 2628 16796 2680 16848
rect 5664 16796 5716 16848
rect 7228 16796 7280 16848
rect 8608 16796 8660 16848
rect 14680 16839 14732 16848
rect 14680 16805 14689 16839
rect 14689 16805 14723 16839
rect 14723 16805 14732 16839
rect 14680 16796 14732 16805
rect 15416 16839 15468 16848
rect 15416 16805 15425 16839
rect 15425 16805 15459 16839
rect 15459 16805 15468 16839
rect 15416 16796 15468 16805
rect 17808 16839 17860 16848
rect 17808 16805 17817 16839
rect 17817 16805 17851 16839
rect 17851 16805 17860 16839
rect 17808 16796 17860 16805
rect 20292 16839 20344 16848
rect 20292 16805 20301 16839
rect 20301 16805 20335 16839
rect 20335 16805 20344 16839
rect 20292 16796 20344 16805
rect 23144 16839 23196 16848
rect 23144 16805 23153 16839
rect 23153 16805 23187 16839
rect 23187 16805 23196 16839
rect 23144 16796 23196 16805
rect 24984 16839 25036 16848
rect 24984 16805 24993 16839
rect 24993 16805 25027 16839
rect 25027 16805 25036 16839
rect 24984 16796 25036 16805
rect 26364 16796 26416 16848
rect 3510 16694 3562 16746
rect 3574 16694 3626 16746
rect 3638 16694 3690 16746
rect 3702 16694 3754 16746
rect 3766 16694 3818 16746
rect 788 16592 840 16644
rect 1800 16635 1852 16644
rect 1800 16601 1809 16635
rect 1809 16601 1843 16635
rect 1843 16601 1852 16635
rect 1800 16592 1852 16601
rect 3272 16592 3324 16644
rect 4100 16592 4152 16644
rect 5572 16635 5624 16644
rect 5572 16601 5581 16635
rect 5581 16601 5615 16635
rect 5615 16601 5624 16635
rect 5572 16592 5624 16601
rect 5664 16592 5716 16644
rect 6952 16592 7004 16644
rect 8976 16592 9028 16644
rect 12380 16592 12432 16644
rect 14588 16635 14640 16644
rect 14588 16601 14597 16635
rect 14597 16601 14631 16635
rect 14631 16601 14640 16635
rect 14588 16592 14640 16601
rect 14680 16592 14732 16644
rect 15140 16635 15192 16644
rect 15140 16601 15149 16635
rect 15149 16601 15183 16635
rect 15183 16601 15192 16635
rect 15140 16592 15192 16601
rect 20476 16635 20528 16644
rect 20476 16601 20485 16635
rect 20485 16601 20519 16635
rect 20519 16601 20528 16635
rect 20476 16592 20528 16601
rect 20660 16635 20712 16644
rect 20660 16601 20669 16635
rect 20669 16601 20703 16635
rect 20703 16601 20712 16635
rect 20660 16592 20712 16601
rect 21120 16592 21172 16644
rect 24064 16592 24116 16644
rect 26456 16635 26508 16644
rect 3916 16567 3968 16576
rect 3916 16533 3925 16567
rect 3925 16533 3959 16567
rect 3959 16533 3968 16567
rect 3916 16524 3968 16533
rect 4284 16567 4336 16576
rect 4284 16533 4293 16567
rect 4293 16533 4327 16567
rect 4327 16533 4336 16567
rect 4284 16524 4336 16533
rect 2536 16499 2588 16508
rect 2536 16465 2542 16499
rect 2542 16465 2588 16499
rect 2536 16456 2588 16465
rect 3364 16456 3416 16508
rect 2628 16388 2680 16440
rect 3272 16388 3324 16440
rect 3916 16388 3968 16440
rect 5940 16524 5992 16576
rect 7228 16524 7280 16576
rect 9068 16499 9120 16508
rect 9068 16465 9077 16499
rect 9077 16465 9111 16499
rect 9111 16465 9120 16499
rect 9068 16456 9120 16465
rect 11184 16456 11236 16508
rect 15416 16499 15468 16508
rect 15416 16465 15425 16499
rect 15425 16465 15459 16499
rect 15459 16465 15468 16499
rect 15416 16456 15468 16465
rect 17808 16524 17860 16576
rect 21212 16524 21264 16576
rect 16428 16456 16480 16508
rect 23144 16524 23196 16576
rect 26456 16601 26465 16635
rect 26465 16601 26499 16635
rect 26499 16601 26508 16635
rect 26456 16592 26508 16601
rect 26364 16567 26416 16576
rect 5480 16388 5532 16440
rect 11828 16431 11880 16440
rect 11828 16397 11837 16431
rect 11837 16397 11871 16431
rect 11871 16397 11880 16431
rect 11828 16388 11880 16397
rect 13116 16388 13168 16440
rect 15140 16388 15192 16440
rect 17164 16388 17216 16440
rect 18544 16388 18596 16440
rect 23328 16456 23380 16508
rect 1248 16252 1300 16304
rect 1616 16252 1668 16304
rect 2996 16295 3048 16304
rect 2996 16261 3005 16295
rect 3005 16261 3039 16295
rect 3039 16261 3048 16295
rect 2996 16252 3048 16261
rect 5756 16295 5808 16304
rect 5756 16261 5765 16295
rect 5765 16261 5799 16295
rect 5799 16261 5808 16295
rect 5756 16252 5808 16261
rect 7228 16295 7280 16304
rect 7228 16261 7237 16295
rect 7237 16261 7271 16295
rect 7271 16261 7280 16295
rect 7228 16252 7280 16261
rect 8240 16295 8292 16304
rect 8240 16261 8249 16295
rect 8249 16261 8283 16295
rect 8283 16261 8292 16295
rect 8976 16320 9028 16372
rect 9344 16320 9396 16372
rect 11736 16320 11788 16372
rect 12104 16320 12156 16372
rect 15324 16320 15376 16372
rect 19280 16388 19332 16440
rect 23236 16388 23288 16440
rect 23788 16456 23840 16508
rect 24984 16499 25036 16508
rect 24984 16465 24993 16499
rect 24993 16465 25027 16499
rect 25027 16465 25036 16499
rect 24984 16456 25036 16465
rect 25812 16456 25864 16508
rect 26364 16533 26373 16567
rect 26373 16533 26407 16567
rect 26407 16533 26416 16567
rect 26364 16524 26416 16533
rect 23696 16320 23748 16372
rect 24064 16431 24116 16440
rect 24064 16397 24073 16431
rect 24073 16397 24107 16431
rect 24107 16397 24116 16431
rect 24064 16388 24116 16397
rect 24248 16388 24300 16440
rect 8240 16252 8292 16261
rect 8608 16295 8660 16304
rect 8608 16261 8617 16295
rect 8617 16261 8651 16295
rect 8651 16261 8660 16295
rect 8608 16252 8660 16261
rect 10264 16252 10316 16304
rect 10908 16295 10960 16304
rect 10908 16261 10917 16295
rect 10917 16261 10951 16295
rect 10951 16261 10960 16295
rect 10908 16252 10960 16261
rect 11184 16295 11236 16304
rect 11184 16261 11193 16295
rect 11193 16261 11227 16295
rect 11227 16261 11236 16295
rect 11184 16252 11236 16261
rect 11460 16295 11512 16304
rect 11460 16261 11469 16295
rect 11469 16261 11503 16295
rect 11503 16261 11512 16295
rect 11460 16252 11512 16261
rect 16704 16295 16756 16304
rect 16704 16261 16713 16295
rect 16713 16261 16747 16295
rect 16747 16261 16756 16295
rect 16704 16252 16756 16261
rect 19372 16252 19424 16304
rect 20292 16252 20344 16304
rect 21488 16295 21540 16304
rect 21488 16261 21497 16295
rect 21497 16261 21531 16295
rect 21531 16261 21540 16295
rect 21488 16252 21540 16261
rect 25812 16320 25864 16372
rect 26272 16320 26324 16372
rect 24708 16295 24760 16304
rect 24708 16261 24717 16295
rect 24717 16261 24751 16295
rect 24751 16261 24760 16295
rect 24708 16252 24760 16261
rect 18870 16150 18922 16202
rect 18934 16150 18986 16202
rect 18998 16150 19050 16202
rect 19062 16150 19114 16202
rect 19126 16150 19178 16202
rect 1708 16091 1760 16100
rect 1708 16057 1717 16091
rect 1717 16057 1751 16091
rect 1751 16057 1760 16091
rect 1708 16048 1760 16057
rect 4284 16048 4336 16100
rect 9068 16048 9120 16100
rect 9344 16048 9396 16100
rect 12104 16091 12156 16100
rect 12104 16057 12113 16091
rect 12113 16057 12147 16091
rect 12147 16057 12156 16091
rect 12104 16048 12156 16057
rect 16428 16048 16480 16100
rect 17900 16048 17952 16100
rect 1800 15980 1852 16032
rect 5480 15980 5532 16032
rect 6216 16023 6268 16032
rect 6216 15989 6225 16023
rect 6225 15989 6259 16023
rect 6259 15989 6268 16023
rect 6216 15980 6268 15989
rect 6584 16023 6636 16032
rect 6584 15989 6593 16023
rect 6593 15989 6627 16023
rect 6627 15989 6636 16023
rect 6584 15980 6636 15989
rect 9528 16023 9580 16032
rect 9528 15989 9537 16023
rect 9537 15989 9571 16023
rect 9571 15989 9580 16023
rect 9528 15980 9580 15989
rect 11460 15980 11512 16032
rect 12196 15980 12248 16032
rect 13116 15980 13168 16032
rect 20660 15980 20712 16032
rect 1800 15844 1852 15896
rect 5940 15912 5992 15964
rect 8608 15912 8660 15964
rect 9712 15912 9764 15964
rect 11368 15955 11420 15964
rect 11368 15921 11377 15955
rect 11377 15921 11411 15955
rect 11411 15921 11420 15955
rect 11368 15912 11420 15921
rect 16612 15955 16664 15964
rect 16612 15921 16621 15955
rect 16621 15921 16655 15955
rect 16655 15921 16664 15955
rect 16612 15912 16664 15921
rect 16980 15955 17032 15964
rect 16980 15921 16989 15955
rect 16989 15921 17023 15955
rect 17023 15921 17032 15955
rect 16980 15912 17032 15921
rect 17072 15912 17124 15964
rect 17808 15912 17860 15964
rect 21028 15955 21080 15964
rect 21028 15921 21037 15955
rect 21037 15921 21071 15955
rect 21071 15921 21080 15955
rect 21028 15912 21080 15921
rect 25720 16048 25772 16100
rect 23420 15980 23472 16032
rect 22684 15912 22736 15964
rect 25812 15955 25864 15964
rect 25812 15921 25821 15955
rect 25821 15921 25855 15955
rect 25855 15921 25864 15955
rect 25812 15912 25864 15921
rect 4928 15844 4980 15896
rect 5848 15887 5900 15896
rect 5848 15853 5857 15887
rect 5857 15853 5891 15887
rect 5891 15853 5900 15887
rect 5848 15844 5900 15853
rect 6676 15844 6728 15896
rect 8240 15844 8292 15896
rect 9160 15887 9212 15896
rect 9160 15853 9169 15887
rect 9169 15853 9203 15887
rect 9203 15853 9212 15887
rect 9160 15844 9212 15853
rect 9804 15844 9856 15896
rect 9988 15844 10040 15896
rect 13392 15844 13444 15896
rect 13668 15887 13720 15896
rect 13668 15853 13677 15887
rect 13677 15853 13711 15887
rect 13711 15853 13720 15887
rect 13668 15844 13720 15853
rect 14680 15844 14732 15896
rect 15232 15844 15284 15896
rect 16704 15844 16756 15896
rect 20200 15887 20252 15896
rect 20200 15853 20209 15887
rect 20209 15853 20243 15887
rect 20243 15853 20252 15887
rect 20200 15844 20252 15853
rect 2076 15776 2128 15828
rect 2996 15776 3048 15828
rect 9620 15776 9672 15828
rect 11828 15776 11880 15828
rect 13576 15819 13628 15828
rect 13576 15785 13585 15819
rect 13585 15785 13619 15819
rect 13619 15785 13628 15819
rect 13576 15776 13628 15785
rect 20292 15776 20344 15828
rect 24248 15844 24300 15896
rect 24708 15844 24760 15896
rect 21488 15776 21540 15828
rect 24064 15819 24116 15828
rect 24064 15785 24073 15819
rect 24073 15785 24107 15819
rect 24107 15785 24116 15819
rect 24064 15776 24116 15785
rect 2168 15751 2220 15760
rect 2168 15717 2177 15751
rect 2177 15717 2211 15751
rect 2211 15717 2220 15751
rect 2168 15708 2220 15717
rect 6308 15708 6360 15760
rect 7780 15751 7832 15760
rect 7780 15717 7789 15751
rect 7789 15717 7823 15751
rect 7823 15717 7832 15751
rect 7780 15708 7832 15717
rect 11552 15751 11604 15760
rect 11552 15717 11561 15751
rect 11561 15717 11595 15751
rect 11595 15717 11604 15751
rect 11552 15708 11604 15717
rect 15324 15751 15376 15760
rect 15324 15717 15333 15751
rect 15333 15717 15367 15751
rect 15367 15717 15376 15751
rect 15324 15708 15376 15717
rect 16888 15708 16940 15760
rect 23236 15708 23288 15760
rect 26272 15708 26324 15760
rect 3510 15606 3562 15658
rect 3574 15606 3626 15658
rect 3638 15606 3690 15658
rect 3702 15606 3754 15658
rect 3766 15606 3818 15658
rect 1800 15547 1852 15556
rect 1800 15513 1809 15547
rect 1809 15513 1843 15547
rect 1843 15513 1852 15547
rect 1800 15504 1852 15513
rect 1892 15547 1944 15556
rect 1892 15513 1901 15547
rect 1901 15513 1935 15547
rect 1935 15513 1944 15547
rect 1892 15504 1944 15513
rect 2444 15504 2496 15556
rect 2996 15547 3048 15556
rect 2996 15513 3005 15547
rect 3005 15513 3039 15547
rect 3039 15513 3048 15547
rect 2996 15504 3048 15513
rect 3916 15504 3968 15556
rect 4008 15504 4060 15556
rect 1708 15436 1760 15488
rect 9620 15504 9672 15556
rect 9804 15547 9856 15556
rect 9804 15513 9813 15547
rect 9813 15513 9847 15547
rect 9847 15513 9856 15547
rect 9804 15504 9856 15513
rect 11368 15547 11420 15556
rect 11368 15513 11377 15547
rect 11377 15513 11411 15547
rect 11411 15513 11420 15547
rect 11368 15504 11420 15513
rect 11552 15547 11604 15556
rect 11552 15513 11561 15547
rect 11561 15513 11595 15547
rect 11595 15513 11604 15547
rect 11552 15504 11604 15513
rect 15232 15547 15284 15556
rect 15232 15513 15241 15547
rect 15241 15513 15275 15547
rect 15275 15513 15284 15547
rect 15232 15504 15284 15513
rect 15416 15504 15468 15556
rect 15876 15504 15928 15556
rect 16888 15547 16940 15556
rect 16888 15513 16897 15547
rect 16897 15513 16931 15547
rect 16931 15513 16940 15547
rect 16888 15504 16940 15513
rect 20292 15547 20344 15556
rect 20292 15513 20301 15547
rect 20301 15513 20335 15547
rect 20335 15513 20344 15547
rect 20292 15504 20344 15513
rect 21028 15504 21080 15556
rect 24064 15547 24116 15556
rect 24064 15513 24073 15547
rect 24073 15513 24107 15547
rect 24107 15513 24116 15547
rect 24064 15504 24116 15513
rect 26272 15547 26324 15556
rect 26272 15513 26281 15547
rect 26281 15513 26315 15547
rect 26315 15513 26324 15547
rect 26272 15504 26324 15513
rect 6952 15436 7004 15488
rect 7780 15436 7832 15488
rect 7964 15479 8016 15488
rect 7964 15445 7973 15479
rect 7973 15445 8007 15479
rect 8007 15445 8016 15479
rect 7964 15436 8016 15445
rect 1892 15368 1944 15420
rect 2628 15368 2680 15420
rect 3272 15368 3324 15420
rect 880 15343 932 15352
rect 880 15309 889 15343
rect 889 15309 923 15343
rect 923 15309 932 15343
rect 880 15300 932 15309
rect 1984 15300 2036 15352
rect 5572 15368 5624 15420
rect 5848 15368 5900 15420
rect 6676 15368 6728 15420
rect 6860 15411 6912 15420
rect 6860 15377 6869 15411
rect 6869 15377 6903 15411
rect 6903 15377 6912 15411
rect 6860 15368 6912 15377
rect 7136 15368 7188 15420
rect 8056 15411 8108 15420
rect 8056 15377 8065 15411
rect 8065 15377 8099 15411
rect 8099 15377 8108 15411
rect 8056 15368 8108 15377
rect 1708 15232 1760 15284
rect 5112 15300 5164 15352
rect 9344 15436 9396 15488
rect 9528 15479 9580 15488
rect 9528 15445 9537 15479
rect 9537 15445 9571 15479
rect 9571 15445 9580 15479
rect 9528 15436 9580 15445
rect 13576 15436 13628 15488
rect 15784 15479 15836 15488
rect 15784 15445 15793 15479
rect 15793 15445 15827 15479
rect 15827 15445 15836 15479
rect 15784 15436 15836 15445
rect 17072 15436 17124 15488
rect 20200 15436 20252 15488
rect 13392 15300 13444 15352
rect 14128 15368 14180 15420
rect 15324 15368 15376 15420
rect 16612 15368 16664 15420
rect 20660 15368 20712 15420
rect 25812 15368 25864 15420
rect 5480 15207 5532 15216
rect 5480 15173 5489 15207
rect 5489 15173 5523 15207
rect 5523 15173 5532 15207
rect 5480 15164 5532 15173
rect 6308 15207 6360 15216
rect 6308 15173 6317 15207
rect 6317 15173 6351 15207
rect 6351 15173 6360 15207
rect 6308 15164 6360 15173
rect 6400 15164 6452 15216
rect 7872 15232 7924 15284
rect 16980 15300 17032 15352
rect 22776 15300 22828 15352
rect 23788 15300 23840 15352
rect 15784 15232 15836 15284
rect 24340 15232 24392 15284
rect 24892 15232 24944 15284
rect 7320 15207 7372 15216
rect 7320 15173 7329 15207
rect 7329 15173 7363 15207
rect 7363 15173 7372 15207
rect 7320 15164 7372 15173
rect 9160 15164 9212 15216
rect 9712 15164 9764 15216
rect 12656 15207 12708 15216
rect 12656 15173 12665 15207
rect 12665 15173 12699 15207
rect 12699 15173 12708 15207
rect 12656 15164 12708 15173
rect 13392 15164 13444 15216
rect 22684 15207 22736 15216
rect 22684 15173 22693 15207
rect 22693 15173 22727 15207
rect 22727 15173 22736 15207
rect 22684 15164 22736 15173
rect 23236 15207 23288 15216
rect 23236 15173 23245 15207
rect 23245 15173 23279 15207
rect 23279 15173 23288 15207
rect 23236 15164 23288 15173
rect 24248 15164 24300 15216
rect 18870 15062 18922 15114
rect 18934 15062 18986 15114
rect 18998 15062 19050 15114
rect 19062 15062 19114 15114
rect 19126 15062 19178 15114
rect 1984 15003 2036 15012
rect 1984 14969 1993 15003
rect 1993 14969 2027 15003
rect 2027 14969 2036 15003
rect 1984 14960 2036 14969
rect 2168 14960 2220 15012
rect 4560 14960 4612 15012
rect 5388 14960 5440 15012
rect 5940 15003 5992 15012
rect 5940 14969 5949 15003
rect 5949 14969 5983 15003
rect 5983 14969 5992 15003
rect 5940 14960 5992 14969
rect 6216 14960 6268 15012
rect 6676 15003 6728 15012
rect 6676 14969 6685 15003
rect 6685 14969 6719 15003
rect 6719 14969 6728 15003
rect 6676 14960 6728 14969
rect 8700 14960 8752 15012
rect 9620 14960 9672 15012
rect 12012 15003 12064 15012
rect 12012 14969 12021 15003
rect 12021 14969 12055 15003
rect 12055 14969 12064 15003
rect 12012 14960 12064 14969
rect 13668 14960 13720 15012
rect 15876 15003 15928 15012
rect 15876 14969 15885 15003
rect 15885 14969 15919 15003
rect 15919 14969 15928 15003
rect 15876 14960 15928 14969
rect 23696 15003 23748 15012
rect 23696 14969 23705 15003
rect 23705 14969 23739 15003
rect 23739 14969 23748 15003
rect 23696 14960 23748 14969
rect 24892 14960 24944 15012
rect 1892 14892 1944 14944
rect 2536 14892 2588 14944
rect 2720 14892 2772 14944
rect 4376 14892 4428 14944
rect 5112 14892 5164 14944
rect 2628 14824 2680 14876
rect 2812 14824 2864 14876
rect 3456 14867 3508 14876
rect 3456 14833 3465 14867
rect 3465 14833 3499 14867
rect 3499 14833 3508 14867
rect 3456 14824 3508 14833
rect 5020 14824 5072 14876
rect 5296 14867 5348 14876
rect 5296 14833 5305 14867
rect 5305 14833 5339 14867
rect 5339 14833 5348 14867
rect 5296 14824 5348 14833
rect 5848 14892 5900 14944
rect 6584 14935 6636 14944
rect 6584 14901 6593 14935
rect 6593 14901 6627 14935
rect 6627 14901 6636 14935
rect 6584 14892 6636 14901
rect 12656 14892 12708 14944
rect 13576 14892 13628 14944
rect 16888 14892 16940 14944
rect 23420 14892 23472 14944
rect 24064 14892 24116 14944
rect 24340 14935 24392 14944
rect 24340 14901 24349 14935
rect 24349 14901 24383 14935
rect 24383 14901 24392 14935
rect 24340 14892 24392 14901
rect 25812 14892 25864 14944
rect 3272 14756 3324 14808
rect 6124 14824 6176 14876
rect 6860 14824 6912 14876
rect 8424 14824 8476 14876
rect 8976 14867 9028 14876
rect 8976 14833 8985 14867
rect 8985 14833 9019 14867
rect 9019 14833 9028 14867
rect 8976 14824 9028 14833
rect 9068 14824 9120 14876
rect 11644 14824 11696 14876
rect 16428 14824 16480 14876
rect 17164 14867 17216 14876
rect 17164 14833 17173 14867
rect 17173 14833 17207 14867
rect 17207 14833 17216 14867
rect 17164 14824 17216 14833
rect 17992 14867 18044 14876
rect 17992 14833 18001 14867
rect 18001 14833 18035 14867
rect 18035 14833 18044 14867
rect 17992 14824 18044 14833
rect 22776 14867 22828 14876
rect 22776 14833 22785 14867
rect 22785 14833 22819 14867
rect 22819 14833 22828 14867
rect 22776 14824 22828 14833
rect 23052 14824 23104 14876
rect 23328 14867 23380 14876
rect 23328 14833 23337 14867
rect 23337 14833 23371 14867
rect 23371 14833 23380 14867
rect 23328 14824 23380 14833
rect 23696 14824 23748 14876
rect 5756 14756 5808 14808
rect 6952 14756 7004 14808
rect 7412 14756 7464 14808
rect 8516 14756 8568 14808
rect 9344 14756 9396 14808
rect 10724 14756 10776 14808
rect 12196 14756 12248 14808
rect 16152 14799 16204 14808
rect 16152 14765 16161 14799
rect 16161 14765 16195 14799
rect 16195 14765 16204 14799
rect 16152 14756 16204 14765
rect 16612 14756 16664 14808
rect 22316 14799 22368 14808
rect 22316 14765 22325 14799
rect 22325 14765 22359 14799
rect 22359 14765 22368 14799
rect 22316 14756 22368 14765
rect 23236 14799 23288 14808
rect 23236 14765 23245 14799
rect 23245 14765 23279 14799
rect 23279 14765 23288 14799
rect 23236 14756 23288 14765
rect 4100 14688 4152 14740
rect 5204 14688 5256 14740
rect 6492 14688 6544 14740
rect 6768 14688 6820 14740
rect 11552 14731 11604 14740
rect 11552 14697 11576 14731
rect 11576 14697 11604 14731
rect 11552 14688 11604 14697
rect 12932 14688 12984 14740
rect 2444 14620 2496 14672
rect 3088 14620 3140 14672
rect 5848 14620 5900 14672
rect 6400 14620 6452 14672
rect 6860 14620 6912 14672
rect 7228 14620 7280 14672
rect 7780 14620 7832 14672
rect 8608 14620 8660 14672
rect 8792 14620 8844 14672
rect 9344 14620 9396 14672
rect 9436 14620 9488 14672
rect 9804 14620 9856 14672
rect 10632 14620 10684 14672
rect 11736 14620 11788 14672
rect 17440 14620 17492 14672
rect 18728 14620 18780 14672
rect 20476 14620 20528 14672
rect 3510 14518 3562 14570
rect 3574 14518 3626 14570
rect 3638 14518 3690 14570
rect 3702 14518 3754 14570
rect 3766 14518 3818 14570
rect 3088 14459 3140 14468
rect 3088 14425 3097 14459
rect 3097 14425 3131 14459
rect 3131 14425 3140 14459
rect 3088 14416 3140 14425
rect 3364 14416 3416 14468
rect 1156 14348 1208 14400
rect 1800 14348 1852 14400
rect 4192 14391 4244 14400
rect 4192 14357 4201 14391
rect 4201 14357 4235 14391
rect 4235 14357 4244 14391
rect 4192 14348 4244 14357
rect 4560 14459 4612 14468
rect 4560 14425 4569 14459
rect 4569 14425 4603 14459
rect 4603 14425 4612 14459
rect 4560 14416 4612 14425
rect 5020 14416 5072 14468
rect 6492 14459 6544 14468
rect 6492 14425 6501 14459
rect 6501 14425 6535 14459
rect 6535 14425 6544 14459
rect 6492 14416 6544 14425
rect 6860 14416 6912 14468
rect 6952 14459 7004 14468
rect 6952 14425 6961 14459
rect 6961 14425 6995 14459
rect 6995 14425 7004 14459
rect 8424 14459 8476 14468
rect 6952 14416 7004 14425
rect 8424 14425 8433 14459
rect 8433 14425 8467 14459
rect 8467 14425 8476 14459
rect 8424 14416 8476 14425
rect 8608 14459 8660 14468
rect 8608 14425 8617 14459
rect 8617 14425 8651 14459
rect 8651 14425 8660 14459
rect 8608 14416 8660 14425
rect 8976 14416 9028 14468
rect 9344 14459 9396 14468
rect 9344 14425 9353 14459
rect 9353 14425 9387 14459
rect 9387 14425 9396 14459
rect 9344 14416 9396 14425
rect 9528 14459 9580 14468
rect 9528 14425 9537 14459
rect 9537 14425 9571 14459
rect 9571 14425 9580 14459
rect 9528 14416 9580 14425
rect 9988 14416 10040 14468
rect 10724 14459 10776 14468
rect 10724 14425 10733 14459
rect 10733 14425 10767 14459
rect 10767 14425 10776 14459
rect 10724 14416 10776 14425
rect 11368 14416 11420 14468
rect 12104 14416 12156 14468
rect 12932 14459 12984 14468
rect 12932 14425 12941 14459
rect 12941 14425 12975 14459
rect 12975 14425 12984 14459
rect 12932 14416 12984 14425
rect 13576 14416 13628 14468
rect 16152 14416 16204 14468
rect 17440 14459 17492 14468
rect 6584 14348 6636 14400
rect 7504 14391 7556 14400
rect 7504 14357 7513 14391
rect 7513 14357 7547 14391
rect 7547 14357 7556 14391
rect 7504 14348 7556 14357
rect 2720 14280 2772 14332
rect 4376 14280 4428 14332
rect 5112 14323 5164 14332
rect 5112 14289 5121 14323
rect 5121 14289 5155 14323
rect 5155 14289 5164 14323
rect 5112 14280 5164 14289
rect 1340 14076 1392 14128
rect 1800 14212 1852 14264
rect 1984 14187 2036 14196
rect 1984 14153 1993 14187
rect 1993 14153 2027 14187
rect 2027 14153 2036 14187
rect 1984 14144 2036 14153
rect 3088 14212 3140 14264
rect 5756 14255 5808 14264
rect 5756 14221 5765 14255
rect 5765 14221 5799 14255
rect 5799 14221 5808 14255
rect 5756 14212 5808 14221
rect 2996 14076 3048 14128
rect 3272 14119 3324 14128
rect 3272 14085 3281 14119
rect 3281 14085 3315 14119
rect 3315 14085 3324 14119
rect 3272 14076 3324 14085
rect 3364 14119 3416 14128
rect 3364 14085 3373 14119
rect 3373 14085 3407 14119
rect 3407 14085 3416 14119
rect 5388 14119 5440 14128
rect 3364 14076 3416 14085
rect 5388 14085 5397 14119
rect 5397 14085 5431 14119
rect 5431 14085 5440 14119
rect 5388 14076 5440 14085
rect 5756 14076 5808 14128
rect 6124 14076 6176 14128
rect 6216 14076 6268 14128
rect 8056 14280 8108 14332
rect 9068 14391 9120 14400
rect 9068 14357 9077 14391
rect 9077 14357 9111 14391
rect 9111 14357 9120 14391
rect 9068 14348 9120 14357
rect 10080 14348 10132 14400
rect 10172 14348 10224 14400
rect 11552 14348 11604 14400
rect 12012 14391 12064 14400
rect 12012 14357 12021 14391
rect 12021 14357 12055 14391
rect 12055 14357 12064 14391
rect 12012 14348 12064 14357
rect 16428 14391 16480 14400
rect 16428 14357 16437 14391
rect 16437 14357 16471 14391
rect 16471 14357 16480 14391
rect 16428 14348 16480 14357
rect 16612 14391 16664 14400
rect 16612 14357 16621 14391
rect 16621 14357 16655 14391
rect 16655 14357 16664 14391
rect 16612 14348 16664 14357
rect 11276 14280 11328 14332
rect 11460 14280 11512 14332
rect 7136 14255 7188 14264
rect 7136 14221 7145 14255
rect 7145 14221 7179 14255
rect 7179 14221 7188 14255
rect 7136 14212 7188 14221
rect 9528 14212 9580 14264
rect 9988 14212 10040 14264
rect 10448 14212 10500 14264
rect 10724 14212 10776 14264
rect 10908 14212 10960 14264
rect 11552 14212 11604 14264
rect 13576 14255 13628 14264
rect 13576 14221 13585 14255
rect 13585 14221 13619 14255
rect 13619 14221 13628 14255
rect 13576 14212 13628 14221
rect 17440 14425 17449 14459
rect 17449 14425 17483 14459
rect 17483 14425 17492 14459
rect 17440 14416 17492 14425
rect 23236 14416 23288 14468
rect 20200 14348 20252 14400
rect 20568 14391 20620 14400
rect 20568 14357 20577 14391
rect 20577 14357 20611 14391
rect 20611 14357 20620 14391
rect 20568 14348 20620 14357
rect 23328 14348 23380 14400
rect 18452 14323 18504 14332
rect 18452 14289 18461 14323
rect 18461 14289 18495 14323
rect 18495 14289 18504 14323
rect 18452 14280 18504 14289
rect 19924 14323 19976 14332
rect 19924 14289 19933 14323
rect 19933 14289 19967 14323
rect 19967 14289 19976 14323
rect 19924 14280 19976 14289
rect 18728 14255 18780 14264
rect 18728 14221 18737 14255
rect 18737 14221 18771 14255
rect 18771 14221 18780 14255
rect 18728 14212 18780 14221
rect 19280 14212 19332 14264
rect 21672 14280 21724 14332
rect 23420 14280 23472 14332
rect 23604 14280 23656 14332
rect 20476 14212 20528 14264
rect 22776 14212 22828 14264
rect 23788 14255 23840 14264
rect 23788 14221 23797 14255
rect 23797 14221 23831 14255
rect 23831 14221 23840 14255
rect 23788 14212 23840 14221
rect 24892 14280 24944 14332
rect 24432 14212 24484 14264
rect 25996 14255 26048 14264
rect 25996 14221 26005 14255
rect 26005 14221 26039 14255
rect 26039 14221 26048 14255
rect 25996 14212 26048 14221
rect 7688 14144 7740 14196
rect 10356 14144 10408 14196
rect 11736 14187 11788 14196
rect 11736 14153 11745 14187
rect 11745 14153 11779 14187
rect 11779 14153 11788 14187
rect 11736 14144 11788 14153
rect 12840 14187 12892 14196
rect 12840 14153 12849 14187
rect 12849 14153 12883 14187
rect 12883 14153 12892 14187
rect 12840 14144 12892 14153
rect 17164 14144 17216 14196
rect 8056 14119 8108 14128
rect 8056 14085 8065 14119
rect 8065 14085 8099 14119
rect 8099 14085 8108 14119
rect 8056 14076 8108 14085
rect 9344 14076 9396 14128
rect 11828 14076 11880 14128
rect 14036 14119 14088 14128
rect 14036 14085 14045 14119
rect 14045 14085 14079 14119
rect 14079 14085 14088 14119
rect 14036 14076 14088 14085
rect 17808 14144 17860 14196
rect 18452 14076 18504 14128
rect 23052 14076 23104 14128
rect 18870 13974 18922 14026
rect 18934 13974 18986 14026
rect 18998 13974 19050 14026
rect 19062 13974 19114 14026
rect 19126 13974 19178 14026
rect 4284 13915 4336 13924
rect 4284 13881 4293 13915
rect 4293 13881 4327 13915
rect 4327 13881 4336 13915
rect 4284 13872 4336 13881
rect 4376 13872 4428 13924
rect 6308 13872 6360 13924
rect 9712 13872 9764 13924
rect 10080 13872 10132 13924
rect 12104 13915 12156 13924
rect 12104 13881 12113 13915
rect 12113 13881 12147 13915
rect 12147 13881 12156 13915
rect 12104 13872 12156 13881
rect 17992 13915 18044 13924
rect 17992 13881 18001 13915
rect 18001 13881 18035 13915
rect 18035 13881 18044 13915
rect 17992 13872 18044 13881
rect 18544 13872 18596 13924
rect 19372 13872 19424 13924
rect 4008 13847 4060 13856
rect 4008 13813 4017 13847
rect 4017 13813 4051 13847
rect 4051 13813 4060 13847
rect 4008 13804 4060 13813
rect 5664 13804 5716 13856
rect 7412 13804 7464 13856
rect 8056 13804 8108 13856
rect 9988 13847 10040 13856
rect 9988 13813 9997 13847
rect 9997 13813 10031 13847
rect 10031 13813 10040 13847
rect 9988 13804 10040 13813
rect 10356 13804 10408 13856
rect 10540 13847 10592 13856
rect 10540 13813 10549 13847
rect 10549 13813 10583 13847
rect 10583 13813 10592 13847
rect 10540 13804 10592 13813
rect 1708 13736 1760 13788
rect 2260 13736 2312 13788
rect 4100 13736 4152 13788
rect 6860 13736 6912 13788
rect 10080 13779 10132 13788
rect 10080 13745 10089 13779
rect 10089 13745 10123 13779
rect 10123 13745 10132 13779
rect 10080 13736 10132 13745
rect 10448 13736 10500 13788
rect 11276 13736 11328 13788
rect 18544 13779 18596 13788
rect 3088 13668 3140 13720
rect 5848 13668 5900 13720
rect 4192 13600 4244 13652
rect 7964 13668 8016 13720
rect 9528 13668 9580 13720
rect 9988 13668 10040 13720
rect 12012 13668 12064 13720
rect 13944 13668 13996 13720
rect 18544 13745 18553 13779
rect 18553 13745 18587 13779
rect 18587 13745 18596 13779
rect 18544 13736 18596 13745
rect 18820 13736 18872 13788
rect 15968 13668 16020 13720
rect 18452 13668 18504 13720
rect 8608 13600 8660 13652
rect 9160 13600 9212 13652
rect 1340 13532 1392 13584
rect 6124 13575 6176 13584
rect 6124 13541 6133 13575
rect 6133 13541 6167 13575
rect 6167 13541 6176 13575
rect 6124 13532 6176 13541
rect 7136 13532 7188 13584
rect 8148 13575 8200 13584
rect 8148 13541 8157 13575
rect 8157 13541 8191 13575
rect 8191 13541 8200 13575
rect 8148 13532 8200 13541
rect 9252 13575 9304 13584
rect 9252 13541 9261 13575
rect 9261 13541 9295 13575
rect 9295 13541 9304 13575
rect 9252 13532 9304 13541
rect 11460 13600 11512 13652
rect 11828 13600 11880 13652
rect 15784 13600 15836 13652
rect 18728 13600 18780 13652
rect 20568 13872 20620 13924
rect 22316 13915 22368 13924
rect 22316 13881 22325 13915
rect 22325 13881 22359 13915
rect 22359 13881 22368 13915
rect 22316 13872 22368 13881
rect 23052 13915 23104 13924
rect 23052 13881 23061 13915
rect 23061 13881 23095 13915
rect 23095 13881 23104 13915
rect 23052 13872 23104 13881
rect 23420 13915 23472 13924
rect 23420 13881 23429 13915
rect 23429 13881 23463 13915
rect 23463 13881 23472 13915
rect 23420 13872 23472 13881
rect 23788 13872 23840 13924
rect 20476 13804 20528 13856
rect 20384 13779 20436 13788
rect 20384 13745 20393 13779
rect 20393 13745 20427 13779
rect 20427 13745 20436 13779
rect 20384 13736 20436 13745
rect 21672 13779 21724 13788
rect 21672 13745 21681 13779
rect 21681 13745 21715 13779
rect 21715 13745 21724 13779
rect 21672 13736 21724 13745
rect 22132 13736 22184 13788
rect 23328 13736 23380 13788
rect 19924 13668 19976 13720
rect 21948 13668 22000 13720
rect 11644 13575 11696 13584
rect 11644 13541 11653 13575
rect 11653 13541 11687 13575
rect 11687 13541 11696 13575
rect 11644 13532 11696 13541
rect 13300 13575 13352 13584
rect 13300 13541 13309 13575
rect 13309 13541 13343 13575
rect 13343 13541 13352 13575
rect 13300 13532 13352 13541
rect 18636 13532 18688 13584
rect 19188 13575 19240 13584
rect 19188 13541 19197 13575
rect 19197 13541 19231 13575
rect 19231 13541 19240 13575
rect 19188 13532 19240 13541
rect 19280 13532 19332 13584
rect 21212 13532 21264 13584
rect 3510 13430 3562 13482
rect 3574 13430 3626 13482
rect 3638 13430 3690 13482
rect 3702 13430 3754 13482
rect 3766 13430 3818 13482
rect 2260 13371 2312 13380
rect 2260 13337 2269 13371
rect 2269 13337 2303 13371
rect 2303 13337 2312 13371
rect 2260 13328 2312 13337
rect 2812 13371 2864 13380
rect 2812 13337 2821 13371
rect 2821 13337 2855 13371
rect 2855 13337 2864 13371
rect 2812 13328 2864 13337
rect 3272 13371 3324 13380
rect 3272 13337 3281 13371
rect 3281 13337 3315 13371
rect 3315 13337 3324 13371
rect 3272 13328 3324 13337
rect 4008 13328 4060 13380
rect 5112 13371 5164 13380
rect 5112 13337 5121 13371
rect 5121 13337 5155 13371
rect 5155 13337 5164 13371
rect 5112 13328 5164 13337
rect 6676 13328 6728 13380
rect 6860 13328 6912 13380
rect 7412 13371 7464 13380
rect 7412 13337 7421 13371
rect 7421 13337 7455 13371
rect 7455 13337 7464 13371
rect 7412 13328 7464 13337
rect 3364 13192 3416 13244
rect 4192 13235 4244 13244
rect 4192 13201 4201 13235
rect 4201 13201 4235 13235
rect 4235 13201 4244 13235
rect 4192 13192 4244 13201
rect 6308 13260 6360 13312
rect 7780 13328 7832 13380
rect 8148 13371 8200 13380
rect 8148 13337 8157 13371
rect 8157 13337 8191 13371
rect 8191 13337 8200 13371
rect 10080 13371 10132 13380
rect 8148 13328 8200 13337
rect 10080 13337 10089 13371
rect 10089 13337 10123 13371
rect 10123 13337 10132 13371
rect 10080 13328 10132 13337
rect 10540 13371 10592 13380
rect 10540 13337 10549 13371
rect 10549 13337 10583 13371
rect 10583 13337 10592 13371
rect 10540 13328 10592 13337
rect 15784 13371 15836 13380
rect 15784 13337 15793 13371
rect 15793 13337 15827 13371
rect 15827 13337 15836 13371
rect 15784 13328 15836 13337
rect 15968 13371 16020 13380
rect 15968 13337 15977 13371
rect 15977 13337 16011 13371
rect 16011 13337 16020 13371
rect 15968 13328 16020 13337
rect 17808 13371 17860 13380
rect 17808 13337 17817 13371
rect 17817 13337 17851 13371
rect 17851 13337 17860 13371
rect 17808 13328 17860 13337
rect 18452 13328 18504 13380
rect 18728 13371 18780 13380
rect 18728 13337 18737 13371
rect 18737 13337 18771 13371
rect 18771 13337 18780 13371
rect 18728 13328 18780 13337
rect 18820 13328 18872 13380
rect 19372 13328 19424 13380
rect 20476 13328 20528 13380
rect 21948 13371 22000 13380
rect 21948 13337 21957 13371
rect 21957 13337 21991 13371
rect 21991 13337 22000 13371
rect 21948 13328 22000 13337
rect 22132 13371 22184 13380
rect 22132 13337 22141 13371
rect 22141 13337 22175 13371
rect 22175 13337 22184 13371
rect 22132 13328 22184 13337
rect 23052 13328 23104 13380
rect 8332 13260 8384 13312
rect 8884 13260 8936 13312
rect 9804 13260 9856 13312
rect 11276 13260 11328 13312
rect 1892 13056 1944 13108
rect 4652 13124 4704 13176
rect 5112 13124 5164 13176
rect 5664 13167 5716 13176
rect 5664 13133 5673 13167
rect 5673 13133 5707 13167
rect 5707 13133 5716 13167
rect 5664 13124 5716 13133
rect 5756 13124 5808 13176
rect 4376 13099 4428 13108
rect 4376 13065 4385 13099
rect 4385 13065 4419 13099
rect 4419 13065 4428 13099
rect 4560 13099 4612 13108
rect 4376 13056 4428 13065
rect 4560 13065 4569 13099
rect 4569 13065 4603 13099
rect 4603 13065 4612 13099
rect 4560 13056 4612 13065
rect 5296 13056 5348 13108
rect 6124 13099 6176 13108
rect 6124 13065 6133 13099
rect 6133 13065 6167 13099
rect 6167 13065 6176 13099
rect 6124 13056 6176 13065
rect 7228 13124 7280 13176
rect 7688 13167 7740 13176
rect 7688 13133 7697 13167
rect 7697 13133 7731 13167
rect 7731 13133 7740 13167
rect 7688 13124 7740 13133
rect 13392 13235 13444 13244
rect 6860 13099 6912 13108
rect 6860 13065 6869 13099
rect 6869 13065 6903 13099
rect 6903 13065 6912 13099
rect 6860 13056 6912 13065
rect 7504 13056 7556 13108
rect 8608 13124 8660 13176
rect 8792 13124 8844 13176
rect 9252 13167 9304 13176
rect 9252 13133 9261 13167
rect 9261 13133 9295 13167
rect 9295 13133 9304 13167
rect 9252 13124 9304 13133
rect 9804 13124 9856 13176
rect 9988 13124 10040 13176
rect 13392 13201 13401 13235
rect 13401 13201 13435 13235
rect 13435 13201 13444 13235
rect 13392 13192 13444 13201
rect 17256 13260 17308 13312
rect 18636 13260 18688 13312
rect 19280 13260 19332 13312
rect 21856 13260 21908 13312
rect 24156 13328 24208 13380
rect 21212 13235 21264 13244
rect 21212 13201 21221 13235
rect 21221 13201 21255 13235
rect 21255 13201 21264 13235
rect 21212 13192 21264 13201
rect 23328 13192 23380 13244
rect 23788 13192 23840 13244
rect 11552 13124 11604 13176
rect 13300 13167 13352 13176
rect 11644 13056 11696 13108
rect 1340 13031 1392 13040
rect 1340 12997 1349 13031
rect 1349 12997 1383 13031
rect 1383 12997 1392 13031
rect 1340 12988 1392 12997
rect 1708 12988 1760 13040
rect 4008 12988 4060 13040
rect 5388 12988 5440 13040
rect 5756 12988 5808 13040
rect 6308 13031 6360 13040
rect 6308 12997 6317 13031
rect 6317 12997 6351 13031
rect 6351 12997 6360 13031
rect 6308 12988 6360 12997
rect 6676 12988 6728 13040
rect 7872 12988 7924 13040
rect 8884 13031 8936 13040
rect 8884 12997 8893 13031
rect 8893 12997 8927 13031
rect 8927 12997 8936 13031
rect 8884 12988 8936 12997
rect 9712 13031 9764 13040
rect 9712 12997 9721 13031
rect 9721 12997 9755 13031
rect 9755 12997 9764 13031
rect 9712 12988 9764 12997
rect 10356 13031 10408 13040
rect 10356 12997 10365 13031
rect 10365 12997 10399 13031
rect 10399 12997 10408 13031
rect 10356 12988 10408 12997
rect 12196 13056 12248 13108
rect 13300 13133 13309 13167
rect 13309 13133 13343 13167
rect 13343 13133 13352 13167
rect 13300 13124 13352 13133
rect 13116 13099 13168 13108
rect 13116 13065 13125 13099
rect 13125 13065 13159 13099
rect 13159 13065 13168 13099
rect 17808 13124 17860 13176
rect 19188 13124 19240 13176
rect 20016 13124 20068 13176
rect 20384 13124 20436 13176
rect 21672 13167 21724 13176
rect 13116 13056 13168 13065
rect 17440 13056 17492 13108
rect 20660 13099 20712 13108
rect 20660 13065 20669 13099
rect 20669 13065 20703 13099
rect 20703 13065 20712 13099
rect 20660 13056 20712 13065
rect 21672 13133 21681 13167
rect 21681 13133 21715 13167
rect 21715 13133 21724 13167
rect 21672 13124 21724 13133
rect 21856 13167 21908 13176
rect 21856 13133 21865 13167
rect 21865 13133 21899 13167
rect 21899 13133 21908 13167
rect 21856 13124 21908 13133
rect 22224 13124 22276 13176
rect 24156 13124 24208 13176
rect 21948 13056 22000 13108
rect 23788 13099 23840 13108
rect 23788 13065 23797 13099
rect 23797 13065 23831 13099
rect 23831 13065 23840 13099
rect 23788 13056 23840 13065
rect 21672 12988 21724 13040
rect 25720 12988 25772 13040
rect 18870 12886 18922 12938
rect 18934 12886 18986 12938
rect 18998 12886 19050 12938
rect 19062 12886 19114 12938
rect 19126 12886 19178 12938
rect 1248 12784 1300 12836
rect 2352 12716 2404 12768
rect 7320 12784 7372 12836
rect 7688 12784 7740 12836
rect 8424 12784 8476 12836
rect 9712 12784 9764 12836
rect 12196 12827 12248 12836
rect 12196 12793 12205 12827
rect 12205 12793 12239 12827
rect 12239 12793 12248 12827
rect 12196 12784 12248 12793
rect 13392 12784 13444 12836
rect 20476 12827 20528 12836
rect 20476 12793 20485 12827
rect 20485 12793 20519 12827
rect 20519 12793 20528 12827
rect 20476 12784 20528 12793
rect 20660 12784 20712 12836
rect 4928 12716 4980 12768
rect 6492 12716 6544 12768
rect 7964 12716 8016 12768
rect 17440 12759 17492 12768
rect 17440 12725 17449 12759
rect 17449 12725 17483 12759
rect 17483 12725 17492 12759
rect 17440 12716 17492 12725
rect 1708 12648 1760 12700
rect 1524 12580 1576 12632
rect 4836 12648 4888 12700
rect 7504 12648 7556 12700
rect 7780 12691 7832 12700
rect 7780 12657 7789 12691
rect 7789 12657 7823 12691
rect 7823 12657 7832 12691
rect 7780 12648 7832 12657
rect 9436 12648 9488 12700
rect 11000 12691 11052 12700
rect 11000 12657 11009 12691
rect 11009 12657 11043 12691
rect 11043 12657 11052 12691
rect 11000 12648 11052 12657
rect 11460 12691 11512 12700
rect 11460 12657 11469 12691
rect 11469 12657 11503 12691
rect 11503 12657 11512 12691
rect 11460 12648 11512 12657
rect 4744 12623 4796 12632
rect 4744 12589 4753 12623
rect 4753 12589 4787 12623
rect 4787 12589 4796 12623
rect 4744 12580 4796 12589
rect 5204 12580 5256 12632
rect 6400 12580 6452 12632
rect 7872 12623 7924 12632
rect 7872 12589 7881 12623
rect 7881 12589 7915 12623
rect 7915 12589 7924 12623
rect 7872 12580 7924 12589
rect 8240 12623 8292 12632
rect 8240 12589 8249 12623
rect 8249 12589 8283 12623
rect 8283 12589 8292 12623
rect 8240 12580 8292 12589
rect 8424 12580 8476 12632
rect 9528 12580 9580 12632
rect 10816 12580 10868 12632
rect 15508 12648 15560 12700
rect 17532 12648 17584 12700
rect 18544 12648 18596 12700
rect 23328 12716 23380 12768
rect 21672 12691 21724 12700
rect 21672 12657 21681 12691
rect 21681 12657 21715 12691
rect 21715 12657 21724 12691
rect 21672 12648 21724 12657
rect 21856 12691 21908 12700
rect 21856 12657 21865 12691
rect 21865 12657 21899 12691
rect 21899 12657 21908 12691
rect 21856 12648 21908 12657
rect 22684 12648 22736 12700
rect 24156 12716 24208 12768
rect 24064 12691 24116 12700
rect 24064 12657 24073 12691
rect 24073 12657 24107 12691
rect 24107 12657 24116 12691
rect 24064 12648 24116 12657
rect 15416 12623 15468 12632
rect 4008 12512 4060 12564
rect 2260 12487 2312 12496
rect 2260 12453 2269 12487
rect 2269 12453 2303 12487
rect 2303 12453 2312 12487
rect 2260 12444 2312 12453
rect 4100 12487 4152 12496
rect 4100 12453 4109 12487
rect 4109 12453 4143 12487
rect 4143 12453 4152 12487
rect 4100 12444 4152 12453
rect 4468 12444 4520 12496
rect 6308 12444 6360 12496
rect 6492 12444 6544 12496
rect 7964 12512 8016 12564
rect 11276 12512 11328 12564
rect 15416 12589 15425 12623
rect 15425 12589 15459 12623
rect 15459 12589 15468 12623
rect 15416 12580 15468 12589
rect 21948 12623 22000 12632
rect 21948 12589 21957 12623
rect 21957 12589 21991 12623
rect 21991 12589 22000 12623
rect 21948 12580 22000 12589
rect 22776 12580 22828 12632
rect 23788 12580 23840 12632
rect 23512 12555 23564 12564
rect 23512 12521 23521 12555
rect 23521 12521 23555 12555
rect 23555 12521 23564 12555
rect 23512 12512 23564 12521
rect 7228 12444 7280 12496
rect 8056 12444 8108 12496
rect 9528 12444 9580 12496
rect 14312 12487 14364 12496
rect 14312 12453 14321 12487
rect 14321 12453 14355 12487
rect 14355 12453 14364 12487
rect 14312 12444 14364 12453
rect 15876 12444 15928 12496
rect 17716 12487 17768 12496
rect 17716 12453 17725 12487
rect 17725 12453 17759 12487
rect 17759 12453 17768 12487
rect 17716 12444 17768 12453
rect 3510 12342 3562 12394
rect 3574 12342 3626 12394
rect 3638 12342 3690 12394
rect 3702 12342 3754 12394
rect 3766 12342 3818 12394
rect 1248 12283 1300 12292
rect 1248 12249 1257 12283
rect 1257 12249 1291 12283
rect 1291 12249 1300 12283
rect 1248 12240 1300 12249
rect 1708 12240 1760 12292
rect 5204 12240 5256 12292
rect 6400 12283 6452 12292
rect 6400 12249 6409 12283
rect 6409 12249 6443 12283
rect 6443 12249 6452 12283
rect 6400 12240 6452 12249
rect 6584 12283 6636 12292
rect 6584 12249 6593 12283
rect 6593 12249 6627 12283
rect 6627 12249 6636 12283
rect 6584 12240 6636 12249
rect 7504 12283 7556 12292
rect 7504 12249 7513 12283
rect 7513 12249 7547 12283
rect 7547 12249 7556 12283
rect 7504 12240 7556 12249
rect 8148 12240 8200 12292
rect 8240 12240 8292 12292
rect 9988 12240 10040 12292
rect 11460 12283 11512 12292
rect 11460 12249 11469 12283
rect 11469 12249 11503 12283
rect 11503 12249 11512 12283
rect 11460 12240 11512 12249
rect 17440 12240 17492 12292
rect 17716 12240 17768 12292
rect 20660 12240 20712 12292
rect 21948 12240 22000 12292
rect 22776 12283 22828 12292
rect 22776 12249 22785 12283
rect 22785 12249 22819 12283
rect 22819 12249 22828 12283
rect 22776 12240 22828 12249
rect 23328 12283 23380 12292
rect 23328 12249 23337 12283
rect 23337 12249 23371 12283
rect 23371 12249 23380 12283
rect 23328 12240 23380 12249
rect 23512 12283 23564 12292
rect 23512 12249 23521 12283
rect 23521 12249 23555 12283
rect 23555 12249 23564 12283
rect 23512 12240 23564 12249
rect 2260 12147 2312 12156
rect 2260 12113 2266 12147
rect 2266 12113 2312 12147
rect 2260 12104 2312 12113
rect 2720 12104 2772 12156
rect 3364 12104 3416 12156
rect 4468 12172 4520 12224
rect 4652 12172 4704 12224
rect 4744 12172 4796 12224
rect 2996 12036 3048 12088
rect 3732 12104 3784 12156
rect 5664 12104 5716 12156
rect 7780 12172 7832 12224
rect 11000 12172 11052 12224
rect 12288 12172 12340 12224
rect 17532 12215 17584 12224
rect 17532 12181 17541 12215
rect 17541 12181 17575 12215
rect 17575 12181 17584 12215
rect 17532 12172 17584 12181
rect 20476 12215 20528 12224
rect 20476 12181 20485 12215
rect 20485 12181 20519 12215
rect 20519 12181 20528 12215
rect 20476 12172 20528 12181
rect 22684 12172 22736 12224
rect 14312 12147 14364 12156
rect 14312 12113 14321 12147
rect 14321 12113 14355 12147
rect 14355 12113 14364 12147
rect 14312 12104 14364 12113
rect 21856 12104 21908 12156
rect 4284 12036 4336 12088
rect 6308 12036 6360 12088
rect 7504 12036 7556 12088
rect 4008 12011 4060 12020
rect 1524 11900 1576 11952
rect 2168 11900 2220 11952
rect 4008 11977 4017 12011
rect 4017 11977 4051 12011
rect 4051 11977 4060 12011
rect 4008 11968 4060 11977
rect 4560 11968 4612 12020
rect 3824 11943 3876 11952
rect 3824 11909 3833 11943
rect 3833 11909 3867 11943
rect 3867 11909 3876 11943
rect 3824 11900 3876 11909
rect 4468 11900 4520 11952
rect 4652 11943 4704 11952
rect 4652 11909 4661 11943
rect 4661 11909 4695 11943
rect 4695 11909 4704 11943
rect 4652 11900 4704 11909
rect 4928 11943 4980 11952
rect 4928 11909 4937 11943
rect 4937 11909 4971 11943
rect 4971 11909 4980 11943
rect 4928 11900 4980 11909
rect 5940 11968 5992 12020
rect 7136 11968 7188 12020
rect 8240 12011 8292 12020
rect 8240 11977 8249 12011
rect 8249 11977 8283 12011
rect 8283 11977 8292 12011
rect 8240 11968 8292 11977
rect 11460 12036 11512 12088
rect 23696 12079 23748 12088
rect 23696 12045 23705 12079
rect 23705 12045 23739 12079
rect 23739 12045 23748 12079
rect 23696 12036 23748 12045
rect 8792 12011 8844 12020
rect 8792 11977 8801 12011
rect 8801 11977 8835 12011
rect 8835 11977 8844 12011
rect 8792 11968 8844 11977
rect 14496 11968 14548 12020
rect 15324 11968 15376 12020
rect 16336 12011 16388 12020
rect 16336 11977 16345 12011
rect 16345 11977 16379 12011
rect 16379 11977 16388 12011
rect 16336 11968 16388 11977
rect 21672 11968 21724 12020
rect 6216 11900 6268 11952
rect 7688 11943 7740 11952
rect 7688 11909 7697 11943
rect 7697 11909 7731 11943
rect 7731 11909 7740 11943
rect 7688 11900 7740 11909
rect 8332 11943 8384 11952
rect 8332 11909 8341 11943
rect 8341 11909 8375 11943
rect 8375 11909 8384 11943
rect 8332 11900 8384 11909
rect 10816 11900 10868 11952
rect 11276 11943 11328 11952
rect 11276 11909 11285 11943
rect 11285 11909 11319 11943
rect 11319 11909 11328 11943
rect 11276 11900 11328 11909
rect 24708 11968 24760 12020
rect 25720 12011 25772 12020
rect 25720 11977 25729 12011
rect 25729 11977 25763 12011
rect 25763 11977 25772 12011
rect 25720 11968 25772 11977
rect 24616 11900 24668 11952
rect 18870 11798 18922 11850
rect 18934 11798 18986 11850
rect 18998 11798 19050 11850
rect 19062 11798 19114 11850
rect 19126 11798 19178 11850
rect 2720 11696 2772 11748
rect 3916 11739 3968 11748
rect 3916 11705 3925 11739
rect 3925 11705 3959 11739
rect 3959 11705 3968 11739
rect 3916 11696 3968 11705
rect 4468 11739 4520 11748
rect 4468 11705 4477 11739
rect 4477 11705 4511 11739
rect 4511 11705 4520 11739
rect 4468 11696 4520 11705
rect 1800 11628 1852 11680
rect 3732 11628 3784 11680
rect 1616 11560 1668 11612
rect 3824 11560 3876 11612
rect 4560 11603 4612 11612
rect 4560 11569 4587 11603
rect 4587 11569 4612 11603
rect 7504 11696 7556 11748
rect 7688 11696 7740 11748
rect 8792 11696 8844 11748
rect 10172 11696 10224 11748
rect 10816 11739 10868 11748
rect 10816 11705 10825 11739
rect 10825 11705 10859 11739
rect 10859 11705 10868 11739
rect 10816 11696 10868 11705
rect 15416 11739 15468 11748
rect 15416 11705 15425 11739
rect 15425 11705 15459 11739
rect 15459 11705 15468 11739
rect 15416 11696 15468 11705
rect 23328 11696 23380 11748
rect 24064 11696 24116 11748
rect 25720 11696 25772 11748
rect 5940 11671 5992 11680
rect 5940 11637 5949 11671
rect 5949 11637 5983 11671
rect 5983 11637 5992 11671
rect 5940 11628 5992 11637
rect 6860 11628 6912 11680
rect 7872 11628 7924 11680
rect 9528 11671 9580 11680
rect 9528 11637 9537 11671
rect 9537 11637 9571 11671
rect 9571 11637 9580 11671
rect 9528 11628 9580 11637
rect 13300 11628 13352 11680
rect 15600 11628 15652 11680
rect 16336 11628 16388 11680
rect 24708 11671 24760 11680
rect 24708 11637 24717 11671
rect 24717 11637 24751 11671
rect 24751 11637 24760 11671
rect 24708 11628 24760 11637
rect 4560 11560 4612 11569
rect 5756 11560 5808 11612
rect 6400 11560 6452 11612
rect 7412 11560 7464 11612
rect 9344 11603 9396 11612
rect 9344 11569 9353 11603
rect 9353 11569 9387 11603
rect 9387 11569 9396 11603
rect 9344 11560 9396 11569
rect 10172 11560 10224 11612
rect 12840 11603 12892 11612
rect 12840 11569 12849 11603
rect 12849 11569 12883 11603
rect 12883 11569 12892 11603
rect 12840 11560 12892 11569
rect 15508 11560 15560 11612
rect 23696 11560 23748 11612
rect 24432 11603 24484 11612
rect 24432 11569 24441 11603
rect 24441 11569 24475 11603
rect 24475 11569 24484 11603
rect 24432 11560 24484 11569
rect 2260 11424 2312 11476
rect 4744 11492 4796 11544
rect 4928 11535 4980 11544
rect 4928 11501 4937 11535
rect 4937 11501 4971 11535
rect 4971 11501 4980 11535
rect 4928 11492 4980 11501
rect 6676 11492 6728 11544
rect 1524 11356 1576 11408
rect 2168 11356 2220 11408
rect 5204 11424 5256 11476
rect 5572 11424 5624 11476
rect 6768 11424 6820 11476
rect 8608 11492 8660 11544
rect 9712 11492 9764 11544
rect 12932 11424 12984 11476
rect 14864 11424 14916 11476
rect 4376 11356 4428 11408
rect 6308 11356 6360 11408
rect 8240 11356 8292 11408
rect 11184 11356 11236 11408
rect 11644 11356 11696 11408
rect 13024 11399 13076 11408
rect 13024 11365 13033 11399
rect 13033 11365 13067 11399
rect 13067 11365 13076 11399
rect 13024 11356 13076 11365
rect 13208 11399 13260 11408
rect 13208 11365 13217 11399
rect 13217 11365 13251 11399
rect 13251 11365 13260 11399
rect 13208 11356 13260 11365
rect 13300 11356 13352 11408
rect 13944 11356 13996 11408
rect 14772 11356 14824 11408
rect 3510 11254 3562 11306
rect 3574 11254 3626 11306
rect 3638 11254 3690 11306
rect 3702 11254 3754 11306
rect 3766 11254 3818 11306
rect 1616 11195 1668 11204
rect 1616 11161 1625 11195
rect 1625 11161 1659 11195
rect 1659 11161 1668 11195
rect 1616 11152 1668 11161
rect 1800 11195 1852 11204
rect 1800 11161 1809 11195
rect 1809 11161 1843 11195
rect 1843 11161 1852 11195
rect 1800 11152 1852 11161
rect 2352 11195 2404 11204
rect 2352 11161 2361 11195
rect 2361 11161 2395 11195
rect 2395 11161 2404 11195
rect 2352 11152 2404 11161
rect 2536 11152 2588 11204
rect 3364 11195 3416 11204
rect 3364 11161 3373 11195
rect 3373 11161 3407 11195
rect 3407 11161 3416 11195
rect 3364 11152 3416 11161
rect 4008 11152 4060 11204
rect 4376 11195 4428 11204
rect 4376 11161 4385 11195
rect 4385 11161 4419 11195
rect 4419 11161 4428 11195
rect 4376 11152 4428 11161
rect 4468 11152 4520 11204
rect 5940 11152 5992 11204
rect 6676 11195 6728 11204
rect 6676 11161 6685 11195
rect 6685 11161 6719 11195
rect 6719 11161 6728 11195
rect 6676 11152 6728 11161
rect 3916 11084 3968 11136
rect 2628 10948 2680 11000
rect 2904 11016 2956 11068
rect 4652 11084 4704 11136
rect 5572 11084 5624 11136
rect 6400 11127 6452 11136
rect 6400 11093 6409 11127
rect 6409 11093 6443 11127
rect 6443 11093 6452 11127
rect 6400 11084 6452 11093
rect 7780 11152 7832 11204
rect 10172 11152 10224 11204
rect 10816 11195 10868 11204
rect 10816 11161 10825 11195
rect 10825 11161 10859 11195
rect 10859 11161 10868 11195
rect 10816 11152 10868 11161
rect 13944 11195 13996 11204
rect 13944 11161 13953 11195
rect 13953 11161 13987 11195
rect 13987 11161 13996 11195
rect 13944 11152 13996 11161
rect 14128 11152 14180 11204
rect 14220 11152 14272 11204
rect 9436 11084 9488 11136
rect 9620 11084 9672 11136
rect 13484 11084 13536 11136
rect 3272 10991 3324 11000
rect 3272 10957 3281 10991
rect 3281 10957 3315 10991
rect 3315 10957 3324 10991
rect 3272 10948 3324 10957
rect 4192 10948 4244 11000
rect 4652 10948 4704 11000
rect 4744 10948 4796 11000
rect 8884 11016 8936 11068
rect 9712 11059 9764 11068
rect 9712 11025 9721 11059
rect 9721 11025 9755 11059
rect 9755 11025 9764 11059
rect 9712 11016 9764 11025
rect 10172 11016 10224 11068
rect 11736 11016 11788 11068
rect 12840 11059 12892 11068
rect 12840 11025 12849 11059
rect 12849 11025 12883 11059
rect 12883 11025 12892 11059
rect 24432 11195 24484 11204
rect 24432 11161 24441 11195
rect 24441 11161 24475 11195
rect 24475 11161 24484 11195
rect 24432 11152 24484 11161
rect 24708 11195 24760 11204
rect 24708 11161 24717 11195
rect 24717 11161 24751 11195
rect 24751 11161 24760 11195
rect 24708 11152 24760 11161
rect 14772 11127 14824 11136
rect 14772 11093 14781 11127
rect 14781 11093 14815 11127
rect 14815 11093 14824 11127
rect 14772 11084 14824 11093
rect 19280 11084 19332 11136
rect 12840 11016 12892 11025
rect 14864 11059 14916 11068
rect 7872 10948 7924 11000
rect 1524 10880 1576 10932
rect 3364 10880 3416 10932
rect 2996 10855 3048 10864
rect 2996 10821 3005 10855
rect 3005 10821 3039 10855
rect 3039 10821 3048 10855
rect 2996 10812 3048 10821
rect 5204 10855 5256 10864
rect 5204 10821 5213 10855
rect 5213 10821 5247 10855
rect 5247 10821 5256 10855
rect 5204 10812 5256 10821
rect 7228 10855 7280 10864
rect 7228 10821 7237 10855
rect 7237 10821 7271 10855
rect 7271 10821 7280 10855
rect 8608 10948 8660 11000
rect 9528 10948 9580 11000
rect 11276 10948 11328 11000
rect 12564 10948 12616 11000
rect 8700 10880 8752 10932
rect 9344 10923 9396 10932
rect 9344 10889 9353 10923
rect 9353 10889 9387 10923
rect 9387 10889 9396 10923
rect 9344 10880 9396 10889
rect 11184 10880 11236 10932
rect 13208 10948 13260 11000
rect 13300 10991 13352 11000
rect 13300 10957 13309 10991
rect 13309 10957 13343 10991
rect 13343 10957 13352 10991
rect 13300 10948 13352 10957
rect 14220 10923 14272 10932
rect 14220 10889 14229 10923
rect 14229 10889 14263 10923
rect 14263 10889 14272 10923
rect 14220 10880 14272 10889
rect 7228 10812 7280 10821
rect 9068 10812 9120 10864
rect 12288 10812 12340 10864
rect 13024 10812 13076 10864
rect 14864 11025 14873 11059
rect 14873 11025 14907 11059
rect 14907 11025 14916 11059
rect 14864 11016 14916 11025
rect 15508 11016 15560 11068
rect 18728 10991 18780 11000
rect 18728 10957 18737 10991
rect 18737 10957 18771 10991
rect 18771 10957 18780 10991
rect 18728 10948 18780 10957
rect 19372 10948 19424 11000
rect 24432 11016 24484 11068
rect 17992 10880 18044 10932
rect 20936 10880 20988 10932
rect 18870 10710 18922 10762
rect 18934 10710 18986 10762
rect 18998 10710 19050 10762
rect 19062 10710 19114 10762
rect 19126 10710 19178 10762
rect 2076 10608 2128 10660
rect 2352 10608 2404 10660
rect 2996 10608 3048 10660
rect 4284 10608 4336 10660
rect 4468 10608 4520 10660
rect 7780 10608 7832 10660
rect 8516 10608 8568 10660
rect 3180 10472 3232 10524
rect 4928 10540 4980 10592
rect 5664 10583 5716 10592
rect 5664 10549 5673 10583
rect 5673 10549 5707 10583
rect 5707 10549 5716 10583
rect 5664 10540 5716 10549
rect 8332 10540 8384 10592
rect 8792 10540 8844 10592
rect 9068 10540 9120 10592
rect 9436 10540 9488 10592
rect 14772 10608 14824 10660
rect 19280 10651 19332 10660
rect 3916 10515 3968 10524
rect 3916 10481 3925 10515
rect 3925 10481 3959 10515
rect 3959 10481 3968 10515
rect 3916 10472 3968 10481
rect 4284 10515 4336 10524
rect 4284 10481 4293 10515
rect 4293 10481 4327 10515
rect 4327 10481 4336 10515
rect 4284 10472 4336 10481
rect 4468 10472 4520 10524
rect 5296 10515 5348 10524
rect 5296 10481 5305 10515
rect 5305 10481 5339 10515
rect 5339 10481 5348 10515
rect 5296 10472 5348 10481
rect 9252 10515 9304 10524
rect 9252 10481 9261 10515
rect 9261 10481 9295 10515
rect 9295 10481 9304 10515
rect 9252 10472 9304 10481
rect 12288 10515 12340 10524
rect 12288 10481 12297 10515
rect 12297 10481 12331 10515
rect 12331 10481 12340 10515
rect 12288 10472 12340 10481
rect 12748 10515 12800 10524
rect 12748 10481 12757 10515
rect 12757 10481 12791 10515
rect 12791 10481 12800 10515
rect 12748 10472 12800 10481
rect 14220 10540 14272 10592
rect 13852 10472 13904 10524
rect 15600 10515 15652 10524
rect 15600 10481 15609 10515
rect 15609 10481 15643 10515
rect 15643 10481 15652 10515
rect 15600 10472 15652 10481
rect 19280 10617 19289 10651
rect 19289 10617 19323 10651
rect 19323 10617 19332 10651
rect 19280 10608 19332 10617
rect 15876 10540 15928 10592
rect 17992 10515 18044 10524
rect 4744 10404 4796 10456
rect 8700 10404 8752 10456
rect 15324 10447 15376 10456
rect 15324 10413 15333 10447
rect 15333 10413 15367 10447
rect 15367 10413 15376 10447
rect 15324 10404 15376 10413
rect 17992 10481 18001 10515
rect 18001 10481 18035 10515
rect 18035 10481 18044 10515
rect 17992 10472 18044 10481
rect 18360 10515 18412 10524
rect 18360 10481 18369 10515
rect 18369 10481 18403 10515
rect 18403 10481 18412 10515
rect 18360 10472 18412 10481
rect 18544 10515 18596 10524
rect 18544 10481 18553 10515
rect 18553 10481 18587 10515
rect 18587 10481 18596 10515
rect 18544 10472 18596 10481
rect 20936 10540 20988 10592
rect 22684 10608 22736 10660
rect 23236 10608 23288 10660
rect 23788 10651 23840 10660
rect 23788 10617 23797 10651
rect 23797 10617 23831 10651
rect 23831 10617 23840 10651
rect 23788 10608 23840 10617
rect 23052 10472 23104 10524
rect 23328 10515 23380 10524
rect 23328 10481 23337 10515
rect 23337 10481 23371 10515
rect 23371 10481 23380 10515
rect 23328 10472 23380 10481
rect 23788 10472 23840 10524
rect 24432 10515 24484 10524
rect 24432 10481 24441 10515
rect 24441 10481 24475 10515
rect 24475 10481 24484 10515
rect 24432 10472 24484 10481
rect 18084 10404 18136 10456
rect 20476 10447 20528 10456
rect 20476 10413 20485 10447
rect 20485 10413 20519 10447
rect 20519 10413 20528 10447
rect 20476 10404 20528 10413
rect 22224 10447 22276 10456
rect 22224 10413 22233 10447
rect 22233 10413 22267 10447
rect 22267 10413 22276 10447
rect 22224 10404 22276 10413
rect 23512 10404 23564 10456
rect 24708 10447 24760 10456
rect 24708 10413 24717 10447
rect 24717 10413 24751 10447
rect 24751 10413 24760 10447
rect 24708 10404 24760 10413
rect 3916 10268 3968 10320
rect 4652 10336 4704 10388
rect 8240 10336 8292 10388
rect 9528 10336 9580 10388
rect 13116 10379 13168 10388
rect 13116 10345 13125 10379
rect 13125 10345 13159 10379
rect 13159 10345 13168 10379
rect 13116 10336 13168 10345
rect 14404 10311 14456 10320
rect 14404 10277 14413 10311
rect 14413 10277 14447 10311
rect 14447 10277 14456 10311
rect 14404 10268 14456 10277
rect 15140 10268 15192 10320
rect 16980 10268 17032 10320
rect 18728 10268 18780 10320
rect 19096 10311 19148 10320
rect 19096 10277 19105 10311
rect 19105 10277 19139 10311
rect 19139 10277 19148 10311
rect 19096 10268 19148 10277
rect 20292 10268 20344 10320
rect 24064 10311 24116 10320
rect 24064 10277 24073 10311
rect 24073 10277 24107 10311
rect 24107 10277 24116 10311
rect 24064 10268 24116 10277
rect 3510 10166 3562 10218
rect 3574 10166 3626 10218
rect 3638 10166 3690 10218
rect 3702 10166 3754 10218
rect 3766 10166 3818 10218
rect 1340 10064 1392 10116
rect 2628 10107 2680 10116
rect 2628 10073 2637 10107
rect 2637 10073 2671 10107
rect 2671 10073 2680 10107
rect 2628 10064 2680 10073
rect 2996 10107 3048 10116
rect 2996 10073 3005 10107
rect 3005 10073 3039 10107
rect 3039 10073 3048 10107
rect 2996 10064 3048 10073
rect 3180 10107 3232 10116
rect 3180 10073 3189 10107
rect 3189 10073 3223 10107
rect 3223 10073 3232 10107
rect 3180 10064 3232 10073
rect 4192 10107 4244 10116
rect 4192 10073 4201 10107
rect 4201 10073 4235 10107
rect 4235 10073 4244 10107
rect 4192 10064 4244 10073
rect 4652 10064 4704 10116
rect 5296 10064 5348 10116
rect 5664 10064 5716 10116
rect 6768 10107 6820 10116
rect 6768 10073 6777 10107
rect 6777 10073 6811 10107
rect 6811 10073 6820 10107
rect 6768 10064 6820 10073
rect 7136 10064 7188 10116
rect 8516 10064 8568 10116
rect 9068 10064 9120 10116
rect 11460 10107 11512 10116
rect 11460 10073 11469 10107
rect 11469 10073 11503 10107
rect 11503 10073 11512 10107
rect 11460 10064 11512 10073
rect 12748 10064 12800 10116
rect 13116 10107 13168 10116
rect 13116 10073 13125 10107
rect 13125 10073 13159 10107
rect 13159 10073 13168 10107
rect 13116 10064 13168 10073
rect 13852 10107 13904 10116
rect 13852 10073 13861 10107
rect 13861 10073 13895 10107
rect 13895 10073 13904 10107
rect 13852 10064 13904 10073
rect 14496 10064 14548 10116
rect 16980 10107 17032 10116
rect 16980 10073 16989 10107
rect 16989 10073 17023 10107
rect 17023 10073 17032 10107
rect 16980 10064 17032 10073
rect 17348 10064 17400 10116
rect 18544 10064 18596 10116
rect 3088 9996 3140 10048
rect 2628 9928 2680 9980
rect 4560 9860 4612 9912
rect 6124 9860 6176 9912
rect 7228 9928 7280 9980
rect 8240 9996 8292 10048
rect 8792 9996 8844 10048
rect 14312 9996 14364 10048
rect 9068 9928 9120 9980
rect 10356 9928 10408 9980
rect 12288 9971 12340 9980
rect 12288 9937 12297 9971
rect 12297 9937 12331 9971
rect 12331 9937 12340 9971
rect 12288 9928 12340 9937
rect 18360 9996 18412 10048
rect 20476 10064 20528 10116
rect 20936 10107 20988 10116
rect 20936 10073 20945 10107
rect 20945 10073 20979 10107
rect 20979 10073 20988 10107
rect 20936 10064 20988 10073
rect 23236 10107 23288 10116
rect 23236 10073 23245 10107
rect 23245 10073 23279 10107
rect 23279 10073 23288 10107
rect 23236 10064 23288 10073
rect 23512 10107 23564 10116
rect 23512 10073 23521 10107
rect 23521 10073 23555 10107
rect 23555 10073 23564 10107
rect 23512 10064 23564 10073
rect 23880 10064 23932 10116
rect 2076 9792 2128 9844
rect 1800 9724 1852 9776
rect 4100 9792 4152 9844
rect 4376 9724 4428 9776
rect 6492 9792 6544 9844
rect 8700 9860 8752 9912
rect 8884 9860 8936 9912
rect 9252 9860 9304 9912
rect 12012 9903 12064 9912
rect 12012 9869 12021 9903
rect 12021 9869 12055 9903
rect 12055 9869 12064 9903
rect 12012 9860 12064 9869
rect 13392 9860 13444 9912
rect 15140 9903 15192 9912
rect 15140 9869 15149 9903
rect 15149 9869 15183 9903
rect 15183 9869 15192 9903
rect 15140 9860 15192 9869
rect 15600 9903 15652 9912
rect 8608 9835 8660 9844
rect 8608 9801 8617 9835
rect 8617 9801 8651 9835
rect 8651 9801 8660 9835
rect 8608 9792 8660 9801
rect 8240 9767 8292 9776
rect 8240 9733 8249 9767
rect 8249 9733 8283 9767
rect 8283 9733 8292 9767
rect 8240 9724 8292 9733
rect 8516 9767 8568 9776
rect 8516 9733 8525 9767
rect 8525 9733 8559 9767
rect 8559 9733 8568 9767
rect 9344 9835 9396 9844
rect 8884 9767 8936 9776
rect 8516 9724 8568 9733
rect 8884 9733 8893 9767
rect 8893 9733 8927 9767
rect 8927 9733 8936 9767
rect 8884 9724 8936 9733
rect 9344 9801 9353 9835
rect 9353 9801 9387 9835
rect 9387 9801 9396 9835
rect 9344 9792 9396 9801
rect 14220 9792 14272 9844
rect 14312 9792 14364 9844
rect 15600 9869 15609 9903
rect 15609 9869 15643 9903
rect 15643 9869 15652 9903
rect 15600 9860 15652 9869
rect 15692 9860 15744 9912
rect 19280 9860 19332 9912
rect 19740 9903 19792 9912
rect 19740 9869 19749 9903
rect 19749 9869 19783 9903
rect 19783 9869 19792 9903
rect 19740 9860 19792 9869
rect 19096 9792 19148 9844
rect 20292 9928 20344 9980
rect 22224 9928 22276 9980
rect 20476 9860 20528 9912
rect 24064 9928 24116 9980
rect 25444 9928 25496 9980
rect 9436 9767 9488 9776
rect 9436 9733 9445 9767
rect 9445 9733 9479 9767
rect 9479 9733 9488 9767
rect 9436 9724 9488 9733
rect 13392 9724 13444 9776
rect 15692 9724 15744 9776
rect 15784 9724 15836 9776
rect 17348 9767 17400 9776
rect 17348 9733 17357 9767
rect 17357 9733 17391 9767
rect 17391 9733 17400 9767
rect 17348 9724 17400 9733
rect 17440 9724 17492 9776
rect 17992 9724 18044 9776
rect 21304 9792 21356 9844
rect 24708 9792 24760 9844
rect 22224 9724 22276 9776
rect 23052 9767 23104 9776
rect 23052 9733 23061 9767
rect 23061 9733 23095 9767
rect 23095 9733 23104 9767
rect 23052 9724 23104 9733
rect 23604 9767 23656 9776
rect 23604 9733 23613 9767
rect 23613 9733 23647 9767
rect 23647 9733 23656 9767
rect 23604 9724 23656 9733
rect 18870 9622 18922 9674
rect 18934 9622 18986 9674
rect 18998 9622 19050 9674
rect 19062 9622 19114 9674
rect 19126 9622 19178 9674
rect 512 9520 564 9572
rect 788 9520 840 9572
rect 1800 9563 1852 9572
rect 1800 9529 1809 9563
rect 1809 9529 1843 9563
rect 1843 9529 1852 9563
rect 1800 9520 1852 9529
rect 1616 9452 1668 9504
rect 2076 9520 2128 9572
rect 3272 9520 3324 9572
rect 3180 9452 3232 9504
rect 5204 9452 5256 9504
rect 7412 9520 7464 9572
rect 9344 9520 9396 9572
rect 12564 9563 12616 9572
rect 12564 9529 12573 9563
rect 12573 9529 12607 9563
rect 12607 9529 12616 9563
rect 12564 9520 12616 9529
rect 15324 9520 15376 9572
rect 18084 9520 18136 9572
rect 19740 9520 19792 9572
rect 20292 9563 20344 9572
rect 20292 9529 20301 9563
rect 20301 9529 20335 9563
rect 20335 9529 20344 9563
rect 20292 9520 20344 9529
rect 23788 9520 23840 9572
rect 24708 9563 24760 9572
rect 6400 9452 6452 9504
rect 14404 9495 14456 9504
rect 14404 9461 14413 9495
rect 14413 9461 14447 9495
rect 14447 9461 14456 9495
rect 14404 9452 14456 9461
rect 15600 9452 15652 9504
rect 19280 9495 19332 9504
rect 19280 9461 19289 9495
rect 19289 9461 19323 9495
rect 19323 9461 19332 9495
rect 19280 9452 19332 9461
rect 23052 9452 23104 9504
rect 24708 9529 24717 9563
rect 24717 9529 24751 9563
rect 24751 9529 24760 9563
rect 24708 9520 24760 9529
rect 2352 9384 2404 9436
rect 3364 9384 3416 9436
rect 4192 9384 4244 9436
rect 4560 9427 4612 9436
rect 4560 9393 4569 9427
rect 4569 9393 4603 9427
rect 4603 9393 4612 9427
rect 4560 9384 4612 9393
rect 6676 9427 6728 9436
rect 2536 9316 2588 9368
rect 2996 9316 3048 9368
rect 6676 9393 6685 9427
rect 6685 9393 6719 9427
rect 6719 9393 6728 9427
rect 6676 9384 6728 9393
rect 6952 9427 7004 9436
rect 6952 9393 6961 9427
rect 6961 9393 6995 9427
rect 6995 9393 7004 9427
rect 6952 9384 7004 9393
rect 9068 9427 9120 9436
rect 9068 9393 9077 9427
rect 9077 9393 9111 9427
rect 9111 9393 9120 9427
rect 9068 9384 9120 9393
rect 11184 9427 11236 9436
rect 11184 9393 11193 9427
rect 11193 9393 11227 9427
rect 11227 9393 11236 9427
rect 11184 9384 11236 9393
rect 12472 9427 12524 9436
rect 12472 9393 12481 9427
rect 12481 9393 12515 9427
rect 12515 9393 12524 9427
rect 12472 9384 12524 9393
rect 13300 9384 13352 9436
rect 14128 9384 14180 9436
rect 14772 9384 14824 9436
rect 16428 9384 16480 9436
rect 17716 9384 17768 9436
rect 18728 9427 18780 9436
rect 18728 9393 18737 9427
rect 18737 9393 18771 9427
rect 18771 9393 18780 9427
rect 18728 9384 18780 9393
rect 18912 9427 18964 9436
rect 18912 9393 18921 9427
rect 18921 9393 18955 9427
rect 18955 9393 18964 9427
rect 18912 9384 18964 9393
rect 19372 9384 19424 9436
rect 23420 9427 23472 9436
rect 23420 9393 23429 9427
rect 23429 9393 23463 9427
rect 23463 9393 23472 9427
rect 23420 9384 23472 9393
rect 23696 9427 23748 9436
rect 23696 9393 23705 9427
rect 23705 9393 23739 9427
rect 23739 9393 23748 9427
rect 23696 9384 23748 9393
rect 25076 9452 25128 9504
rect 24156 9427 24208 9436
rect 24156 9393 24165 9427
rect 24165 9393 24199 9427
rect 24199 9393 24208 9427
rect 24156 9384 24208 9393
rect 5112 9359 5164 9368
rect 5112 9325 5121 9359
rect 5121 9325 5155 9359
rect 5155 9325 5164 9359
rect 5112 9316 5164 9325
rect 3916 9248 3968 9300
rect 4376 9248 4428 9300
rect 3088 9180 3140 9232
rect 4284 9180 4336 9232
rect 4928 9180 4980 9232
rect 6768 9316 6820 9368
rect 7136 9359 7188 9368
rect 7136 9325 7145 9359
rect 7145 9325 7179 9359
rect 7179 9325 7188 9359
rect 7136 9316 7188 9325
rect 11092 9359 11144 9368
rect 6676 9248 6728 9300
rect 8608 9248 8660 9300
rect 11092 9325 11101 9359
rect 11101 9325 11135 9359
rect 11135 9325 11144 9359
rect 11092 9316 11144 9325
rect 13852 9316 13904 9368
rect 15324 9316 15376 9368
rect 9344 9248 9396 9300
rect 23328 9316 23380 9368
rect 25168 9316 25220 9368
rect 16520 9248 16572 9300
rect 23052 9248 23104 9300
rect 23604 9248 23656 9300
rect 6584 9180 6636 9232
rect 7872 9180 7924 9232
rect 9252 9223 9304 9232
rect 9252 9189 9261 9223
rect 9261 9189 9295 9223
rect 9295 9189 9304 9223
rect 9252 9180 9304 9189
rect 11276 9180 11328 9232
rect 14864 9223 14916 9232
rect 14864 9189 14873 9223
rect 14873 9189 14907 9223
rect 14907 9189 14916 9223
rect 14864 9180 14916 9189
rect 15232 9223 15284 9232
rect 15232 9189 15241 9223
rect 15241 9189 15275 9223
rect 15275 9189 15284 9223
rect 15232 9180 15284 9189
rect 22776 9180 22828 9232
rect 23696 9180 23748 9232
rect 3510 9078 3562 9130
rect 3574 9078 3626 9130
rect 3638 9078 3690 9130
rect 3702 9078 3754 9130
rect 3766 9078 3818 9130
rect 2076 9019 2128 9028
rect 2076 8985 2085 9019
rect 2085 8985 2119 9019
rect 2119 8985 2128 9019
rect 2076 8976 2128 8985
rect 2996 9019 3048 9028
rect 2996 8985 3005 9019
rect 3005 8985 3039 9019
rect 3039 8985 3048 9019
rect 2996 8976 3048 8985
rect 3180 9019 3232 9028
rect 3180 8985 3189 9019
rect 3189 8985 3223 9019
rect 3223 8985 3232 9019
rect 3180 8976 3232 8985
rect 3916 8976 3968 9028
rect 4284 9019 4336 9028
rect 4284 8985 4293 9019
rect 4293 8985 4327 9019
rect 4327 8985 4336 9019
rect 4928 9019 4980 9028
rect 4284 8976 4336 8985
rect 4928 8985 4937 9019
rect 4937 8985 4971 9019
rect 4971 8985 4980 9019
rect 4928 8976 4980 8985
rect 6952 8976 7004 9028
rect 9068 9019 9120 9028
rect 9068 8985 9077 9019
rect 9077 8985 9111 9019
rect 9111 8985 9120 9019
rect 9068 8976 9120 8985
rect 9252 9019 9304 9028
rect 9252 8985 9261 9019
rect 9261 8985 9295 9019
rect 9295 8985 9304 9019
rect 9252 8976 9304 8985
rect 9344 9019 9396 9028
rect 9344 8985 9353 9019
rect 9353 8985 9387 9019
rect 9387 8985 9396 9019
rect 9344 8976 9396 8985
rect 11092 8976 11144 9028
rect 11460 8976 11512 9028
rect 12564 8976 12616 9028
rect 2352 8908 2404 8960
rect 3088 8908 3140 8960
rect 4560 8908 4612 8960
rect 696 8840 748 8892
rect 4192 8840 4244 8892
rect 6768 8908 6820 8960
rect 8884 8908 8936 8960
rect 12472 8908 12524 8960
rect 788 8815 840 8824
rect 788 8781 797 8815
rect 797 8781 831 8815
rect 831 8781 840 8815
rect 788 8772 840 8781
rect 1616 8815 1668 8824
rect 1616 8781 1625 8815
rect 1625 8781 1659 8815
rect 1659 8781 1668 8815
rect 1616 8772 1668 8781
rect 880 8747 932 8756
rect 880 8713 889 8747
rect 889 8713 923 8747
rect 923 8713 932 8747
rect 880 8704 932 8713
rect 2536 8636 2588 8688
rect 4376 8772 4428 8824
rect 6216 8840 6268 8892
rect 8240 8840 8292 8892
rect 9068 8840 9120 8892
rect 11184 8840 11236 8892
rect 13392 8951 13444 8960
rect 13392 8917 13401 8951
rect 13401 8917 13435 8951
rect 13435 8917 13444 8951
rect 13392 8908 13444 8917
rect 11276 8815 11328 8824
rect 4192 8704 4244 8756
rect 6216 8704 6268 8756
rect 6492 8747 6544 8756
rect 6492 8713 6501 8747
rect 6501 8713 6535 8747
rect 6535 8713 6544 8747
rect 6492 8704 6544 8713
rect 6860 8747 6912 8756
rect 6860 8713 6869 8747
rect 6869 8713 6903 8747
rect 6903 8713 6912 8747
rect 6860 8704 6912 8713
rect 11276 8781 11285 8815
rect 11285 8781 11319 8815
rect 11319 8781 11328 8815
rect 11276 8772 11328 8781
rect 13116 8815 13168 8824
rect 13116 8781 13125 8815
rect 13125 8781 13159 8815
rect 13159 8781 13168 8815
rect 13116 8772 13168 8781
rect 8516 8747 8568 8756
rect 8516 8713 8525 8747
rect 8525 8713 8559 8747
rect 8559 8713 8568 8747
rect 8516 8704 8568 8713
rect 11368 8704 11420 8756
rect 13024 8704 13076 8756
rect 14864 8976 14916 9028
rect 15324 9019 15376 9028
rect 15324 8985 15333 9019
rect 15333 8985 15367 9019
rect 15367 8985 15376 9019
rect 15324 8976 15376 8985
rect 16428 9019 16480 9028
rect 16428 8985 16437 9019
rect 16437 8985 16471 9019
rect 16471 8985 16480 9019
rect 16428 8976 16480 8985
rect 16520 9019 16572 9028
rect 16520 8985 16529 9019
rect 16529 8985 16563 9019
rect 16563 8985 16572 9019
rect 16520 8976 16572 8985
rect 18728 8976 18780 9028
rect 19280 9019 19332 9028
rect 19280 8985 19289 9019
rect 19289 8985 19323 9019
rect 19323 8985 19332 9019
rect 19280 8976 19332 8985
rect 20476 8976 20528 9028
rect 21488 8976 21540 9028
rect 22224 9019 22276 9028
rect 22224 8985 22233 9019
rect 22233 8985 22267 9019
rect 22267 8985 22276 9019
rect 22224 8976 22276 8985
rect 22776 9019 22828 9028
rect 22776 8985 22785 9019
rect 22785 8985 22819 9019
rect 22819 8985 22828 9019
rect 22776 8976 22828 8985
rect 23052 9019 23104 9028
rect 23052 8985 23061 9019
rect 23061 8985 23095 9019
rect 23095 8985 23104 9019
rect 23052 8976 23104 8985
rect 23420 9019 23472 9028
rect 23420 8985 23429 9019
rect 23429 8985 23463 9019
rect 23463 8985 23472 9019
rect 23420 8976 23472 8985
rect 25444 9019 25496 9028
rect 25444 8985 25453 9019
rect 25453 8985 25487 9019
rect 25487 8985 25496 9019
rect 25444 8976 25496 8985
rect 14220 8951 14272 8960
rect 14220 8917 14229 8951
rect 14229 8917 14263 8951
rect 14263 8917 14272 8951
rect 14220 8908 14272 8917
rect 18912 8951 18964 8960
rect 18912 8917 18921 8951
rect 18921 8917 18955 8951
rect 18955 8917 18964 8951
rect 18912 8908 18964 8917
rect 15232 8840 15284 8892
rect 14680 8815 14732 8824
rect 14680 8781 14689 8815
rect 14689 8781 14723 8815
rect 14723 8781 14732 8815
rect 14680 8772 14732 8781
rect 16520 8772 16572 8824
rect 17716 8772 17768 8824
rect 18268 8840 18320 8892
rect 14496 8747 14548 8756
rect 14496 8713 14505 8747
rect 14505 8713 14539 8747
rect 14539 8713 14548 8747
rect 14496 8704 14548 8713
rect 18452 8815 18504 8824
rect 18452 8781 18461 8815
rect 18461 8781 18495 8815
rect 18495 8781 18504 8815
rect 21304 8815 21356 8824
rect 18452 8772 18504 8781
rect 21304 8781 21313 8815
rect 21313 8781 21347 8815
rect 21347 8781 21356 8815
rect 21304 8772 21356 8781
rect 18360 8704 18412 8756
rect 4744 8679 4796 8688
rect 4744 8645 4753 8679
rect 4753 8645 4787 8679
rect 4787 8645 4796 8679
rect 4744 8636 4796 8645
rect 6308 8679 6360 8688
rect 6308 8645 6317 8679
rect 6317 8645 6351 8679
rect 6351 8645 6360 8679
rect 6308 8636 6360 8645
rect 6676 8636 6728 8688
rect 18268 8636 18320 8688
rect 23328 8772 23380 8824
rect 23512 8704 23564 8756
rect 25168 8883 25220 8892
rect 25168 8849 25177 8883
rect 25177 8849 25211 8883
rect 25211 8849 25220 8883
rect 25168 8840 25220 8849
rect 25444 8772 25496 8824
rect 18870 8534 18922 8586
rect 18934 8534 18986 8586
rect 18998 8534 19050 8586
rect 19062 8534 19114 8586
rect 19126 8534 19178 8586
rect 696 8475 748 8484
rect 696 8441 705 8475
rect 705 8441 739 8475
rect 739 8441 748 8475
rect 696 8432 748 8441
rect 880 8475 932 8484
rect 880 8441 889 8475
rect 889 8441 923 8475
rect 923 8441 932 8475
rect 880 8432 932 8441
rect 3364 8432 3416 8484
rect 4376 8364 4428 8416
rect 4652 8432 4704 8484
rect 5296 8432 5348 8484
rect 6860 8432 6912 8484
rect 9068 8475 9120 8484
rect 9068 8441 9077 8475
rect 9077 8441 9111 8475
rect 9111 8441 9120 8475
rect 9068 8432 9120 8441
rect 13392 8432 13444 8484
rect 14772 8432 14824 8484
rect 23328 8432 23380 8484
rect 6400 8407 6452 8416
rect 6400 8373 6409 8407
rect 6409 8373 6443 8407
rect 6443 8373 6452 8407
rect 6400 8364 6452 8373
rect 6676 8407 6728 8416
rect 6676 8373 6685 8407
rect 6685 8373 6719 8407
rect 6719 8373 6728 8407
rect 6676 8364 6728 8373
rect 11368 8364 11420 8416
rect 12012 8364 12064 8416
rect 1524 8296 1576 8348
rect 1616 8339 1668 8348
rect 1616 8305 1625 8339
rect 1625 8305 1659 8339
rect 1659 8305 1668 8339
rect 1616 8296 1668 8305
rect 4008 8296 4060 8348
rect 4192 8296 4244 8348
rect 4744 8296 4796 8348
rect 5756 8339 5808 8348
rect 5756 8305 5765 8339
rect 5765 8305 5799 8339
rect 5799 8305 5808 8339
rect 5756 8296 5808 8305
rect 8424 8296 8476 8348
rect 8976 8339 9028 8348
rect 8976 8305 8985 8339
rect 8985 8305 9019 8339
rect 9019 8305 9028 8339
rect 8976 8296 9028 8305
rect 11460 8339 11512 8348
rect 11460 8305 11469 8339
rect 11469 8305 11503 8339
rect 11503 8305 11512 8339
rect 11460 8296 11512 8305
rect 9068 8228 9120 8280
rect 14680 8228 14732 8280
rect 14772 8271 14824 8280
rect 14772 8237 14781 8271
rect 14781 8237 14815 8271
rect 14815 8237 14824 8271
rect 15324 8296 15376 8348
rect 15600 8339 15652 8348
rect 15600 8305 15609 8339
rect 15609 8305 15643 8339
rect 15643 8305 15652 8339
rect 15600 8296 15652 8305
rect 16428 8296 16480 8348
rect 17716 8339 17768 8348
rect 17716 8305 17725 8339
rect 17725 8305 17759 8339
rect 17759 8305 17768 8339
rect 17716 8296 17768 8305
rect 18268 8339 18320 8348
rect 18268 8305 18277 8339
rect 18277 8305 18311 8339
rect 18311 8305 18320 8339
rect 18268 8296 18320 8305
rect 23420 8296 23472 8348
rect 24248 8339 24300 8348
rect 24248 8305 24257 8339
rect 24257 8305 24291 8339
rect 24291 8305 24300 8339
rect 24248 8296 24300 8305
rect 26180 8296 26232 8348
rect 14772 8228 14824 8237
rect 15692 8228 15744 8280
rect 23512 8271 23564 8280
rect 23512 8237 23521 8271
rect 23521 8237 23555 8271
rect 23555 8237 23564 8271
rect 23512 8228 23564 8237
rect 23972 8271 24024 8280
rect 23972 8237 23981 8271
rect 23981 8237 24015 8271
rect 24015 8237 24024 8271
rect 23972 8228 24024 8237
rect 13116 8160 13168 8212
rect 23696 8160 23748 8212
rect 1708 8135 1760 8144
rect 1708 8101 1717 8135
rect 1717 8101 1751 8135
rect 1751 8101 1760 8135
rect 1708 8092 1760 8101
rect 6124 8092 6176 8144
rect 12932 8092 12984 8144
rect 17808 8135 17860 8144
rect 17808 8101 17817 8135
rect 17817 8101 17851 8135
rect 17851 8101 17860 8135
rect 17808 8092 17860 8101
rect 18636 8092 18688 8144
rect 18820 8135 18872 8144
rect 18820 8101 18829 8135
rect 18829 8101 18863 8135
rect 18863 8101 18872 8135
rect 18820 8092 18872 8101
rect 26272 8092 26324 8144
rect 3510 7990 3562 8042
rect 3574 7990 3626 8042
rect 3638 7990 3690 8042
rect 3702 7990 3754 8042
rect 3766 7990 3818 8042
rect 1524 7888 1576 7940
rect 1708 7888 1760 7940
rect 4192 7931 4244 7940
rect 4192 7897 4201 7931
rect 4201 7897 4235 7931
rect 4235 7897 4244 7931
rect 4192 7888 4244 7897
rect 4376 7931 4428 7940
rect 4376 7897 4385 7931
rect 4385 7897 4419 7931
rect 4419 7897 4428 7931
rect 4376 7888 4428 7897
rect 5756 7931 5808 7940
rect 5756 7897 5765 7931
rect 5765 7897 5799 7931
rect 5799 7897 5808 7931
rect 5756 7888 5808 7897
rect 6124 7931 6176 7940
rect 6124 7897 6133 7931
rect 6133 7897 6167 7931
rect 6167 7897 6176 7931
rect 6124 7888 6176 7897
rect 9068 7931 9120 7940
rect 9068 7897 9077 7931
rect 9077 7897 9111 7931
rect 9111 7897 9120 7931
rect 9068 7888 9120 7897
rect 11460 7888 11512 7940
rect 12012 7888 12064 7940
rect 13392 7888 13444 7940
rect 15232 7931 15284 7940
rect 15232 7897 15241 7931
rect 15241 7897 15275 7931
rect 15275 7897 15284 7931
rect 15232 7888 15284 7897
rect 17808 7888 17860 7940
rect 20936 7931 20988 7940
rect 20936 7897 20945 7931
rect 20945 7897 20979 7931
rect 20979 7897 20988 7931
rect 20936 7888 20988 7897
rect 21488 7931 21540 7940
rect 21488 7897 21497 7931
rect 21497 7897 21531 7931
rect 21531 7897 21540 7931
rect 21488 7888 21540 7897
rect 23420 7888 23472 7940
rect 23696 7931 23748 7940
rect 23696 7897 23705 7931
rect 23705 7897 23739 7931
rect 23739 7897 23748 7931
rect 23696 7888 23748 7897
rect 23972 7931 24024 7940
rect 23972 7897 23981 7931
rect 23981 7897 24015 7931
rect 24015 7897 24024 7931
rect 23972 7888 24024 7897
rect 26272 7931 26324 7940
rect 26272 7897 26281 7931
rect 26281 7897 26315 7931
rect 26315 7897 26324 7931
rect 26272 7888 26324 7897
rect 8976 7820 9028 7872
rect 15600 7820 15652 7872
rect 1616 7752 1668 7804
rect 12932 7795 12984 7804
rect 12932 7761 12941 7795
rect 12941 7761 12975 7795
rect 12975 7761 12984 7795
rect 12932 7752 12984 7761
rect 13484 7752 13536 7804
rect 17624 7752 17676 7804
rect 18360 7752 18412 7804
rect 18820 7752 18872 7804
rect 20016 7752 20068 7804
rect 12564 7616 12616 7668
rect 13024 7727 13076 7736
rect 13024 7693 13033 7727
rect 13033 7693 13067 7727
rect 13067 7693 13076 7727
rect 13392 7727 13444 7736
rect 13024 7684 13076 7693
rect 13392 7693 13401 7727
rect 13401 7693 13435 7727
rect 13435 7693 13444 7727
rect 13392 7684 13444 7693
rect 15876 7727 15928 7736
rect 15876 7693 15885 7727
rect 15885 7693 15919 7727
rect 15919 7693 15928 7727
rect 15876 7684 15928 7693
rect 18452 7727 18504 7736
rect 18452 7693 18461 7727
rect 18461 7693 18495 7727
rect 18495 7693 18504 7727
rect 18452 7684 18504 7693
rect 18636 7727 18688 7736
rect 18636 7693 18645 7727
rect 18645 7693 18679 7727
rect 18679 7693 18688 7727
rect 18636 7684 18688 7693
rect 19464 7727 19516 7736
rect 14772 7616 14824 7668
rect 15784 7659 15836 7668
rect 15784 7625 15793 7659
rect 15793 7625 15827 7659
rect 15827 7625 15836 7659
rect 15784 7616 15836 7625
rect 17900 7659 17952 7668
rect 17900 7625 17909 7659
rect 17909 7625 17943 7659
rect 17943 7625 17952 7659
rect 17900 7616 17952 7625
rect 18084 7616 18136 7668
rect 19464 7693 19473 7727
rect 19473 7693 19507 7727
rect 19507 7693 19516 7727
rect 19464 7684 19516 7693
rect 21488 7684 21540 7736
rect 23880 7684 23932 7736
rect 24892 7616 24944 7668
rect 26180 7659 26232 7668
rect 26180 7625 26189 7659
rect 26189 7625 26223 7659
rect 26223 7625 26232 7659
rect 26180 7616 26232 7625
rect 11368 7548 11420 7600
rect 14864 7591 14916 7600
rect 14864 7557 14873 7591
rect 14873 7557 14907 7591
rect 14907 7557 14916 7591
rect 14864 7548 14916 7557
rect 15692 7548 15744 7600
rect 17532 7591 17584 7600
rect 17532 7557 17541 7591
rect 17541 7557 17575 7591
rect 17575 7557 17584 7591
rect 17532 7548 17584 7557
rect 17624 7548 17676 7600
rect 19464 7548 19516 7600
rect 23512 7591 23564 7600
rect 23512 7557 23521 7591
rect 23521 7557 23555 7591
rect 23555 7557 23564 7591
rect 23512 7548 23564 7557
rect 24248 7548 24300 7600
rect 18870 7446 18922 7498
rect 18934 7446 18986 7498
rect 18998 7446 19050 7498
rect 19062 7446 19114 7498
rect 19126 7446 19178 7498
rect 880 7208 932 7260
rect 1340 7208 1392 7260
rect 5848 7208 5900 7260
rect 6584 7276 6636 7328
rect 8424 7276 8476 7328
rect 9896 7344 9948 7396
rect 13024 7344 13076 7396
rect 15600 7344 15652 7396
rect 17716 7387 17768 7396
rect 17716 7353 17725 7387
rect 17725 7353 17759 7387
rect 17759 7353 17768 7387
rect 17716 7344 17768 7353
rect 18084 7387 18136 7396
rect 18084 7353 18093 7387
rect 18093 7353 18127 7387
rect 18127 7353 18136 7387
rect 18084 7344 18136 7353
rect 19464 7344 19516 7396
rect 21304 7344 21356 7396
rect 23880 7344 23932 7396
rect 26180 7344 26232 7396
rect 12564 7319 12616 7328
rect 12564 7285 12573 7319
rect 12573 7285 12607 7319
rect 12607 7285 12616 7319
rect 12564 7276 12616 7285
rect 6676 7251 6728 7260
rect 6676 7217 6685 7251
rect 6685 7217 6719 7251
rect 6719 7217 6728 7251
rect 6676 7208 6728 7217
rect 8884 7208 8936 7260
rect 9620 7251 9672 7260
rect 9620 7217 9629 7251
rect 9629 7217 9663 7251
rect 9663 7217 9672 7251
rect 9620 7208 9672 7217
rect 9896 7251 9948 7260
rect 9896 7217 9905 7251
rect 9905 7217 9939 7251
rect 9939 7217 9948 7251
rect 9896 7208 9948 7217
rect 11184 7208 11236 7260
rect 12840 7251 12892 7260
rect 12840 7217 12849 7251
rect 12849 7217 12883 7251
rect 12883 7217 12892 7251
rect 12840 7208 12892 7217
rect 14220 7208 14272 7260
rect 17440 7276 17492 7328
rect 16152 7251 16204 7260
rect 16152 7217 16161 7251
rect 16161 7217 16195 7251
rect 16195 7217 16204 7251
rect 16152 7208 16204 7217
rect 972 7140 1024 7192
rect 3364 7140 3416 7192
rect 9528 7140 9580 7192
rect 10080 7183 10132 7192
rect 10080 7149 10089 7183
rect 10089 7149 10123 7183
rect 10123 7149 10132 7183
rect 10080 7140 10132 7149
rect 12748 7183 12800 7192
rect 2076 7115 2128 7124
rect 2076 7081 2085 7115
rect 2085 7081 2119 7115
rect 2119 7081 2128 7115
rect 2076 7072 2128 7081
rect 6584 7072 6636 7124
rect 9252 7072 9304 7124
rect 12748 7149 12757 7183
rect 12757 7149 12791 7183
rect 12791 7149 12800 7183
rect 12748 7140 12800 7149
rect 15692 7183 15744 7192
rect 15692 7149 15701 7183
rect 15701 7149 15735 7183
rect 15735 7149 15744 7183
rect 17624 7208 17676 7260
rect 24892 7276 24944 7328
rect 15692 7140 15744 7149
rect 17532 7140 17584 7192
rect 18268 7183 18320 7192
rect 18268 7149 18277 7183
rect 18277 7149 18311 7183
rect 18311 7149 18320 7183
rect 18268 7140 18320 7149
rect 18636 7140 18688 7192
rect 18176 7072 18228 7124
rect 19648 7208 19700 7260
rect 20016 7208 20068 7260
rect 19280 7183 19332 7192
rect 19280 7149 19289 7183
rect 19289 7149 19323 7183
rect 19323 7149 19332 7183
rect 19280 7140 19332 7149
rect 20108 7140 20160 7192
rect 20384 7072 20436 7124
rect 11368 7047 11420 7056
rect 11368 7013 11377 7047
rect 11377 7013 11411 7047
rect 11411 7013 11420 7047
rect 11368 7004 11420 7013
rect 13116 7004 13168 7056
rect 15048 7047 15100 7056
rect 15048 7013 15057 7047
rect 15057 7013 15091 7047
rect 15091 7013 15100 7047
rect 15048 7004 15100 7013
rect 19648 7004 19700 7056
rect 22040 7208 22092 7260
rect 21672 7047 21724 7056
rect 21672 7013 21681 7047
rect 21681 7013 21715 7047
rect 21715 7013 21724 7047
rect 21672 7004 21724 7013
rect 3510 6902 3562 6954
rect 3574 6902 3626 6954
rect 3638 6902 3690 6954
rect 3702 6902 3754 6954
rect 3766 6902 3818 6954
rect 972 6843 1024 6852
rect 972 6809 981 6843
rect 981 6809 1015 6843
rect 1015 6809 1024 6843
rect 972 6800 1024 6809
rect 1340 6843 1392 6852
rect 1340 6809 1349 6843
rect 1349 6809 1383 6843
rect 1383 6809 1392 6843
rect 1340 6800 1392 6809
rect 5848 6800 5900 6852
rect 6676 6800 6728 6852
rect 8608 6843 8660 6852
rect 8608 6809 8617 6843
rect 8617 6809 8651 6843
rect 8651 6809 8660 6843
rect 8608 6800 8660 6809
rect 8884 6843 8936 6852
rect 8884 6809 8893 6843
rect 8893 6809 8927 6843
rect 8927 6809 8936 6843
rect 8884 6800 8936 6809
rect 9252 6843 9304 6852
rect 9252 6809 9261 6843
rect 9261 6809 9295 6843
rect 9295 6809 9304 6843
rect 9252 6800 9304 6809
rect 9528 6843 9580 6852
rect 9528 6809 9537 6843
rect 9537 6809 9571 6843
rect 9571 6809 9580 6843
rect 9528 6800 9580 6809
rect 10356 6800 10408 6852
rect 12564 6800 12616 6852
rect 13116 6843 13168 6852
rect 13116 6809 13125 6843
rect 13125 6809 13159 6843
rect 13159 6809 13168 6843
rect 13116 6800 13168 6809
rect 14496 6800 14548 6852
rect 16152 6800 16204 6852
rect 6492 6732 6544 6784
rect 9620 6732 9672 6784
rect 11184 6732 11236 6784
rect 15600 6732 15652 6784
rect 15692 6732 15744 6784
rect 10080 6664 10132 6716
rect 16060 6664 16112 6716
rect 17992 6732 18044 6784
rect 19280 6800 19332 6852
rect 20016 6800 20068 6852
rect 22040 6843 22092 6852
rect 22040 6809 22049 6843
rect 22049 6809 22083 6843
rect 22083 6809 22092 6843
rect 22040 6800 22092 6809
rect 21212 6732 21264 6784
rect 1340 6596 1392 6648
rect 2076 6639 2128 6648
rect 2076 6605 2085 6639
rect 2085 6605 2119 6639
rect 2119 6605 2128 6639
rect 2076 6596 2128 6605
rect 6032 6596 6084 6648
rect 7320 6639 7372 6648
rect 7320 6605 7329 6639
rect 7329 6605 7363 6639
rect 7363 6605 7372 6639
rect 7320 6596 7372 6605
rect 8608 6596 8660 6648
rect 9896 6639 9948 6648
rect 9896 6605 9905 6639
rect 9905 6605 9939 6639
rect 9939 6605 9948 6639
rect 10724 6639 10776 6648
rect 9896 6596 9948 6605
rect 10724 6605 10733 6639
rect 10733 6605 10767 6639
rect 10767 6605 10776 6639
rect 10724 6596 10776 6605
rect 12840 6596 12892 6648
rect 2352 6571 2404 6580
rect 2352 6537 2361 6571
rect 2361 6537 2395 6571
rect 2395 6537 2404 6571
rect 2352 6528 2404 6537
rect 2996 6528 3048 6580
rect 6584 6528 6636 6580
rect 7228 6460 7280 6512
rect 9804 6528 9856 6580
rect 14864 6571 14916 6580
rect 14864 6537 14873 6571
rect 14873 6537 14907 6571
rect 14907 6537 14916 6571
rect 14864 6528 14916 6537
rect 15140 6639 15192 6648
rect 15140 6605 15149 6639
rect 15149 6605 15183 6639
rect 15183 6605 15192 6639
rect 15140 6596 15192 6605
rect 15692 6596 15744 6648
rect 21304 6664 21356 6716
rect 23512 6664 23564 6716
rect 15232 6528 15284 6580
rect 15784 6528 15836 6580
rect 16152 6528 16204 6580
rect 10356 6460 10408 6512
rect 11368 6503 11420 6512
rect 11368 6469 11377 6503
rect 11377 6469 11411 6503
rect 11411 6469 11420 6503
rect 12748 6503 12800 6512
rect 11368 6460 11420 6469
rect 12748 6469 12757 6503
rect 12757 6469 12791 6503
rect 12791 6469 12800 6503
rect 12748 6460 12800 6469
rect 14220 6503 14272 6512
rect 14220 6469 14229 6503
rect 14229 6469 14263 6503
rect 14263 6469 14272 6503
rect 14220 6460 14272 6469
rect 15140 6460 15192 6512
rect 17440 6503 17492 6512
rect 17440 6469 17449 6503
rect 17449 6469 17483 6503
rect 17483 6469 17492 6503
rect 17440 6460 17492 6469
rect 18544 6596 18596 6648
rect 20936 6639 20988 6648
rect 20936 6605 20945 6639
rect 20945 6605 20979 6639
rect 20979 6605 20988 6639
rect 20936 6596 20988 6605
rect 21672 6639 21724 6648
rect 20108 6571 20160 6580
rect 20108 6537 20117 6571
rect 20117 6537 20151 6571
rect 20151 6537 20160 6571
rect 20108 6528 20160 6537
rect 21672 6605 21681 6639
rect 21681 6605 21715 6639
rect 21715 6605 21724 6639
rect 21672 6596 21724 6605
rect 22316 6528 22368 6580
rect 24892 6664 24944 6716
rect 25076 6596 25128 6648
rect 19648 6503 19700 6512
rect 19648 6469 19657 6503
rect 19657 6469 19691 6503
rect 19691 6469 19700 6503
rect 19648 6460 19700 6469
rect 24616 6503 24668 6512
rect 24616 6469 24625 6503
rect 24625 6469 24659 6503
rect 24659 6469 24668 6503
rect 24616 6460 24668 6469
rect 18870 6358 18922 6410
rect 18934 6358 18986 6410
rect 18998 6358 19050 6410
rect 19062 6358 19114 6410
rect 19126 6358 19178 6410
rect 1156 6256 1208 6308
rect 1708 6256 1760 6308
rect 2076 6256 2128 6308
rect 3364 6299 3416 6308
rect 3364 6265 3373 6299
rect 3373 6265 3407 6299
rect 3407 6265 3416 6299
rect 3364 6256 3416 6265
rect 10356 6299 10408 6308
rect 10356 6265 10365 6299
rect 10365 6265 10399 6299
rect 10399 6265 10408 6299
rect 10356 6256 10408 6265
rect 11184 6256 11236 6308
rect 12840 6256 12892 6308
rect 15048 6256 15100 6308
rect 19648 6256 19700 6308
rect 20936 6299 20988 6308
rect 20936 6265 20945 6299
rect 20945 6265 20979 6299
rect 20979 6265 20988 6299
rect 20936 6256 20988 6265
rect 880 6188 932 6240
rect 6584 6188 6636 6240
rect 12288 6188 12340 6240
rect 14220 6188 14272 6240
rect 14588 6231 14640 6240
rect 14588 6197 14597 6231
rect 14597 6197 14631 6231
rect 14631 6197 14640 6231
rect 14588 6188 14640 6197
rect 15232 6231 15284 6240
rect 15232 6197 15241 6231
rect 15241 6197 15275 6231
rect 15275 6197 15284 6231
rect 15232 6188 15284 6197
rect 18636 6231 18688 6240
rect 18636 6197 18645 6231
rect 18645 6197 18679 6231
rect 18679 6197 18688 6231
rect 18636 6188 18688 6197
rect 1248 6052 1300 6104
rect 2352 6120 2404 6172
rect 3272 6120 3324 6172
rect 5664 6120 5716 6172
rect 6400 6163 6452 6172
rect 6400 6129 6409 6163
rect 6409 6129 6443 6163
rect 6443 6129 6452 6163
rect 6400 6120 6452 6129
rect 7136 6163 7188 6172
rect 7136 6129 7145 6163
rect 7145 6129 7179 6163
rect 7179 6129 7188 6163
rect 7136 6120 7188 6129
rect 7320 6163 7372 6172
rect 7320 6129 7329 6163
rect 7329 6129 7363 6163
rect 7363 6129 7372 6163
rect 7320 6120 7372 6129
rect 8976 6120 9028 6172
rect 10724 6120 10776 6172
rect 14772 6163 14824 6172
rect 14772 6129 14781 6163
rect 14781 6129 14815 6163
rect 14815 6129 14824 6163
rect 14772 6120 14824 6129
rect 16060 6163 16112 6172
rect 16060 6129 16069 6163
rect 16069 6129 16103 6163
rect 16103 6129 16112 6163
rect 16060 6120 16112 6129
rect 17624 6163 17676 6172
rect 17624 6129 17633 6163
rect 17633 6129 17667 6163
rect 17667 6129 17676 6163
rect 20292 6188 20344 6240
rect 21672 6188 21724 6240
rect 20384 6163 20436 6172
rect 17624 6120 17676 6129
rect 20384 6129 20393 6163
rect 20393 6129 20427 6163
rect 20427 6129 20436 6163
rect 20384 6120 20436 6129
rect 22500 6120 22552 6172
rect 24248 6163 24300 6172
rect 24248 6129 24257 6163
rect 24257 6129 24291 6163
rect 24291 6129 24300 6163
rect 24248 6120 24300 6129
rect 1800 6052 1852 6104
rect 4836 6095 4888 6104
rect 4836 6061 4845 6095
rect 4845 6061 4879 6095
rect 4879 6061 4888 6095
rect 4836 6052 4888 6061
rect 5388 6095 5440 6104
rect 5388 6061 5397 6095
rect 5397 6061 5431 6095
rect 5431 6061 5440 6095
rect 5388 6052 5440 6061
rect 9804 6052 9856 6104
rect 12380 5984 12432 6036
rect 15232 6052 15284 6104
rect 15968 6095 16020 6104
rect 15968 6061 15977 6095
rect 15977 6061 16011 6095
rect 16011 6061 16020 6095
rect 15968 6052 16020 6061
rect 16520 6052 16572 6104
rect 17808 6095 17860 6104
rect 17808 6061 17814 6095
rect 17814 6061 17860 6095
rect 17808 6052 17860 6061
rect 17992 6095 18044 6104
rect 17992 6061 18001 6095
rect 18001 6061 18035 6095
rect 18035 6061 18044 6095
rect 17992 6052 18044 6061
rect 18176 6052 18228 6104
rect 22592 6052 22644 6104
rect 23420 6052 23472 6104
rect 24616 6120 24668 6172
rect 25904 6120 25956 6172
rect 17440 5984 17492 6036
rect 24616 5984 24668 6036
rect 4192 5959 4244 5968
rect 4192 5925 4201 5959
rect 4201 5925 4235 5959
rect 4235 5925 4244 5959
rect 4192 5916 4244 5925
rect 8700 5959 8752 5968
rect 8700 5925 8709 5959
rect 8709 5925 8743 5959
rect 8743 5925 8752 5959
rect 8700 5916 8752 5925
rect 16244 5959 16296 5968
rect 16244 5925 16253 5959
rect 16253 5925 16287 5959
rect 16287 5925 16296 5959
rect 16244 5916 16296 5925
rect 18176 5916 18228 5968
rect 20476 5959 20528 5968
rect 20476 5925 20485 5959
rect 20485 5925 20519 5959
rect 20519 5925 20528 5959
rect 20476 5916 20528 5925
rect 22316 5916 22368 5968
rect 23788 5916 23840 5968
rect 24156 5916 24208 5968
rect 3510 5814 3562 5866
rect 3574 5814 3626 5866
rect 3638 5814 3690 5866
rect 3702 5814 3754 5866
rect 3766 5814 3818 5866
rect 880 5755 932 5764
rect 880 5721 889 5755
rect 889 5721 923 5755
rect 923 5721 932 5755
rect 880 5712 932 5721
rect 1156 5755 1208 5764
rect 1156 5721 1165 5755
rect 1165 5721 1199 5755
rect 1199 5721 1208 5755
rect 1156 5712 1208 5721
rect 3272 5712 3324 5764
rect 4836 5712 4888 5764
rect 5388 5712 5440 5764
rect 5664 5755 5716 5764
rect 5664 5721 5673 5755
rect 5673 5721 5707 5755
rect 5707 5721 5716 5755
rect 5664 5712 5716 5721
rect 6032 5712 6084 5764
rect 6400 5755 6452 5764
rect 6400 5721 6409 5755
rect 6409 5721 6443 5755
rect 6443 5721 6452 5755
rect 6400 5712 6452 5721
rect 9528 5712 9580 5764
rect 15968 5755 16020 5764
rect 15968 5721 15977 5755
rect 15977 5721 16011 5755
rect 16011 5721 16020 5755
rect 15968 5712 16020 5721
rect 16060 5712 16112 5764
rect 16244 5712 16296 5764
rect 17624 5755 17676 5764
rect 17624 5721 17633 5755
rect 17633 5721 17667 5755
rect 17667 5721 17676 5755
rect 17624 5712 17676 5721
rect 17900 5755 17952 5764
rect 17900 5721 17909 5755
rect 17909 5721 17943 5755
rect 17943 5721 17952 5755
rect 17900 5712 17952 5721
rect 20292 5755 20344 5764
rect 20292 5721 20301 5755
rect 20301 5721 20335 5755
rect 20335 5721 20344 5755
rect 20292 5712 20344 5721
rect 20476 5755 20528 5764
rect 20476 5721 20485 5755
rect 20485 5721 20519 5755
rect 20519 5721 20528 5755
rect 20476 5712 20528 5721
rect 22316 5755 22368 5764
rect 22316 5721 22325 5755
rect 22325 5721 22359 5755
rect 22359 5721 22368 5755
rect 22316 5712 22368 5721
rect 23420 5755 23472 5764
rect 23420 5721 23429 5755
rect 23429 5721 23463 5755
rect 23463 5721 23472 5755
rect 23420 5712 23472 5721
rect 24248 5712 24300 5764
rect 1800 5644 1852 5696
rect 2076 5644 2128 5696
rect 4744 5644 4796 5696
rect 2996 5619 3048 5628
rect 2996 5585 3005 5619
rect 3005 5585 3039 5619
rect 3039 5585 3048 5619
rect 2996 5576 3048 5585
rect 1064 5508 1116 5560
rect 4192 5551 4244 5560
rect 3272 5440 3324 5492
rect 4192 5517 4201 5551
rect 4201 5517 4235 5551
rect 4235 5517 4244 5551
rect 4192 5508 4244 5517
rect 4008 5440 4060 5492
rect 4468 5576 4520 5628
rect 6492 5644 6544 5696
rect 7136 5687 7188 5696
rect 7136 5653 7145 5687
rect 7145 5653 7179 5687
rect 7179 5653 7188 5687
rect 7136 5644 7188 5653
rect 14220 5687 14272 5696
rect 14220 5653 14229 5687
rect 14229 5653 14263 5687
rect 14263 5653 14272 5687
rect 14220 5644 14272 5653
rect 14772 5644 14824 5696
rect 15600 5644 15652 5696
rect 4744 5508 4796 5560
rect 6124 5576 6176 5628
rect 7228 5619 7280 5628
rect 7228 5585 7237 5619
rect 7237 5585 7271 5619
rect 7271 5585 7280 5619
rect 7228 5576 7280 5585
rect 8976 5576 9028 5628
rect 10724 5619 10776 5628
rect 10724 5585 10733 5619
rect 10733 5585 10767 5619
rect 10767 5585 10776 5619
rect 10724 5576 10776 5585
rect 23788 5687 23840 5696
rect 23788 5653 23797 5687
rect 23797 5653 23831 5687
rect 23831 5653 23840 5687
rect 23788 5644 23840 5653
rect 6308 5508 6360 5560
rect 8700 5551 8752 5560
rect 8700 5517 8709 5551
rect 8709 5517 8743 5551
rect 8743 5517 8752 5551
rect 8700 5508 8752 5517
rect 11368 5551 11420 5560
rect 11368 5517 11377 5551
rect 11377 5517 11411 5551
rect 11411 5517 11420 5551
rect 11368 5508 11420 5517
rect 12380 5551 12432 5560
rect 12380 5517 12389 5551
rect 12389 5517 12423 5551
rect 12423 5517 12432 5551
rect 12380 5508 12432 5517
rect 12748 5551 12800 5560
rect 12748 5517 12757 5551
rect 12757 5517 12791 5551
rect 12791 5517 12800 5551
rect 12748 5508 12800 5517
rect 12840 5551 12892 5560
rect 12840 5517 12849 5551
rect 12849 5517 12883 5551
rect 12883 5517 12892 5551
rect 12840 5508 12892 5517
rect 14220 5508 14272 5560
rect 14956 5551 15008 5560
rect 14956 5517 14965 5551
rect 14965 5517 14999 5551
rect 14999 5517 15008 5551
rect 14956 5508 15008 5517
rect 15140 5551 15192 5560
rect 15140 5517 15149 5551
rect 15149 5517 15183 5551
rect 15183 5517 15192 5551
rect 15140 5508 15192 5517
rect 18360 5576 18412 5628
rect 20384 5576 20436 5628
rect 23880 5619 23932 5628
rect 23880 5585 23889 5619
rect 23889 5585 23923 5619
rect 23923 5585 23932 5619
rect 23880 5576 23932 5585
rect 24156 5619 24208 5628
rect 24156 5585 24165 5619
rect 24165 5585 24199 5619
rect 24199 5585 24208 5619
rect 24156 5576 24208 5585
rect 25904 5619 25956 5628
rect 25904 5585 25913 5619
rect 25913 5585 25947 5619
rect 25947 5585 25956 5619
rect 25904 5576 25956 5585
rect 15600 5551 15652 5560
rect 15600 5517 15609 5551
rect 15609 5517 15643 5551
rect 15643 5517 15652 5551
rect 15600 5508 15652 5517
rect 15876 5508 15928 5560
rect 17440 5551 17492 5560
rect 17440 5517 17449 5551
rect 17449 5517 17483 5551
rect 17483 5517 17492 5551
rect 17440 5508 17492 5517
rect 17992 5551 18044 5560
rect 17992 5517 18001 5551
rect 18001 5517 18035 5551
rect 18035 5517 18044 5551
rect 17992 5508 18044 5517
rect 19372 5508 19424 5560
rect 19832 5508 19884 5560
rect 1248 5415 1300 5424
rect 1248 5381 1257 5415
rect 1257 5381 1291 5415
rect 1291 5381 1300 5415
rect 1248 5372 1300 5381
rect 4468 5372 4520 5424
rect 8976 5483 9028 5492
rect 8976 5449 8985 5483
rect 8985 5449 9019 5483
rect 9019 5449 9028 5483
rect 8976 5440 9028 5449
rect 9436 5440 9488 5492
rect 11184 5440 11236 5492
rect 14496 5483 14548 5492
rect 14496 5449 14505 5483
rect 14505 5449 14539 5483
rect 14539 5449 14548 5483
rect 14496 5440 14548 5449
rect 17072 5483 17124 5492
rect 17072 5449 17081 5483
rect 17081 5449 17115 5483
rect 17115 5449 17124 5483
rect 17072 5440 17124 5449
rect 17900 5440 17952 5492
rect 13668 5415 13720 5424
rect 13668 5381 13677 5415
rect 13677 5381 13711 5415
rect 13711 5381 13720 5415
rect 13668 5372 13720 5381
rect 21304 5372 21356 5424
rect 21764 5372 21816 5424
rect 22500 5415 22552 5424
rect 22500 5381 22509 5415
rect 22509 5381 22543 5415
rect 22543 5381 22552 5415
rect 22500 5372 22552 5381
rect 24616 5440 24668 5492
rect 24432 5372 24484 5424
rect 25076 5372 25128 5424
rect 18870 5270 18922 5322
rect 18934 5270 18986 5322
rect 18998 5270 19050 5322
rect 19062 5270 19114 5322
rect 19126 5270 19178 5322
rect 3364 5211 3416 5220
rect 3364 5177 3373 5211
rect 3373 5177 3407 5211
rect 3407 5177 3416 5211
rect 3364 5168 3416 5177
rect 4468 5168 4520 5220
rect 6492 5211 6544 5220
rect 6492 5177 6501 5211
rect 6501 5177 6535 5211
rect 6535 5177 6544 5211
rect 6492 5168 6544 5177
rect 8608 5168 8660 5220
rect 8976 5168 9028 5220
rect 9804 5168 9856 5220
rect 10724 5168 10776 5220
rect 13668 5168 13720 5220
rect 5388 5100 5440 5152
rect 6952 5100 7004 5152
rect 9436 5100 9488 5152
rect 10356 5100 10408 5152
rect 11184 5143 11236 5152
rect 11184 5109 11193 5143
rect 11193 5109 11227 5143
rect 11227 5109 11236 5143
rect 11184 5100 11236 5109
rect 11920 5100 11972 5152
rect 12840 5100 12892 5152
rect 14588 5168 14640 5220
rect 15232 5211 15284 5220
rect 15232 5177 15241 5211
rect 15241 5177 15275 5211
rect 15275 5177 15284 5211
rect 15232 5168 15284 5177
rect 17808 5168 17860 5220
rect 18360 5211 18412 5220
rect 18360 5177 18369 5211
rect 18369 5177 18403 5211
rect 18403 5177 18412 5211
rect 23880 5211 23932 5220
rect 18360 5168 18412 5177
rect 15140 5100 15192 5152
rect 18084 5100 18136 5152
rect 6032 5032 6084 5084
rect 9068 5075 9120 5084
rect 9068 5041 9077 5075
rect 9077 5041 9111 5075
rect 9111 5041 9120 5075
rect 9068 5032 9120 5041
rect 15048 5032 15100 5084
rect 15876 5075 15928 5084
rect 15876 5041 15885 5075
rect 15885 5041 15919 5075
rect 15919 5041 15928 5075
rect 15876 5032 15928 5041
rect 23880 5177 23889 5211
rect 23889 5177 23923 5211
rect 23923 5177 23932 5211
rect 23880 5168 23932 5177
rect 24156 5168 24208 5220
rect 18820 5100 18872 5152
rect 19280 5100 19332 5152
rect 21212 5100 21264 5152
rect 21764 5100 21816 5152
rect 24616 5100 24668 5152
rect 18912 5032 18964 5084
rect 24432 5075 24484 5084
rect 24432 5041 24441 5075
rect 24441 5041 24475 5075
rect 24475 5041 24484 5075
rect 24432 5032 24484 5041
rect 10908 5007 10960 5016
rect 10908 4973 10917 5007
rect 10917 4973 10951 5007
rect 10951 4973 10960 5007
rect 10908 4964 10960 4973
rect 15968 4964 16020 5016
rect 17992 4964 18044 5016
rect 21028 5007 21080 5016
rect 21028 4973 21037 5007
rect 21037 4973 21071 5007
rect 21071 4973 21080 5007
rect 21028 4964 21080 4973
rect 22500 4964 22552 5016
rect 5664 4939 5716 4948
rect 5664 4905 5673 4939
rect 5673 4905 5707 4939
rect 5707 4905 5716 4939
rect 5664 4896 5716 4905
rect 18820 4896 18872 4948
rect 2444 4871 2496 4880
rect 2444 4837 2453 4871
rect 2453 4837 2487 4871
rect 2487 4837 2496 4871
rect 2444 4828 2496 4837
rect 14588 4828 14640 4880
rect 16152 4828 16204 4880
rect 3510 4726 3562 4778
rect 3574 4726 3626 4778
rect 3638 4726 3690 4778
rect 3702 4726 3754 4778
rect 3766 4726 3818 4778
rect 2352 4624 2404 4676
rect 4468 4667 4520 4676
rect 4468 4633 4477 4667
rect 4477 4633 4511 4667
rect 4511 4633 4520 4667
rect 4468 4624 4520 4633
rect 6032 4624 6084 4676
rect 6492 4624 6544 4676
rect 6952 4667 7004 4676
rect 6952 4633 6961 4667
rect 6961 4633 6995 4667
rect 6995 4633 7004 4667
rect 6952 4624 7004 4633
rect 9436 4624 9488 4676
rect 11184 4624 11236 4676
rect 12748 4624 12800 4676
rect 15140 4624 15192 4676
rect 15876 4624 15928 4676
rect 16152 4667 16204 4676
rect 16152 4633 16161 4667
rect 16161 4633 16195 4667
rect 16195 4633 16204 4667
rect 16152 4624 16204 4633
rect 18728 4667 18780 4676
rect 18728 4633 18737 4667
rect 18737 4633 18771 4667
rect 18771 4633 18780 4667
rect 18728 4624 18780 4633
rect 18820 4624 18872 4676
rect 19372 4624 19424 4676
rect 21304 4667 21356 4676
rect 21304 4633 21313 4667
rect 21313 4633 21347 4667
rect 21347 4633 21356 4667
rect 21304 4624 21356 4633
rect 22500 4624 22552 4676
rect 24432 4667 24484 4676
rect 24432 4633 24441 4667
rect 24441 4633 24475 4667
rect 24475 4633 24484 4667
rect 24432 4624 24484 4633
rect 24616 4667 24668 4676
rect 24616 4633 24625 4667
rect 24625 4633 24659 4667
rect 24659 4633 24668 4667
rect 24616 4624 24668 4633
rect 12840 4556 12892 4608
rect 15048 4556 15100 4608
rect 18912 4599 18964 4608
rect 18912 4565 18921 4599
rect 18921 4565 18955 4599
rect 18955 4565 18964 4599
rect 18912 4556 18964 4565
rect 19832 4599 19884 4608
rect 2444 4463 2496 4472
rect 2444 4429 2453 4463
rect 2453 4429 2487 4463
rect 2487 4429 2496 4463
rect 2444 4420 2496 4429
rect 6124 4488 6176 4540
rect 10172 4488 10224 4540
rect 11920 4488 11972 4540
rect 15968 4488 16020 4540
rect 18728 4488 18780 4540
rect 12380 4420 12432 4472
rect 17900 4420 17952 4472
rect 19832 4565 19841 4599
rect 19841 4565 19875 4599
rect 19875 4565 19884 4599
rect 19832 4556 19884 4565
rect 21028 4556 21080 4608
rect 23880 4556 23932 4608
rect 21304 4488 21356 4540
rect 4008 4395 4060 4404
rect 4008 4361 4017 4395
rect 4017 4361 4051 4395
rect 4051 4361 4060 4395
rect 4008 4352 4060 4361
rect 8700 4352 8752 4404
rect 10908 4352 10960 4404
rect 6216 4284 6268 4336
rect 9068 4327 9120 4336
rect 9068 4293 9077 4327
rect 9077 4293 9111 4327
rect 9111 4293 9120 4327
rect 9068 4284 9120 4293
rect 12380 4327 12432 4336
rect 12380 4293 12389 4327
rect 12389 4293 12423 4327
rect 12423 4293 12432 4327
rect 12380 4284 12432 4293
rect 15508 4284 15560 4336
rect 18870 4182 18922 4234
rect 18934 4182 18986 4234
rect 18998 4182 19050 4234
rect 19062 4182 19114 4234
rect 19126 4182 19178 4234
rect 23604 4080 23656 4132
rect 25352 4080 25404 4132
rect 1340 4012 1392 4064
rect 2720 4012 2772 4064
rect 3272 4012 3324 4064
rect 14496 4012 14548 4064
rect 15232 4012 15284 4064
rect 15968 4012 16020 4064
rect 22684 4012 22736 4064
rect 788 3944 840 3996
rect 1248 3944 1300 3996
rect 1524 3944 1576 3996
rect 9160 3987 9212 3996
rect 3364 3876 3416 3928
rect 9160 3953 9169 3987
rect 9169 3953 9203 3987
rect 9203 3953 9212 3987
rect 9160 3944 9212 3953
rect 22776 3987 22828 3996
rect 22776 3953 22785 3987
rect 22785 3953 22819 3987
rect 22819 3953 22828 3987
rect 22776 3944 22828 3953
rect 15508 3876 15560 3928
rect 15876 3876 15928 3928
rect 17072 3876 17124 3928
rect 2444 3808 2496 3860
rect 3916 3808 3968 3860
rect 9160 3783 9212 3792
rect 9160 3749 9169 3783
rect 9169 3749 9203 3783
rect 9203 3749 9212 3783
rect 9160 3740 9212 3749
rect 22500 3740 22552 3792
rect 23880 3783 23932 3792
rect 23880 3749 23889 3783
rect 23889 3749 23923 3783
rect 23923 3749 23932 3783
rect 23880 3740 23932 3749
rect 24340 3740 24392 3792
rect 3510 3638 3562 3690
rect 3574 3638 3626 3690
rect 3638 3638 3690 3690
rect 3702 3638 3754 3690
rect 3766 3638 3818 3690
rect 788 3579 840 3588
rect 788 3545 797 3579
rect 797 3545 831 3579
rect 831 3545 840 3579
rect 788 3536 840 3545
rect 3272 3536 3324 3588
rect 3916 3536 3968 3588
rect 4008 3536 4060 3588
rect 1340 3511 1392 3520
rect 1340 3477 1349 3511
rect 1349 3477 1383 3511
rect 1383 3477 1392 3511
rect 1340 3468 1392 3477
rect 8700 3536 8752 3588
rect 15232 3579 15284 3588
rect 15232 3545 15241 3579
rect 15241 3545 15275 3579
rect 15275 3545 15284 3579
rect 15232 3536 15284 3545
rect 15876 3579 15928 3588
rect 15876 3545 15885 3579
rect 15885 3545 15919 3579
rect 15919 3545 15928 3579
rect 15876 3536 15928 3545
rect 21028 3579 21080 3588
rect 21028 3545 21037 3579
rect 21037 3545 21071 3579
rect 21071 3545 21080 3579
rect 21028 3536 21080 3545
rect 22500 3579 22552 3588
rect 22500 3545 22509 3579
rect 22509 3545 22543 3579
rect 22543 3545 22552 3579
rect 22500 3536 22552 3545
rect 22776 3536 22828 3588
rect 9068 3468 9120 3520
rect 15968 3468 16020 3520
rect 3364 3332 3416 3384
rect 1616 3264 1668 3316
rect 6124 3375 6176 3384
rect 6124 3341 6133 3375
rect 6133 3341 6167 3375
rect 6167 3341 6176 3375
rect 6124 3332 6176 3341
rect 23880 3536 23932 3588
rect 23880 3400 23932 3452
rect 9160 3332 9212 3384
rect 12380 3332 12432 3384
rect 17900 3375 17952 3384
rect 17900 3341 17909 3375
rect 17909 3341 17943 3375
rect 17943 3341 17952 3375
rect 17900 3332 17952 3341
rect 23604 3375 23656 3384
rect 23604 3341 23613 3375
rect 23613 3341 23647 3375
rect 23647 3341 23656 3375
rect 23604 3332 23656 3341
rect 12472 3264 12524 3316
rect 15508 3264 15560 3316
rect 17992 3264 18044 3316
rect 3272 3196 3324 3248
rect 5112 3239 5164 3248
rect 5112 3205 5121 3239
rect 5121 3205 5155 3239
rect 5155 3205 5164 3239
rect 5112 3196 5164 3205
rect 6216 3239 6268 3248
rect 6216 3205 6225 3239
rect 6225 3205 6259 3239
rect 6259 3205 6268 3239
rect 6216 3196 6268 3205
rect 11368 3196 11420 3248
rect 22684 3239 22736 3248
rect 22684 3205 22693 3239
rect 22693 3205 22727 3239
rect 22727 3205 22736 3239
rect 22684 3196 22736 3205
rect 23512 3239 23564 3248
rect 23512 3205 23521 3239
rect 23521 3205 23555 3239
rect 23555 3205 23564 3239
rect 24340 3264 24392 3316
rect 23512 3196 23564 3205
rect 18870 3094 18922 3146
rect 18934 3094 18986 3146
rect 18998 3094 19050 3146
rect 19062 3094 19114 3146
rect 19126 3094 19178 3146
rect 1340 2992 1392 3044
rect 9068 3035 9120 3044
rect 9068 3001 9077 3035
rect 9077 3001 9111 3035
rect 9111 3001 9120 3035
rect 9068 2992 9120 3001
rect 22684 2992 22736 3044
rect 24156 2992 24208 3044
rect 25260 2992 25312 3044
rect 1616 2967 1668 2976
rect 1616 2933 1625 2967
rect 1625 2933 1659 2967
rect 1659 2933 1668 2967
rect 1616 2924 1668 2933
rect 18084 2967 18136 2976
rect 18084 2933 18093 2967
rect 18093 2933 18127 2967
rect 18127 2933 18136 2967
rect 18084 2924 18136 2933
rect 20936 2924 20988 2976
rect 1432 2899 1484 2908
rect 1432 2865 1441 2899
rect 1441 2865 1475 2899
rect 1475 2865 1484 2899
rect 1432 2856 1484 2865
rect 5112 2856 5164 2908
rect 6676 2856 6728 2908
rect 10264 2856 10316 2908
rect 11828 2856 11880 2908
rect 13208 2899 13260 2908
rect 13208 2865 13217 2899
rect 13217 2865 13251 2899
rect 13251 2865 13260 2899
rect 13208 2856 13260 2865
rect 14036 2856 14088 2908
rect 14404 2856 14456 2908
rect 15968 2856 16020 2908
rect 18636 2856 18688 2908
rect 22132 2899 22184 2908
rect 1524 2788 1576 2840
rect 7504 2831 7556 2840
rect 7504 2797 7513 2831
rect 7513 2797 7547 2831
rect 7547 2797 7556 2831
rect 7504 2788 7556 2797
rect 13300 2831 13352 2840
rect 13300 2797 13309 2831
rect 13309 2797 13343 2831
rect 13343 2797 13352 2831
rect 13300 2788 13352 2797
rect 14956 2831 15008 2840
rect 14956 2797 14965 2831
rect 14965 2797 14999 2831
rect 14999 2797 15008 2831
rect 14956 2788 15008 2797
rect 17992 2831 18044 2840
rect 17992 2797 18001 2831
rect 18001 2797 18035 2831
rect 18035 2797 18044 2831
rect 17992 2788 18044 2797
rect 18176 2788 18228 2840
rect 20476 2831 20528 2840
rect 20476 2797 20485 2831
rect 20485 2797 20519 2831
rect 20519 2797 20528 2831
rect 20476 2788 20528 2797
rect 22132 2865 22141 2899
rect 22141 2865 22175 2899
rect 22175 2865 22184 2899
rect 22132 2856 22184 2865
rect 22408 2899 22460 2908
rect 22408 2865 22417 2899
rect 22417 2865 22451 2899
rect 22451 2865 22460 2899
rect 22408 2856 22460 2865
rect 23512 2899 23564 2908
rect 23512 2865 23521 2899
rect 23521 2865 23555 2899
rect 23555 2865 23564 2899
rect 23512 2856 23564 2865
rect 23880 2856 23932 2908
rect 22500 2788 22552 2840
rect 20752 2763 20804 2772
rect 4744 2652 4796 2704
rect 7136 2652 7188 2704
rect 10816 2652 10868 2704
rect 20752 2729 20761 2763
rect 20761 2729 20795 2763
rect 20795 2729 20804 2763
rect 20752 2720 20804 2729
rect 15692 2695 15744 2704
rect 15692 2661 15701 2695
rect 15701 2661 15735 2695
rect 15735 2661 15744 2695
rect 15692 2652 15744 2661
rect 22408 2652 22460 2704
rect 24064 2652 24116 2704
rect 24432 2695 24484 2704
rect 24432 2661 24441 2695
rect 24441 2661 24475 2695
rect 24475 2661 24484 2695
rect 24432 2652 24484 2661
rect 3510 2550 3562 2602
rect 3574 2550 3626 2602
rect 3638 2550 3690 2602
rect 3702 2550 3754 2602
rect 3766 2550 3818 2602
rect 1524 2448 1576 2500
rect 1432 2312 1484 2364
rect 5112 2491 5164 2500
rect 5112 2457 5121 2491
rect 5121 2457 5155 2491
rect 5155 2457 5164 2491
rect 5112 2448 5164 2457
rect 6676 2491 6728 2500
rect 6676 2457 6685 2491
rect 6685 2457 6719 2491
rect 6719 2457 6728 2491
rect 6676 2448 6728 2457
rect 11828 2491 11880 2500
rect 11828 2457 11837 2491
rect 11837 2457 11871 2491
rect 11871 2457 11880 2491
rect 11828 2448 11880 2457
rect 14404 2491 14456 2500
rect 14404 2457 14413 2491
rect 14413 2457 14447 2491
rect 14447 2457 14456 2491
rect 14404 2448 14456 2457
rect 7136 2380 7188 2432
rect 1616 2176 1668 2228
rect 13760 2380 13812 2432
rect 6676 2244 6728 2296
rect 7780 2287 7832 2296
rect 7780 2253 7789 2287
rect 7789 2253 7823 2287
rect 7823 2253 7832 2287
rect 7780 2244 7832 2253
rect 12472 2355 12524 2364
rect 12472 2321 12481 2355
rect 12481 2321 12515 2355
rect 12515 2321 12524 2355
rect 12472 2312 12524 2321
rect 1340 2108 1392 2160
rect 3088 2151 3140 2160
rect 3088 2117 3097 2151
rect 3097 2117 3131 2151
rect 3131 2117 3140 2151
rect 3088 2108 3140 2117
rect 4744 2151 4796 2160
rect 4744 2117 4753 2151
rect 4753 2117 4787 2151
rect 4787 2117 4796 2151
rect 4744 2108 4796 2117
rect 6216 2151 6268 2160
rect 6216 2117 6225 2151
rect 6225 2117 6259 2151
rect 6259 2117 6268 2151
rect 6216 2108 6268 2117
rect 9804 2151 9856 2160
rect 9804 2117 9813 2151
rect 9813 2117 9847 2151
rect 9847 2117 9856 2151
rect 11276 2244 11328 2296
rect 10816 2219 10868 2228
rect 10816 2185 10825 2219
rect 10825 2185 10859 2219
rect 10859 2185 10868 2219
rect 10816 2176 10868 2185
rect 13300 2244 13352 2296
rect 14956 2448 15008 2500
rect 17440 2491 17492 2500
rect 17440 2457 17449 2491
rect 17449 2457 17483 2491
rect 17483 2457 17492 2491
rect 17440 2448 17492 2457
rect 18084 2448 18136 2500
rect 22132 2491 22184 2500
rect 22132 2457 22141 2491
rect 22141 2457 22175 2491
rect 22175 2457 22184 2491
rect 22132 2448 22184 2457
rect 22500 2448 22552 2500
rect 23604 2448 23656 2500
rect 22408 2380 22460 2432
rect 18636 2312 18688 2364
rect 20752 2312 20804 2364
rect 21120 2312 21172 2364
rect 16520 2287 16572 2296
rect 9804 2108 9856 2117
rect 10908 2108 10960 2160
rect 15508 2176 15560 2228
rect 16520 2253 16529 2287
rect 16529 2253 16563 2287
rect 16563 2253 16572 2287
rect 16520 2244 16572 2253
rect 17900 2244 17952 2296
rect 19556 2244 19608 2296
rect 21028 2244 21080 2296
rect 16704 2176 16756 2228
rect 17440 2176 17492 2228
rect 18176 2176 18228 2228
rect 19280 2176 19332 2228
rect 24156 2355 24208 2364
rect 24156 2321 24165 2355
rect 24165 2321 24199 2355
rect 24199 2321 24208 2355
rect 24156 2312 24208 2321
rect 24432 2448 24484 2500
rect 20936 2108 20988 2160
rect 23880 2176 23932 2228
rect 24340 2176 24392 2228
rect 24892 2176 24944 2228
rect 23420 2108 23472 2160
rect 23512 2151 23564 2160
rect 23512 2117 23521 2151
rect 23521 2117 23555 2151
rect 23555 2117 23564 2151
rect 23512 2108 23564 2117
rect 18870 2006 18922 2058
rect 18934 2006 18986 2058
rect 18998 2006 19050 2058
rect 19062 2006 19114 2058
rect 19126 2006 19178 2058
rect 7504 1904 7556 1956
rect 10816 1904 10868 1956
rect 12196 1904 12248 1956
rect 13208 1904 13260 1956
rect 17992 1904 18044 1956
rect 4192 1836 4244 1888
rect 1340 1768 1392 1820
rect 2076 1768 2128 1820
rect 2536 1768 2588 1820
rect 3364 1768 3416 1820
rect 6216 1836 6268 1888
rect 7136 1879 7188 1888
rect 5848 1811 5900 1820
rect 5848 1777 5857 1811
rect 5857 1777 5891 1811
rect 5891 1777 5900 1811
rect 5848 1768 5900 1777
rect 6584 1811 6636 1820
rect 6584 1777 6593 1811
rect 6593 1777 6627 1811
rect 6627 1777 6636 1811
rect 6584 1768 6636 1777
rect 7136 1845 7145 1879
rect 7145 1845 7179 1879
rect 7179 1845 7188 1879
rect 7136 1836 7188 1845
rect 8884 1836 8936 1888
rect 9804 1836 9856 1888
rect 11368 1879 11420 1888
rect 11368 1845 11377 1879
rect 11377 1845 11411 1879
rect 11411 1845 11420 1879
rect 11368 1836 11420 1845
rect 15508 1879 15560 1888
rect 15508 1845 15517 1879
rect 15517 1845 15551 1879
rect 15551 1845 15560 1879
rect 15508 1836 15560 1845
rect 15692 1879 15744 1888
rect 15692 1845 15701 1879
rect 15701 1845 15735 1879
rect 15735 1845 15744 1879
rect 15692 1836 15744 1845
rect 16704 1836 16756 1888
rect 18176 1836 18228 1888
rect 19556 1904 19608 1956
rect 20752 1904 20804 1956
rect 22132 1904 22184 1956
rect 23052 1904 23104 1956
rect 23880 1947 23932 1956
rect 23880 1913 23889 1947
rect 23889 1913 23923 1947
rect 23923 1913 23932 1947
rect 23880 1904 23932 1913
rect 24064 1904 24116 1956
rect 24340 1904 24392 1956
rect 24708 1904 24760 1956
rect 26364 1904 26416 1956
rect 19464 1836 19516 1888
rect 23236 1879 23288 1888
rect 23236 1845 23245 1879
rect 23245 1845 23279 1879
rect 23279 1845 23288 1879
rect 23236 1836 23288 1845
rect 23604 1836 23656 1888
rect 24156 1879 24208 1888
rect 24156 1845 24165 1879
rect 24165 1845 24199 1879
rect 24199 1845 24208 1879
rect 24156 1836 24208 1845
rect 7780 1811 7832 1820
rect 7780 1777 7789 1811
rect 7789 1777 7823 1811
rect 7823 1777 7832 1811
rect 7780 1768 7832 1777
rect 8148 1768 8200 1820
rect 9712 1768 9764 1820
rect 9896 1811 9948 1820
rect 9896 1777 9905 1811
rect 9905 1777 9939 1811
rect 9939 1777 9948 1811
rect 9896 1768 9948 1777
rect 10172 1768 10224 1820
rect 12288 1768 12340 1820
rect 13392 1811 13444 1820
rect 13392 1777 13401 1811
rect 13401 1777 13435 1811
rect 13435 1777 13444 1811
rect 13392 1768 13444 1777
rect 14588 1811 14640 1820
rect 14588 1777 14597 1811
rect 14597 1777 14631 1811
rect 14631 1777 14640 1811
rect 14588 1768 14640 1777
rect 15232 1811 15284 1820
rect 15232 1777 15241 1811
rect 15241 1777 15275 1811
rect 15275 1777 15284 1811
rect 15232 1768 15284 1777
rect 16520 1811 16572 1820
rect 16520 1777 16529 1811
rect 16529 1777 16563 1811
rect 16563 1777 16572 1811
rect 16520 1768 16572 1777
rect 18912 1811 18964 1820
rect 1248 1700 1300 1752
rect 2168 1700 2220 1752
rect 2352 1743 2404 1752
rect 2352 1709 2361 1743
rect 2361 1709 2395 1743
rect 2395 1709 2404 1743
rect 2352 1700 2404 1709
rect 3916 1700 3968 1752
rect 4284 1700 4336 1752
rect 9988 1743 10040 1752
rect 9988 1709 9997 1743
rect 9997 1709 10031 1743
rect 10031 1709 10040 1743
rect 9988 1700 10040 1709
rect 10908 1743 10960 1752
rect 10908 1709 10917 1743
rect 10917 1709 10951 1743
rect 10951 1709 10960 1743
rect 10908 1700 10960 1709
rect 11460 1743 11512 1752
rect 11460 1709 11469 1743
rect 11469 1709 11503 1743
rect 11503 1709 11512 1743
rect 11460 1700 11512 1709
rect 13024 1700 13076 1752
rect 13484 1743 13536 1752
rect 13484 1709 13493 1743
rect 13493 1709 13527 1743
rect 13527 1709 13536 1743
rect 13484 1700 13536 1709
rect 14404 1700 14456 1752
rect 18084 1700 18136 1752
rect 18912 1777 18921 1811
rect 18921 1777 18955 1811
rect 18955 1777 18964 1811
rect 18912 1768 18964 1777
rect 20844 1811 20896 1820
rect 20844 1777 20853 1811
rect 20853 1777 20887 1811
rect 20887 1777 20896 1811
rect 20844 1768 20896 1777
rect 23420 1811 23472 1820
rect 23420 1777 23429 1811
rect 23429 1777 23463 1811
rect 23463 1777 23472 1811
rect 23420 1768 23472 1777
rect 26272 1768 26324 1820
rect 19004 1700 19056 1752
rect 20476 1700 20528 1752
rect 21764 1743 21816 1752
rect 21764 1709 21773 1743
rect 21773 1709 21807 1743
rect 21807 1709 21816 1743
rect 21764 1700 21816 1709
rect 7596 1607 7648 1616
rect 7596 1573 7605 1607
rect 7605 1573 7639 1607
rect 7639 1573 7648 1607
rect 7596 1564 7648 1573
rect 11828 1564 11880 1616
rect 15692 1564 15744 1616
rect 16336 1607 16388 1616
rect 16336 1573 16345 1607
rect 16345 1573 16379 1607
rect 16379 1573 16388 1607
rect 16336 1564 16388 1573
rect 17900 1607 17952 1616
rect 17900 1573 17909 1607
rect 17909 1573 17943 1607
rect 17943 1573 17952 1607
rect 17900 1564 17952 1573
rect 3510 1462 3562 1514
rect 3574 1462 3626 1514
rect 3638 1462 3690 1514
rect 3702 1462 3754 1514
rect 3766 1462 3818 1514
rect 1248 1403 1300 1412
rect 1248 1369 1257 1403
rect 1257 1369 1291 1403
rect 1291 1369 1300 1403
rect 1248 1360 1300 1369
rect 2076 1403 2128 1412
rect 2076 1369 2085 1403
rect 2085 1369 2119 1403
rect 2119 1369 2128 1403
rect 2076 1360 2128 1369
rect 2352 1360 2404 1412
rect 3272 1360 3324 1412
rect 4192 1335 4244 1344
rect 4192 1301 4201 1335
rect 4201 1301 4235 1335
rect 4235 1301 4244 1335
rect 4192 1292 4244 1301
rect 420 1224 472 1276
rect 7596 1360 7648 1412
rect 7872 1360 7924 1412
rect 8884 1403 8936 1412
rect 8884 1369 8893 1403
rect 8893 1369 8927 1403
rect 8927 1369 8936 1403
rect 8884 1360 8936 1369
rect 9712 1403 9764 1412
rect 9712 1369 9721 1403
rect 9721 1369 9755 1403
rect 9755 1369 9764 1403
rect 9712 1360 9764 1369
rect 10908 1403 10960 1412
rect 10908 1369 10917 1403
rect 10917 1369 10951 1403
rect 10951 1369 10960 1403
rect 10908 1360 10960 1369
rect 11460 1360 11512 1412
rect 12196 1403 12248 1412
rect 12196 1369 12205 1403
rect 12205 1369 12239 1403
rect 12239 1369 12248 1403
rect 12196 1360 12248 1369
rect 13484 1360 13536 1412
rect 16336 1403 16388 1412
rect 1340 1199 1392 1208
rect 1340 1165 1349 1199
rect 1349 1165 1383 1199
rect 1383 1165 1392 1199
rect 1340 1156 1392 1165
rect 7504 1224 7556 1276
rect 8332 1224 8384 1276
rect 9896 1224 9948 1276
rect 3916 1156 3968 1208
rect 5848 1199 5900 1208
rect 5848 1165 5857 1199
rect 5857 1165 5891 1199
rect 5891 1165 5900 1199
rect 5848 1156 5900 1165
rect 9988 1156 10040 1208
rect 1616 1088 1668 1140
rect 3088 1088 3140 1140
rect 6584 1131 6636 1140
rect 6584 1097 6593 1131
rect 6593 1097 6627 1131
rect 6627 1097 6636 1131
rect 6584 1088 6636 1097
rect 11828 1292 11880 1344
rect 12288 1292 12340 1344
rect 13024 1335 13076 1344
rect 13024 1301 13033 1335
rect 13033 1301 13067 1335
rect 13067 1301 13076 1335
rect 13024 1292 13076 1301
rect 11368 1267 11420 1276
rect 11368 1233 11377 1267
rect 11377 1233 11411 1267
rect 11411 1233 11420 1267
rect 11368 1224 11420 1233
rect 12196 1156 12248 1208
rect 16336 1369 16345 1403
rect 16345 1369 16379 1403
rect 16379 1369 16388 1403
rect 16336 1360 16388 1369
rect 16612 1360 16664 1412
rect 19004 1403 19056 1412
rect 19004 1369 19013 1403
rect 19013 1369 19047 1403
rect 19047 1369 19056 1403
rect 19004 1360 19056 1369
rect 20844 1360 20896 1412
rect 21028 1360 21080 1412
rect 23052 1403 23104 1412
rect 23052 1369 23061 1403
rect 23061 1369 23095 1403
rect 23095 1369 23104 1403
rect 23052 1360 23104 1369
rect 23236 1403 23288 1412
rect 23236 1369 23245 1403
rect 23245 1369 23279 1403
rect 23279 1369 23288 1403
rect 23236 1360 23288 1369
rect 23420 1403 23472 1412
rect 23420 1369 23429 1403
rect 23429 1369 23463 1403
rect 23463 1369 23472 1403
rect 23420 1360 23472 1369
rect 24156 1360 24208 1412
rect 26364 1403 26416 1412
rect 26364 1369 26373 1403
rect 26373 1369 26407 1403
rect 26407 1369 26416 1403
rect 26364 1360 26416 1369
rect 15968 1335 16020 1344
rect 15968 1301 15977 1335
rect 15977 1301 16011 1335
rect 16011 1301 16020 1335
rect 15968 1292 16020 1301
rect 19464 1335 19516 1344
rect 19464 1301 19473 1335
rect 19473 1301 19507 1335
rect 19507 1301 19516 1335
rect 19464 1292 19516 1301
rect 21764 1292 21816 1344
rect 14588 1156 14640 1208
rect 18452 1224 18504 1276
rect 15232 1088 15284 1140
rect 16428 1156 16480 1208
rect 20936 1224 20988 1276
rect 16704 1088 16756 1140
rect 18912 1088 18964 1140
rect 20476 1088 20528 1140
rect 3916 1063 3968 1072
rect 3916 1029 3925 1063
rect 3925 1029 3959 1063
rect 3959 1029 3968 1063
rect 3916 1020 3968 1029
rect 4284 1020 4336 1072
rect 9896 1020 9948 1072
rect 13392 1020 13444 1072
rect 17900 1020 17952 1072
rect 18636 1063 18688 1072
rect 18636 1029 18645 1063
rect 18645 1029 18679 1063
rect 18679 1029 18688 1063
rect 18636 1020 18688 1029
rect 25628 1156 25680 1208
rect 24892 1088 24944 1140
rect 24524 1020 24576 1072
rect 26272 1063 26324 1072
rect 26272 1029 26281 1063
rect 26281 1029 26315 1063
rect 26315 1029 26324 1063
rect 26272 1020 26324 1029
rect 18870 918 18922 970
rect 18934 918 18986 970
rect 18998 918 19050 970
rect 19062 918 19114 970
rect 19126 918 19178 970
rect 1340 859 1392 868
rect 1340 825 1349 859
rect 1349 825 1383 859
rect 1383 825 1392 859
rect 1340 816 1392 825
rect 1616 859 1668 868
rect 1616 825 1625 859
rect 1625 825 1659 859
rect 1659 825 1668 859
rect 1616 816 1668 825
rect 3364 816 3416 868
rect 3824 859 3876 868
rect 3824 825 3833 859
rect 3833 825 3867 859
rect 3867 825 3876 859
rect 3824 816 3876 825
rect 3916 816 3968 868
rect 6216 816 6268 868
rect 15508 816 15560 868
rect 25628 816 25680 868
rect 16428 748 16480 800
rect 24892 748 24944 800
rect 11644 544 11696 596
rect 12380 544 12432 596
rect 3510 374 3562 426
rect 3574 374 3626 426
rect 3638 374 3690 426
rect 3702 374 3754 426
rect 3766 374 3818 426
<< metal2 >>
rect 2216 27315 2356 27735
rect 4240 27315 4380 27735
rect 6264 27315 6404 27735
rect 8288 27315 8428 27735
rect 10312 27339 10452 27735
rect 10092 27315 10452 27339
rect 12152 27315 12292 27735
rect 14176 27315 14316 27735
rect 16200 27315 16340 27735
rect 18224 27315 18364 27735
rect 20248 27315 20388 27735
rect 22272 27315 22412 27735
rect 24296 27315 24436 27735
rect 25444 27320 25496 27326
rect 878 27016 934 27025
rect 878 26951 934 26960
rect 892 24810 920 26951
rect 2168 26232 2220 26238
rect 2168 26174 2220 26180
rect 1708 26096 1760 26102
rect 1708 26038 1760 26044
rect 972 25756 1024 25762
rect 972 25698 1024 25704
rect 984 25150 1012 25698
rect 1720 25218 1748 26038
rect 2180 25830 2208 26174
rect 2168 25824 2220 25830
rect 2168 25766 2220 25772
rect 1892 25756 1944 25762
rect 1892 25698 1944 25704
rect 1708 25212 1760 25218
rect 1708 25154 1760 25160
rect 972 25144 1024 25150
rect 972 25086 1024 25092
rect 880 24804 932 24810
rect 880 24746 932 24752
rect 892 24198 920 24746
rect 880 24192 932 24198
rect 880 24134 932 24140
rect 788 24056 840 24062
rect 788 23998 840 24004
rect 800 23382 828 23998
rect 788 23376 840 23382
rect 788 23318 840 23324
rect 878 21032 934 21041
rect 878 20967 934 20976
rect 788 20248 840 20254
rect 788 20190 840 20196
rect 892 20236 920 20967
rect 984 20338 1012 25086
rect 1904 25082 1932 25698
rect 1892 25076 1944 25082
rect 1892 25018 1944 25024
rect 1904 24810 1932 25018
rect 1892 24804 1944 24810
rect 1892 24746 1944 24752
rect 2180 24742 2208 25766
rect 2168 24736 2220 24742
rect 2168 24678 2220 24684
rect 1064 24464 1116 24470
rect 1064 24406 1116 24412
rect 1076 24130 1104 24406
rect 1064 24124 1116 24130
rect 1064 24066 1116 24072
rect 1076 23586 1104 24066
rect 1524 24056 1576 24062
rect 1430 24024 1486 24033
rect 1524 23998 1576 24004
rect 1430 23959 1486 23968
rect 1064 23580 1116 23586
rect 1064 23522 1116 23528
rect 1076 23178 1104 23522
rect 1156 23376 1208 23382
rect 1156 23318 1208 23324
rect 1064 23172 1116 23178
rect 1064 23114 1116 23120
rect 1076 22974 1104 23114
rect 1064 22968 1116 22974
rect 1064 22910 1116 22916
rect 984 20310 1104 20338
rect 972 20248 1024 20254
rect 892 20208 972 20236
rect 800 19846 828 20190
rect 892 19914 920 20208
rect 972 20190 1024 20196
rect 880 19908 932 19914
rect 880 19850 932 19856
rect 788 19840 840 19846
rect 788 19782 840 19788
rect 512 19568 564 19574
rect 512 19510 564 19516
rect 524 18554 552 19510
rect 800 18826 828 19782
rect 788 18820 840 18826
rect 788 18762 840 18768
rect 880 18684 932 18690
rect 880 18626 932 18632
rect 512 18548 564 18554
rect 512 18490 564 18496
rect 524 17942 552 18490
rect 892 18486 920 18626
rect 880 18480 932 18486
rect 880 18422 932 18428
rect 892 18049 920 18422
rect 1076 18060 1104 20310
rect 878 18040 934 18049
rect 878 17975 934 17984
rect 984 18032 1104 18060
rect 512 17936 564 17942
rect 512 17878 564 17884
rect 788 17936 840 17942
rect 788 17878 840 17884
rect 524 17534 552 17878
rect 800 17602 828 17878
rect 984 17602 1012 18032
rect 1064 17936 1116 17942
rect 1064 17878 1116 17884
rect 788 17596 840 17602
rect 788 17538 840 17544
rect 972 17596 1024 17602
rect 972 17538 1024 17544
rect 512 17528 564 17534
rect 512 17470 564 17476
rect 524 9578 552 17470
rect 696 17460 748 17466
rect 696 17402 748 17408
rect 708 16854 736 17402
rect 800 16922 828 17538
rect 984 17194 1012 17538
rect 972 17188 1024 17194
rect 972 17130 1024 17136
rect 788 16916 840 16922
rect 788 16858 840 16864
rect 696 16848 748 16854
rect 696 16790 748 16796
rect 708 12065 736 16790
rect 800 16650 828 16858
rect 788 16644 840 16650
rect 788 16586 840 16592
rect 880 15352 932 15358
rect 880 15294 932 15300
rect 892 15057 920 15294
rect 878 15048 934 15057
rect 878 14983 934 14992
rect 694 12056 750 12065
rect 694 11991 750 12000
rect 512 9572 564 9578
rect 512 9514 564 9520
rect 788 9572 840 9578
rect 788 9514 840 9520
rect 694 9064 750 9073
rect 694 8999 750 9008
rect 708 8898 736 8999
rect 696 8892 748 8898
rect 696 8834 748 8840
rect 708 8490 736 8834
rect 800 8830 828 9514
rect 788 8824 840 8830
rect 788 8766 840 8772
rect 880 8756 932 8762
rect 880 8698 932 8704
rect 892 8490 920 8698
rect 696 8484 748 8490
rect 696 8426 748 8432
rect 880 8484 932 8490
rect 880 8426 932 8432
rect 892 7266 920 8426
rect 880 7260 932 7266
rect 880 7202 932 7208
rect 972 7192 1024 7198
rect 972 7134 1024 7140
rect 984 6858 1012 7134
rect 972 6852 1024 6858
rect 972 6794 1024 6800
rect 880 6240 932 6246
rect 880 6182 932 6188
rect 892 6081 920 6182
rect 878 6072 934 6081
rect 878 6007 934 6016
rect 892 5770 920 6007
rect 880 5764 932 5770
rect 880 5706 932 5712
rect 1076 5566 1104 17878
rect 1168 14406 1196 23318
rect 1248 22424 1300 22430
rect 1248 22366 1300 22372
rect 1260 21750 1288 22366
rect 1248 21744 1300 21750
rect 1248 21686 1300 21692
rect 1260 21206 1288 21686
rect 1248 21200 1300 21206
rect 1248 21142 1300 21148
rect 1260 20322 1288 21142
rect 1248 20316 1300 20322
rect 1248 20258 1300 20264
rect 1260 19914 1288 20258
rect 1248 19908 1300 19914
rect 1248 19850 1300 19856
rect 1340 19364 1392 19370
rect 1340 19306 1392 19312
rect 1352 18622 1380 19306
rect 1340 18616 1392 18622
rect 1340 18558 1392 18564
rect 1248 18548 1300 18554
rect 1248 18490 1300 18496
rect 1260 17942 1288 18490
rect 1248 17936 1300 17942
rect 1248 17878 1300 17884
rect 1248 16984 1300 16990
rect 1248 16926 1300 16932
rect 1260 16310 1288 16926
rect 1248 16304 1300 16310
rect 1248 16246 1300 16252
rect 1156 14400 1208 14406
rect 1156 14342 1208 14348
rect 1260 12842 1288 16246
rect 1340 14128 1392 14134
rect 1340 14070 1392 14076
rect 1352 13590 1380 14070
rect 1340 13584 1392 13590
rect 1340 13526 1392 13532
rect 1352 13046 1380 13526
rect 1340 13040 1392 13046
rect 1340 12982 1392 12988
rect 1248 12836 1300 12842
rect 1248 12778 1300 12784
rect 1260 12298 1288 12778
rect 1248 12292 1300 12298
rect 1248 12234 1300 12240
rect 1352 10122 1380 12982
rect 1340 10116 1392 10122
rect 1340 10058 1392 10064
rect 1340 7260 1392 7266
rect 1340 7202 1392 7208
rect 1352 6858 1380 7202
rect 1340 6852 1392 6858
rect 1340 6794 1392 6800
rect 1352 6654 1380 6794
rect 1340 6648 1392 6654
rect 1340 6590 1392 6596
rect 1156 6308 1208 6314
rect 1156 6250 1208 6256
rect 1168 5770 1196 6250
rect 1248 6104 1300 6110
rect 1248 6046 1300 6052
rect 1156 5764 1208 5770
rect 1156 5706 1208 5712
rect 1064 5560 1116 5566
rect 1064 5502 1116 5508
rect 1260 5430 1288 6046
rect 1248 5424 1300 5430
rect 1248 5366 1300 5372
rect 1260 4002 1288 5366
rect 1340 4064 1392 4070
rect 1340 4006 1392 4012
rect 788 3996 840 4002
rect 788 3938 840 3944
rect 1248 3996 1300 4002
rect 1248 3938 1300 3944
rect 800 3594 828 3938
rect 788 3588 840 3594
rect 788 3530 840 3536
rect 1352 3526 1380 4006
rect 1444 3905 1472 23959
rect 1536 20322 1564 23998
rect 2168 23988 2220 23994
rect 2168 23930 2220 23936
rect 1892 23580 1944 23586
rect 1892 23522 1944 23528
rect 1800 23512 1852 23518
rect 1800 23454 1852 23460
rect 1812 23110 1840 23454
rect 1800 23104 1852 23110
rect 1800 23046 1852 23052
rect 1812 22634 1840 23046
rect 1904 22906 1932 23522
rect 1984 23376 2036 23382
rect 1984 23318 2036 23324
rect 1996 22974 2024 23318
rect 1984 22968 2036 22974
rect 2036 22928 2116 22956
rect 1984 22910 2036 22916
rect 1892 22900 1944 22906
rect 1892 22842 1944 22848
rect 1800 22628 1852 22634
rect 1800 22570 1852 22576
rect 1904 21410 1932 22842
rect 1984 22424 2036 22430
rect 1984 22366 2036 22372
rect 1996 21546 2024 22366
rect 2088 21886 2116 22928
rect 2180 22634 2208 23930
rect 2168 22628 2220 22634
rect 2168 22570 2220 22576
rect 2180 22022 2208 22570
rect 2168 22016 2220 22022
rect 2168 21958 2220 21964
rect 2076 21880 2128 21886
rect 2076 21822 2128 21828
rect 1984 21540 2036 21546
rect 1984 21482 2036 21488
rect 1892 21404 1944 21410
rect 1892 21346 1944 21352
rect 1904 21002 1932 21346
rect 1996 21002 2024 21482
rect 2088 21478 2116 21822
rect 2076 21472 2128 21478
rect 2076 21414 2128 21420
rect 1892 20996 1944 21002
rect 1892 20938 1944 20944
rect 1984 20996 2036 21002
rect 1984 20938 2036 20944
rect 1524 20316 1576 20322
rect 1524 20258 1576 20264
rect 1536 19574 1564 20258
rect 2088 19914 2116 21414
rect 2076 19908 2128 19914
rect 2076 19850 2128 19856
rect 2272 19734 2300 27315
rect 3504 26540 3824 26560
rect 3504 26538 3516 26540
rect 3572 26538 3596 26540
rect 3652 26538 3676 26540
rect 3732 26538 3756 26540
rect 3812 26538 3824 26540
rect 3504 26486 3510 26538
rect 3572 26486 3574 26538
rect 3754 26486 3756 26538
rect 3818 26486 3824 26538
rect 3504 26484 3516 26486
rect 3572 26484 3596 26486
rect 3652 26484 3676 26486
rect 3732 26484 3756 26486
rect 3812 26484 3824 26486
rect 3504 26464 3824 26484
rect 4296 26374 4324 27315
rect 6216 26776 6268 26782
rect 6216 26718 6268 26724
rect 3916 26368 3968 26374
rect 3916 26310 3968 26316
rect 4284 26368 4336 26374
rect 4284 26310 4336 26316
rect 2996 26300 3048 26306
rect 2996 26242 3048 26248
rect 3008 25354 3036 26242
rect 3364 26232 3416 26238
rect 3364 26174 3416 26180
rect 3376 25762 3404 26174
rect 3364 25756 3416 25762
rect 3364 25698 3416 25704
rect 3376 25354 3404 25698
rect 3504 25452 3824 25472
rect 3504 25450 3516 25452
rect 3572 25450 3596 25452
rect 3652 25450 3676 25452
rect 3732 25450 3756 25452
rect 3812 25450 3824 25452
rect 3504 25398 3510 25450
rect 3572 25398 3574 25450
rect 3754 25398 3756 25450
rect 3818 25398 3824 25450
rect 3504 25396 3516 25398
rect 3572 25396 3596 25398
rect 3652 25396 3676 25398
rect 3732 25396 3756 25398
rect 3812 25396 3824 25398
rect 3504 25376 3824 25396
rect 3928 25354 3956 26310
rect 6228 26102 6256 26718
rect 4192 26096 4244 26102
rect 4192 26038 4244 26044
rect 6216 26096 6268 26102
rect 6216 26038 6268 26044
rect 4204 25626 4232 26038
rect 4284 25756 4336 25762
rect 4284 25698 4336 25704
rect 4192 25620 4244 25626
rect 4192 25562 4244 25568
rect 2996 25348 3048 25354
rect 2996 25290 3048 25296
rect 3364 25348 3416 25354
rect 3364 25290 3416 25296
rect 3916 25348 3968 25354
rect 3916 25290 3968 25296
rect 3504 24364 3824 24384
rect 3504 24362 3516 24364
rect 3572 24362 3596 24364
rect 3652 24362 3676 24364
rect 3732 24362 3756 24364
rect 3812 24362 3824 24364
rect 3504 24310 3510 24362
rect 3572 24310 3574 24362
rect 3754 24310 3756 24362
rect 3818 24310 3824 24362
rect 3504 24308 3516 24310
rect 3572 24308 3596 24310
rect 3652 24308 3676 24310
rect 3732 24308 3756 24310
rect 3812 24308 3824 24310
rect 3504 24288 3824 24308
rect 3928 24266 3956 25290
rect 4204 25082 4232 25562
rect 4296 25354 4324 25698
rect 6228 25694 6256 26038
rect 5388 25688 5440 25694
rect 5388 25630 5440 25636
rect 6216 25688 6268 25694
rect 6216 25630 6268 25636
rect 4284 25348 4336 25354
rect 4284 25290 4336 25296
rect 4192 25076 4244 25082
rect 4192 25018 4244 25024
rect 4204 24674 4232 25018
rect 5400 25014 5428 25630
rect 6228 25150 6256 25630
rect 6216 25144 6268 25150
rect 6216 25086 6268 25092
rect 5388 25008 5440 25014
rect 5388 24950 5440 24956
rect 5480 25008 5532 25014
rect 5480 24950 5532 24956
rect 4192 24668 4244 24674
rect 4192 24610 4244 24616
rect 3916 24260 3968 24266
rect 3916 24202 3968 24208
rect 4204 24198 4232 24610
rect 4284 24464 4336 24470
rect 4284 24406 4336 24412
rect 4296 24266 4324 24406
rect 4284 24260 4336 24266
rect 4284 24202 4336 24208
rect 4192 24192 4244 24198
rect 4192 24134 4244 24140
rect 4296 23586 4324 24202
rect 4192 23580 4244 23586
rect 4192 23522 4244 23528
rect 4284 23580 4336 23586
rect 4284 23522 4336 23528
rect 3504 23276 3824 23296
rect 3504 23274 3516 23276
rect 3572 23274 3596 23276
rect 3652 23274 3676 23276
rect 3732 23274 3756 23276
rect 3812 23274 3824 23276
rect 3504 23222 3510 23274
rect 3572 23222 3574 23274
rect 3754 23222 3756 23274
rect 3818 23222 3824 23274
rect 3504 23220 3516 23222
rect 3572 23220 3596 23222
rect 3652 23220 3676 23222
rect 3732 23220 3756 23222
rect 3812 23220 3824 23222
rect 3504 23200 3824 23220
rect 4204 23178 4232 23522
rect 4192 23172 4244 23178
rect 4192 23114 4244 23120
rect 4296 23110 4324 23522
rect 4284 23104 4336 23110
rect 4284 23046 4336 23052
rect 4296 22498 4324 23046
rect 5204 22900 5256 22906
rect 5204 22842 5256 22848
rect 5216 22566 5244 22842
rect 5204 22560 5256 22566
rect 5204 22502 5256 22508
rect 4284 22492 4336 22498
rect 4284 22434 4336 22440
rect 4928 22492 4980 22498
rect 4928 22434 4980 22440
rect 4008 22288 4060 22294
rect 4008 22230 4060 22236
rect 3504 22188 3824 22208
rect 3504 22186 3516 22188
rect 3572 22186 3596 22188
rect 3652 22186 3676 22188
rect 3732 22186 3756 22188
rect 3812 22186 3824 22188
rect 3504 22134 3510 22186
rect 3572 22134 3574 22186
rect 3754 22134 3756 22186
rect 3818 22134 3824 22186
rect 3504 22132 3516 22134
rect 3572 22132 3596 22134
rect 3652 22132 3676 22134
rect 3732 22132 3756 22134
rect 3812 22132 3824 22134
rect 3504 22112 3824 22132
rect 4020 22090 4048 22230
rect 4008 22084 4060 22090
rect 4008 22026 4060 22032
rect 4020 21410 4048 22026
rect 4296 22022 4324 22434
rect 4284 22016 4336 22022
rect 4284 21958 4336 21964
rect 4296 21546 4324 21958
rect 4940 21818 4968 22434
rect 5216 22090 5244 22502
rect 5204 22084 5256 22090
rect 5204 22026 5256 22032
rect 4928 21812 4980 21818
rect 4928 21754 4980 21760
rect 4560 21744 4612 21750
rect 4560 21686 4612 21692
rect 4284 21540 4336 21546
rect 4284 21482 4336 21488
rect 4008 21404 4060 21410
rect 4008 21346 4060 21352
rect 4572 21342 4600 21686
rect 4940 21478 4968 21754
rect 4928 21472 4980 21478
rect 4928 21414 4980 21420
rect 4744 21404 4796 21410
rect 4744 21346 4796 21352
rect 4560 21336 4612 21342
rect 4560 21278 4612 21284
rect 3504 21100 3824 21120
rect 3504 21098 3516 21100
rect 3572 21098 3596 21100
rect 3652 21098 3676 21100
rect 3732 21098 3756 21100
rect 3812 21098 3824 21100
rect 3504 21046 3510 21098
rect 3572 21046 3574 21098
rect 3754 21046 3756 21098
rect 3818 21046 3824 21098
rect 3504 21044 3516 21046
rect 3572 21044 3596 21046
rect 3652 21044 3676 21046
rect 3732 21044 3756 21046
rect 3812 21044 3824 21046
rect 3504 21024 3824 21044
rect 4572 20866 4600 21278
rect 4756 21002 4784 21346
rect 4940 21002 4968 21414
rect 4744 20996 4796 21002
rect 4744 20938 4796 20944
rect 4928 20996 4980 21002
rect 4928 20938 4980 20944
rect 4560 20860 4612 20866
rect 4560 20802 4612 20808
rect 4560 20316 4612 20322
rect 4560 20258 4612 20264
rect 4376 20112 4428 20118
rect 4376 20054 4428 20060
rect 3504 20012 3824 20032
rect 3504 20010 3516 20012
rect 3572 20010 3596 20012
rect 3652 20010 3676 20012
rect 3732 20010 3756 20012
rect 3812 20010 3824 20012
rect 3504 19958 3510 20010
rect 3572 19958 3574 20010
rect 3754 19958 3756 20010
rect 3818 19958 3824 20010
rect 3504 19956 3516 19958
rect 3572 19956 3596 19958
rect 3652 19956 3676 19958
rect 3732 19956 3756 19958
rect 3812 19956 3824 19958
rect 3504 19936 3824 19956
rect 4388 19778 4416 20054
rect 4376 19772 4428 19778
rect 2272 19706 2392 19734
rect 4376 19714 4428 19720
rect 1708 19636 1760 19642
rect 1708 19578 1760 19584
rect 1524 19568 1576 19574
rect 1524 19510 1576 19516
rect 1720 19370 1748 19578
rect 2260 19568 2312 19574
rect 2260 19510 2312 19516
rect 1708 19364 1760 19370
rect 1708 19306 1760 19312
rect 1708 18820 1760 18826
rect 1708 18762 1760 18768
rect 1720 17126 1748 18762
rect 1708 17120 1760 17126
rect 1760 17080 1840 17108
rect 1708 17062 1760 17068
rect 1708 16848 1760 16854
rect 1708 16790 1760 16796
rect 1616 16304 1668 16310
rect 1616 16246 1668 16252
rect 1524 12632 1576 12638
rect 1524 12574 1576 12580
rect 1536 11958 1564 12574
rect 1524 11952 1576 11958
rect 1524 11894 1576 11900
rect 1536 11414 1564 11894
rect 1628 11618 1656 16246
rect 1720 16106 1748 16790
rect 1812 16650 1840 17080
rect 1800 16644 1852 16650
rect 1800 16586 1852 16592
rect 1708 16100 1760 16106
rect 1708 16042 1760 16048
rect 1720 15494 1748 16042
rect 1812 16038 1840 16586
rect 1800 16032 1852 16038
rect 1852 15992 1932 16020
rect 1800 15974 1852 15980
rect 1800 15896 1852 15902
rect 1800 15838 1852 15844
rect 1812 15562 1840 15838
rect 1904 15562 1932 15992
rect 2076 15828 2128 15834
rect 2076 15770 2128 15776
rect 1800 15556 1852 15562
rect 1800 15498 1852 15504
rect 1892 15556 1944 15562
rect 1892 15498 1944 15504
rect 1708 15488 1760 15494
rect 1708 15430 1760 15436
rect 1982 15456 2038 15465
rect 1892 15420 1944 15426
rect 1982 15391 2038 15400
rect 1892 15362 1944 15368
rect 1708 15284 1760 15290
rect 1708 15226 1760 15232
rect 1720 15193 1748 15226
rect 1706 15184 1762 15193
rect 1706 15119 1762 15128
rect 1904 14950 1932 15362
rect 1996 15358 2024 15391
rect 1984 15352 2036 15358
rect 1984 15294 2036 15300
rect 1984 15012 2036 15018
rect 1984 14954 2036 14960
rect 1892 14944 1944 14950
rect 1892 14886 1944 14892
rect 1800 14400 1852 14406
rect 1800 14342 1852 14348
rect 1812 14270 1840 14342
rect 1800 14264 1852 14270
rect 1800 14206 1852 14212
rect 1996 14202 2024 14954
rect 1984 14196 2036 14202
rect 1984 14138 2036 14144
rect 1708 13788 1760 13794
rect 1708 13730 1760 13736
rect 1720 13046 1748 13730
rect 1892 13108 1944 13114
rect 1892 13050 1944 13056
rect 1708 13040 1760 13046
rect 1708 12982 1760 12988
rect 1720 12706 1748 12982
rect 1708 12700 1760 12706
rect 1708 12642 1760 12648
rect 1720 12298 1748 12642
rect 1708 12292 1760 12298
rect 1708 12234 1760 12240
rect 1800 11680 1852 11686
rect 1904 11668 1932 13050
rect 1852 11640 1932 11668
rect 1800 11622 1852 11628
rect 1616 11612 1668 11618
rect 1616 11554 1668 11560
rect 1524 11408 1576 11414
rect 1524 11350 1576 11356
rect 1536 10938 1564 11350
rect 1628 11210 1656 11554
rect 1812 11210 1840 11622
rect 1616 11204 1668 11210
rect 1616 11146 1668 11152
rect 1800 11204 1852 11210
rect 1800 11146 1852 11152
rect 1524 10932 1576 10938
rect 1524 10874 1576 10880
rect 1536 8354 1564 10874
rect 2088 10666 2116 15770
rect 2168 15760 2220 15766
rect 2168 15702 2220 15708
rect 2180 15018 2208 15702
rect 2168 15012 2220 15018
rect 2168 14954 2220 14960
rect 2272 14214 2300 19510
rect 2364 17641 2392 19706
rect 4572 19658 4600 20258
rect 4652 20112 4704 20118
rect 4652 20054 4704 20060
rect 4296 19630 4600 19658
rect 4192 19568 4244 19574
rect 4296 19556 4324 19630
rect 4664 19574 4692 20054
rect 5020 19840 5072 19846
rect 5020 19782 5072 19788
rect 4244 19528 4324 19556
rect 4468 19568 4520 19574
rect 4192 19510 4244 19516
rect 4468 19510 4520 19516
rect 4652 19568 4704 19574
rect 4652 19510 4704 19516
rect 3504 18924 3824 18944
rect 3504 18922 3516 18924
rect 3572 18922 3596 18924
rect 3652 18922 3676 18924
rect 3732 18922 3756 18924
rect 3812 18922 3824 18924
rect 3504 18870 3510 18922
rect 3572 18870 3574 18922
rect 3754 18870 3756 18922
rect 3818 18870 3824 18922
rect 3504 18868 3516 18870
rect 3572 18868 3596 18870
rect 3652 18868 3676 18870
rect 3732 18868 3756 18870
rect 3812 18868 3824 18870
rect 3504 18848 3824 18868
rect 3364 18616 3416 18622
rect 3364 18558 3416 18564
rect 2350 17632 2406 17641
rect 2350 17567 2406 17576
rect 3272 17596 3324 17602
rect 3272 17538 3324 17544
rect 2628 17392 2680 17398
rect 2628 17334 2680 17340
rect 2640 17194 2668 17334
rect 2628 17188 2680 17194
rect 2628 17130 2680 17136
rect 2536 16916 2588 16922
rect 2536 16858 2588 16864
rect 2548 16514 2576 16858
rect 2640 16854 2668 17130
rect 2628 16848 2680 16854
rect 2628 16790 2680 16796
rect 2536 16508 2588 16514
rect 2536 16450 2588 16456
rect 2640 16446 2668 16790
rect 3284 16650 3312 17538
rect 3272 16644 3324 16650
rect 3272 16586 3324 16592
rect 3376 16514 3404 18558
rect 3916 18276 3968 18282
rect 3916 18218 3968 18224
rect 3504 17836 3824 17856
rect 3504 17834 3516 17836
rect 3572 17834 3596 17836
rect 3652 17834 3676 17836
rect 3732 17834 3756 17836
rect 3812 17834 3824 17836
rect 3504 17782 3510 17834
rect 3572 17782 3574 17834
rect 3754 17782 3756 17834
rect 3818 17782 3824 17834
rect 3504 17780 3516 17782
rect 3572 17780 3596 17782
rect 3652 17780 3676 17782
rect 3732 17780 3756 17782
rect 3812 17780 3824 17782
rect 3504 17760 3824 17780
rect 3504 16748 3824 16768
rect 3504 16746 3516 16748
rect 3572 16746 3596 16748
rect 3652 16746 3676 16748
rect 3732 16746 3756 16748
rect 3812 16746 3824 16748
rect 3504 16694 3510 16746
rect 3572 16694 3574 16746
rect 3754 16694 3756 16746
rect 3818 16694 3824 16746
rect 3504 16692 3516 16694
rect 3572 16692 3596 16694
rect 3652 16692 3676 16694
rect 3732 16692 3756 16694
rect 3812 16692 3824 16694
rect 3504 16672 3824 16692
rect 3928 16582 3956 18218
rect 4100 18140 4152 18146
rect 4100 18082 4152 18088
rect 4008 17528 4060 17534
rect 4008 17470 4060 17476
rect 4020 17398 4048 17470
rect 4008 17392 4060 17398
rect 4008 17334 4060 17340
rect 3916 16576 3968 16582
rect 3916 16518 3968 16524
rect 3364 16508 3416 16514
rect 3364 16450 3416 16456
rect 3928 16446 3956 16518
rect 2628 16440 2680 16446
rect 2628 16382 2680 16388
rect 3272 16440 3324 16446
rect 3272 16382 3324 16388
rect 3916 16440 3968 16446
rect 3916 16382 3968 16388
rect 2996 16304 3048 16310
rect 2996 16246 3048 16252
rect 3008 15834 3036 16246
rect 2996 15828 3048 15834
rect 2996 15770 3048 15776
rect 2444 15556 2496 15562
rect 2444 15498 2496 15504
rect 2996 15556 3048 15562
rect 2996 15498 3048 15504
rect 2456 14678 2484 15498
rect 3008 15465 3036 15498
rect 2994 15456 3050 15465
rect 2628 15420 2680 15426
rect 2628 15362 2680 15368
rect 2916 15414 2994 15442
rect 2536 14944 2588 14950
rect 2536 14886 2588 14892
rect 2444 14672 2496 14678
rect 2444 14614 2496 14620
rect 2272 14186 2484 14214
rect 2260 13788 2312 13794
rect 2260 13730 2312 13736
rect 2272 13386 2300 13730
rect 2260 13380 2312 13386
rect 2260 13322 2312 13328
rect 2352 12768 2404 12774
rect 2352 12710 2404 12716
rect 2260 12496 2312 12502
rect 2260 12438 2312 12444
rect 2272 12162 2300 12438
rect 2260 12156 2312 12162
rect 2260 12098 2312 12104
rect 2168 11952 2220 11958
rect 2168 11894 2220 11900
rect 2180 11414 2208 11894
rect 2272 11482 2300 12098
rect 2260 11476 2312 11482
rect 2260 11418 2312 11424
rect 2168 11408 2220 11414
rect 2168 11350 2220 11356
rect 2076 10660 2128 10666
rect 2076 10602 2128 10608
rect 2088 9850 2116 10602
rect 2076 9844 2128 9850
rect 2076 9786 2128 9792
rect 1800 9776 1852 9782
rect 1800 9718 1852 9724
rect 1812 9578 1840 9718
rect 2088 9578 2116 9786
rect 1800 9572 1852 9578
rect 1800 9514 1852 9520
rect 2076 9572 2128 9578
rect 2076 9514 2128 9520
rect 1616 9504 1668 9510
rect 1616 9446 1668 9452
rect 1628 8830 1656 9446
rect 2088 9034 2116 9514
rect 2076 9028 2128 9034
rect 2076 8970 2128 8976
rect 1616 8824 1668 8830
rect 1668 8784 1840 8812
rect 1616 8766 1668 8772
rect 1524 8348 1576 8354
rect 1524 8290 1576 8296
rect 1616 8348 1668 8354
rect 1616 8290 1668 8296
rect 1536 7946 1564 8290
rect 1524 7940 1576 7946
rect 1524 7882 1576 7888
rect 1628 7810 1656 8290
rect 1708 8144 1760 8150
rect 1708 8086 1760 8092
rect 1720 7946 1748 8086
rect 1708 7940 1760 7946
rect 1708 7882 1760 7888
rect 1616 7804 1668 7810
rect 1616 7746 1668 7752
rect 1720 6314 1748 7882
rect 1708 6308 1760 6314
rect 1708 6250 1760 6256
rect 1812 6110 1840 8784
rect 2076 7124 2128 7130
rect 2076 7066 2128 7072
rect 2088 6654 2116 7066
rect 2076 6648 2128 6654
rect 2076 6590 2128 6596
rect 2088 6314 2116 6590
rect 2076 6308 2128 6314
rect 2076 6250 2128 6256
rect 1800 6104 1852 6110
rect 1800 6046 1852 6052
rect 1812 5702 1840 6046
rect 1800 5696 1852 5702
rect 1800 5638 1852 5644
rect 2076 5696 2128 5702
rect 2076 5638 2128 5644
rect 1524 3996 1576 4002
rect 1524 3938 1576 3944
rect 1430 3896 1486 3905
rect 1430 3831 1486 3840
rect 1340 3520 1392 3526
rect 1340 3462 1392 3468
rect 418 3080 474 3089
rect 1352 3050 1380 3462
rect 418 3015 474 3024
rect 1340 3044 1392 3050
rect 432 1865 460 3015
rect 1340 2986 1392 2992
rect 1432 2908 1484 2914
rect 1432 2850 1484 2856
rect 1444 2370 1472 2850
rect 1536 2846 1564 3938
rect 1616 3316 1668 3322
rect 1616 3258 1668 3264
rect 1628 2982 1656 3258
rect 1616 2976 1668 2982
rect 1616 2918 1668 2924
rect 1524 2840 1576 2846
rect 1524 2782 1576 2788
rect 1536 2506 1564 2782
rect 1524 2500 1576 2506
rect 1524 2442 1576 2448
rect 1432 2364 1484 2370
rect 1432 2306 1484 2312
rect 1616 2228 1668 2234
rect 1616 2170 1668 2176
rect 1340 2160 1392 2166
rect 1340 2102 1392 2108
rect 418 1856 474 1865
rect 1352 1826 1380 2102
rect 418 1791 474 1800
rect 1340 1820 1392 1826
rect 1340 1762 1392 1768
rect 1248 1752 1300 1758
rect 1248 1694 1300 1700
rect 1260 1418 1288 1694
rect 1248 1412 1300 1418
rect 1248 1354 1300 1360
rect 420 1276 472 1282
rect 420 1218 472 1224
rect 432 420 460 1218
rect 1352 1214 1380 1762
rect 1340 1208 1392 1214
rect 1340 1150 1392 1156
rect 1352 874 1380 1150
rect 1628 1146 1656 2170
rect 2088 1826 2116 5638
rect 2076 1820 2128 1826
rect 2076 1762 2128 1768
rect 2088 1418 2116 1762
rect 2180 1758 2208 11350
rect 2364 11210 2392 12710
rect 2352 11204 2404 11210
rect 2352 11146 2404 11152
rect 2364 10666 2392 11146
rect 2352 10660 2404 10666
rect 2352 10602 2404 10608
rect 2364 9442 2392 10602
rect 2456 9458 2484 14186
rect 2548 11210 2576 14886
rect 2640 14882 2668 15362
rect 2720 14944 2772 14950
rect 2720 14886 2772 14892
rect 2628 14876 2680 14882
rect 2628 14818 2680 14824
rect 2732 14338 2760 14886
rect 2812 14876 2864 14882
rect 2812 14818 2864 14824
rect 2720 14332 2772 14338
rect 2720 14274 2772 14280
rect 2732 12162 2760 14274
rect 2824 13386 2852 14818
rect 2812 13380 2864 13386
rect 2812 13322 2864 13328
rect 2720 12156 2772 12162
rect 2720 12098 2772 12104
rect 2732 11754 2760 12098
rect 2720 11748 2772 11754
rect 2720 11690 2772 11696
rect 2536 11204 2588 11210
rect 2536 11146 2588 11152
rect 2916 11074 2944 15414
rect 3284 15426 3312 16382
rect 3504 15660 3824 15680
rect 3504 15658 3516 15660
rect 3572 15658 3596 15660
rect 3652 15658 3676 15660
rect 3732 15658 3756 15660
rect 3812 15658 3824 15660
rect 3504 15606 3510 15658
rect 3572 15606 3574 15658
rect 3754 15606 3756 15658
rect 3818 15606 3824 15658
rect 3504 15604 3516 15606
rect 3572 15604 3596 15606
rect 3652 15604 3676 15606
rect 3732 15604 3756 15606
rect 3812 15604 3824 15606
rect 3504 15584 3824 15604
rect 3928 15562 3956 16382
rect 4020 15562 4048 17334
rect 4112 17194 4140 18082
rect 4204 18078 4232 19510
rect 4480 18486 4508 19510
rect 4560 19296 4612 19302
rect 4560 19238 4612 19244
rect 4572 18826 4600 19238
rect 4744 19228 4796 19234
rect 4744 19170 4796 19176
rect 4560 18820 4612 18826
rect 4560 18762 4612 18768
rect 4756 18758 4784 19170
rect 5032 19030 5060 19782
rect 5204 19772 5256 19778
rect 5204 19714 5256 19720
rect 5020 19024 5072 19030
rect 5020 18966 5072 18972
rect 4744 18752 4796 18758
rect 4744 18694 4796 18700
rect 4468 18480 4520 18486
rect 4468 18422 4520 18428
rect 4192 18072 4244 18078
rect 4192 18014 4244 18020
rect 4480 17942 4508 18422
rect 4192 17936 4244 17942
rect 4192 17878 4244 17884
rect 4468 17936 4520 17942
rect 4468 17878 4520 17884
rect 4560 17936 4612 17942
rect 4560 17878 4612 17884
rect 4100 17188 4152 17194
rect 4100 17130 4152 17136
rect 4112 16650 4140 17130
rect 4204 16990 4232 17878
rect 4480 17602 4508 17878
rect 4468 17596 4520 17602
rect 4468 17538 4520 17544
rect 4376 17392 4428 17398
rect 4376 17334 4428 17340
rect 4192 16984 4244 16990
rect 4192 16926 4244 16932
rect 4100 16644 4152 16650
rect 4100 16586 4152 16592
rect 4284 16576 4336 16582
rect 4284 16518 4336 16524
rect 4296 16106 4324 16518
rect 4284 16100 4336 16106
rect 4284 16042 4336 16048
rect 3916 15556 3968 15562
rect 3916 15498 3968 15504
rect 4008 15556 4060 15562
rect 4008 15498 4060 15504
rect 2994 15391 3050 15400
rect 3272 15420 3324 15426
rect 3272 15362 3324 15368
rect 4388 14950 4416 17334
rect 4572 17194 4600 17878
rect 4756 17534 4784 18694
rect 4928 18480 4980 18486
rect 4928 18422 4980 18428
rect 4940 18282 4968 18422
rect 4928 18276 4980 18282
rect 4928 18218 4980 18224
rect 4928 18072 4980 18078
rect 4928 18014 4980 18020
rect 4940 17738 4968 18014
rect 5032 17942 5060 18966
rect 5020 17936 5072 17942
rect 5020 17878 5072 17884
rect 4928 17732 4980 17738
rect 4928 17674 4980 17680
rect 4940 17534 4968 17674
rect 4744 17528 4796 17534
rect 4744 17470 4796 17476
rect 4928 17528 4980 17534
rect 4928 17470 4980 17476
rect 4560 17188 4612 17194
rect 4560 17130 4612 17136
rect 4928 15896 4980 15902
rect 5032 15884 5060 17878
rect 4980 15856 5060 15884
rect 4928 15838 4980 15844
rect 4560 15012 4612 15018
rect 4560 14954 4612 14960
rect 4376 14944 4428 14950
rect 4376 14886 4428 14892
rect 3456 14876 3508 14882
rect 3376 14836 3456 14864
rect 3272 14808 3324 14814
rect 3272 14750 3324 14756
rect 3088 14672 3140 14678
rect 3088 14614 3140 14620
rect 3100 14474 3128 14614
rect 3088 14468 3140 14474
rect 3088 14410 3140 14416
rect 3284 14354 3312 14750
rect 3376 14474 3404 14836
rect 3456 14818 3508 14824
rect 4100 14740 4152 14746
rect 4100 14682 4152 14688
rect 3504 14572 3824 14592
rect 3504 14570 3516 14572
rect 3572 14570 3596 14572
rect 3652 14570 3676 14572
rect 3732 14570 3756 14572
rect 3812 14570 3824 14572
rect 3504 14518 3510 14570
rect 3572 14518 3574 14570
rect 3754 14518 3756 14570
rect 3818 14518 3824 14570
rect 3504 14516 3516 14518
rect 3572 14516 3596 14518
rect 3652 14516 3676 14518
rect 3732 14516 3756 14518
rect 3812 14516 3824 14518
rect 3504 14496 3824 14516
rect 3364 14468 3416 14474
rect 3364 14410 3416 14416
rect 3284 14326 3404 14354
rect 3088 14264 3140 14270
rect 3088 14206 3140 14212
rect 3270 14232 3326 14241
rect 2996 14128 3048 14134
rect 2996 14070 3048 14076
rect 3008 12094 3036 14070
rect 3100 13726 3128 14206
rect 3270 14167 3326 14176
rect 3284 14134 3312 14167
rect 3376 14134 3404 14326
rect 3272 14128 3324 14134
rect 3272 14070 3324 14076
rect 3364 14128 3416 14134
rect 3364 14070 3416 14076
rect 3088 13720 3140 13726
rect 3088 13662 3140 13668
rect 3284 13386 3312 14070
rect 3272 13380 3324 13386
rect 3272 13322 3324 13328
rect 3376 13250 3404 14070
rect 4008 13856 4060 13862
rect 4008 13798 4060 13804
rect 3504 13484 3824 13504
rect 3504 13482 3516 13484
rect 3572 13482 3596 13484
rect 3652 13482 3676 13484
rect 3732 13482 3756 13484
rect 3812 13482 3824 13484
rect 3504 13430 3510 13482
rect 3572 13430 3574 13482
rect 3754 13430 3756 13482
rect 3818 13430 3824 13482
rect 3504 13428 3516 13430
rect 3572 13428 3596 13430
rect 3652 13428 3676 13430
rect 3732 13428 3756 13430
rect 3812 13428 3824 13430
rect 3504 13408 3824 13428
rect 4020 13386 4048 13798
rect 4112 13794 4140 14682
rect 4192 14400 4244 14406
rect 4244 14360 4324 14388
rect 4192 14342 4244 14348
rect 4296 14241 4324 14360
rect 4388 14338 4416 14886
rect 4572 14474 4600 14954
rect 4940 14649 4968 15838
rect 5112 15352 5164 15358
rect 5112 15294 5164 15300
rect 5124 14950 5152 15294
rect 5112 14944 5164 14950
rect 5112 14886 5164 14892
rect 5020 14876 5072 14882
rect 5020 14818 5072 14824
rect 4926 14640 4982 14649
rect 4926 14575 4982 14584
rect 5032 14474 5060 14818
rect 4560 14468 4612 14474
rect 4560 14410 4612 14416
rect 5020 14468 5072 14474
rect 5020 14410 5072 14416
rect 5124 14338 5152 14886
rect 5216 14746 5244 19714
rect 5400 15018 5428 24950
rect 5492 24674 5520 24950
rect 6228 24810 6256 25086
rect 6216 24804 6268 24810
rect 6216 24746 6268 24752
rect 5480 24668 5532 24674
rect 5480 24610 5532 24616
rect 5492 24062 5520 24610
rect 5572 24600 5624 24606
rect 5572 24542 5624 24548
rect 5664 24600 5716 24606
rect 5664 24542 5716 24548
rect 5584 24198 5612 24542
rect 5676 24266 5704 24542
rect 5664 24260 5716 24266
rect 5664 24202 5716 24208
rect 5572 24192 5624 24198
rect 5572 24134 5624 24140
rect 5480 24056 5532 24062
rect 5480 23998 5532 24004
rect 5480 20316 5532 20322
rect 5480 20258 5532 20264
rect 5492 19914 5520 20258
rect 5584 20118 5612 24134
rect 5676 23178 5704 24202
rect 5756 23512 5808 23518
rect 5756 23454 5808 23460
rect 5664 23172 5716 23178
rect 5664 23114 5716 23120
rect 5768 22974 5796 23454
rect 5756 22968 5808 22974
rect 5756 22910 5808 22916
rect 5768 21886 5796 22910
rect 5756 21880 5808 21886
rect 5756 21822 5808 21828
rect 6032 21744 6084 21750
rect 6032 21686 6084 21692
rect 5756 20248 5808 20254
rect 5756 20190 5808 20196
rect 5940 20248 5992 20254
rect 5940 20190 5992 20196
rect 5572 20112 5624 20118
rect 5572 20054 5624 20060
rect 5480 19908 5532 19914
rect 5480 19850 5532 19856
rect 5768 19642 5796 20190
rect 5952 19710 5980 20190
rect 5940 19704 5992 19710
rect 5940 19646 5992 19652
rect 5756 19636 5808 19642
rect 5756 19578 5808 19584
rect 5952 19574 5980 19646
rect 5940 19568 5992 19574
rect 5940 19510 5992 19516
rect 5572 18548 5624 18554
rect 5572 18490 5624 18496
rect 5584 17738 5612 18490
rect 5572 17732 5624 17738
rect 5572 17674 5624 17680
rect 5584 17466 5612 17674
rect 5572 17460 5624 17466
rect 5572 17402 5624 17408
rect 5584 17176 5612 17402
rect 5584 17148 5704 17176
rect 5572 17052 5624 17058
rect 5572 16994 5624 17000
rect 5584 16650 5612 16994
rect 5676 16854 5704 17148
rect 5756 17120 5808 17126
rect 5756 17062 5808 17068
rect 5664 16848 5716 16854
rect 5664 16790 5716 16796
rect 5676 16650 5704 16790
rect 5572 16644 5624 16650
rect 5572 16586 5624 16592
rect 5664 16644 5716 16650
rect 5664 16586 5716 16592
rect 5480 16440 5532 16446
rect 5480 16382 5532 16388
rect 5492 16038 5520 16382
rect 5768 16310 5796 17062
rect 5952 16582 5980 19510
rect 5940 16576 5992 16582
rect 5940 16518 5992 16524
rect 5756 16304 5808 16310
rect 5756 16246 5808 16252
rect 5480 16032 5532 16038
rect 5480 15974 5532 15980
rect 5492 15222 5520 15974
rect 5572 15420 5624 15426
rect 5572 15362 5624 15368
rect 5480 15216 5532 15222
rect 5480 15158 5532 15164
rect 5388 15012 5440 15018
rect 5388 14954 5440 14960
rect 5296 14876 5348 14882
rect 5492 14864 5520 15158
rect 5348 14836 5520 14864
rect 5296 14818 5348 14824
rect 5204 14740 5256 14746
rect 5204 14682 5256 14688
rect 5202 14640 5258 14649
rect 5202 14575 5258 14584
rect 4376 14332 4428 14338
rect 4376 14274 4428 14280
rect 5112 14332 5164 14338
rect 5112 14274 5164 14280
rect 4282 14232 4338 14241
rect 4388 14214 4416 14274
rect 4388 14186 4508 14214
rect 4282 14167 4338 14176
rect 4296 13930 4324 14167
rect 4284 13924 4336 13930
rect 4284 13866 4336 13872
rect 4376 13924 4428 13930
rect 4376 13866 4428 13872
rect 4100 13788 4152 13794
rect 4100 13730 4152 13736
rect 4008 13380 4060 13386
rect 3928 13340 4008 13368
rect 3364 13244 3416 13250
rect 3364 13186 3416 13192
rect 3376 12162 3404 13186
rect 3504 12396 3824 12416
rect 3504 12394 3516 12396
rect 3572 12394 3596 12396
rect 3652 12394 3676 12396
rect 3732 12394 3756 12396
rect 3812 12394 3824 12396
rect 3504 12342 3510 12394
rect 3572 12342 3574 12394
rect 3754 12342 3756 12394
rect 3818 12342 3824 12394
rect 3504 12340 3516 12342
rect 3572 12340 3596 12342
rect 3652 12340 3676 12342
rect 3732 12340 3756 12342
rect 3812 12340 3824 12342
rect 3504 12320 3824 12340
rect 3364 12156 3416 12162
rect 3364 12098 3416 12104
rect 3732 12156 3784 12162
rect 3732 12098 3784 12104
rect 2996 12088 3048 12094
rect 2996 12030 3048 12036
rect 3744 11686 3772 12098
rect 3824 11952 3876 11958
rect 3824 11894 3876 11900
rect 3732 11680 3784 11686
rect 3732 11622 3784 11628
rect 3836 11618 3864 11894
rect 3928 11754 3956 13340
rect 4008 13322 4060 13328
rect 4008 13040 4060 13046
rect 4008 12982 4060 12988
rect 4020 12570 4048 12982
rect 4008 12564 4060 12570
rect 4008 12506 4060 12512
rect 4020 12026 4048 12506
rect 4112 12502 4140 13730
rect 4192 13652 4244 13658
rect 4192 13594 4244 13600
rect 4204 13250 4232 13594
rect 4192 13244 4244 13250
rect 4192 13186 4244 13192
rect 4388 13114 4416 13866
rect 4376 13108 4428 13114
rect 4376 13050 4428 13056
rect 4480 12502 4508 14186
rect 5124 13386 5152 14274
rect 5112 13380 5164 13386
rect 5112 13322 5164 13328
rect 5124 13182 5152 13322
rect 4652 13176 4704 13182
rect 4652 13118 4704 13124
rect 5112 13176 5164 13182
rect 5112 13118 5164 13124
rect 4560 13108 4612 13114
rect 4560 13050 4612 13056
rect 4100 12496 4152 12502
rect 4100 12438 4152 12444
rect 4468 12496 4520 12502
rect 4468 12438 4520 12444
rect 4008 12020 4060 12026
rect 4008 11962 4060 11968
rect 3916 11748 3968 11754
rect 3916 11690 3968 11696
rect 3824 11612 3876 11618
rect 3824 11554 3876 11560
rect 3504 11308 3824 11328
rect 3504 11306 3516 11308
rect 3572 11306 3596 11308
rect 3652 11306 3676 11308
rect 3732 11306 3756 11308
rect 3812 11306 3824 11308
rect 3504 11254 3510 11306
rect 3572 11254 3574 11306
rect 3754 11254 3756 11306
rect 3818 11254 3824 11306
rect 3504 11252 3516 11254
rect 3572 11252 3596 11254
rect 3652 11252 3676 11254
rect 3732 11252 3756 11254
rect 3812 11252 3824 11254
rect 3504 11232 3824 11252
rect 3364 11204 3416 11210
rect 3364 11146 3416 11152
rect 2904 11068 2956 11074
rect 2904 11010 2956 11016
rect 2628 11000 2680 11006
rect 2628 10942 2680 10948
rect 3272 11000 3324 11006
rect 3272 10942 3324 10948
rect 2640 10122 2668 10942
rect 2996 10864 3048 10870
rect 2996 10806 3048 10812
rect 3008 10666 3036 10806
rect 2996 10660 3048 10666
rect 2996 10602 3048 10608
rect 3008 10122 3036 10602
rect 3180 10524 3232 10530
rect 3180 10466 3232 10472
rect 3192 10122 3220 10466
rect 2628 10116 2680 10122
rect 2628 10058 2680 10064
rect 2996 10116 3048 10122
rect 2996 10058 3048 10064
rect 3180 10116 3232 10122
rect 3180 10058 3232 10064
rect 2640 9986 2668 10058
rect 3088 10048 3140 10054
rect 3088 9990 3140 9996
rect 2628 9980 2680 9986
rect 2628 9922 2680 9928
rect 2352 9436 2404 9442
rect 2456 9430 2668 9458
rect 2352 9378 2404 9384
rect 2364 8966 2392 9378
rect 2536 9368 2588 9374
rect 2536 9310 2588 9316
rect 2352 8960 2404 8966
rect 2352 8902 2404 8908
rect 2548 8694 2576 9310
rect 2536 8688 2588 8694
rect 2536 8630 2588 8636
rect 2352 6580 2404 6586
rect 2352 6522 2404 6528
rect 2364 6178 2392 6522
rect 2352 6172 2404 6178
rect 2352 6114 2404 6120
rect 2364 4682 2392 6114
rect 2444 4880 2496 4886
rect 2444 4822 2496 4828
rect 2352 4676 2404 4682
rect 2352 4618 2404 4624
rect 2456 4478 2484 4822
rect 2444 4472 2496 4478
rect 2444 4414 2496 4420
rect 2456 3866 2484 4414
rect 2444 3860 2496 3866
rect 2444 3802 2496 3808
rect 2548 1826 2576 8630
rect 2640 4554 2668 9430
rect 2996 9368 3048 9374
rect 2996 9310 3048 9316
rect 3008 9034 3036 9310
rect 3100 9238 3128 9990
rect 3284 9578 3312 10942
rect 3376 10938 3404 11146
rect 3928 11142 3956 11690
rect 4020 11210 4048 11962
rect 4008 11204 4060 11210
rect 4008 11146 4060 11152
rect 3916 11136 3968 11142
rect 3916 11078 3968 11084
rect 4112 10988 4140 12438
rect 4468 12224 4520 12230
rect 4468 12166 4520 12172
rect 4284 12088 4336 12094
rect 4284 12030 4336 12036
rect 3928 10960 4140 10988
rect 4192 11000 4244 11006
rect 3364 10932 3416 10938
rect 3364 10874 3416 10880
rect 3272 9572 3324 9578
rect 3272 9514 3324 9520
rect 3180 9504 3232 9510
rect 3180 9446 3232 9452
rect 3088 9232 3140 9238
rect 3088 9174 3140 9180
rect 2996 9028 3048 9034
rect 2996 8970 3048 8976
rect 3100 8966 3128 9174
rect 3192 9034 3220 9446
rect 3376 9442 3404 10874
rect 3928 10530 3956 10960
rect 4192 10942 4244 10948
rect 3916 10524 3968 10530
rect 3916 10466 3968 10472
rect 3928 10326 3956 10466
rect 3916 10320 3968 10326
rect 3916 10262 3968 10268
rect 3504 10220 3824 10240
rect 3504 10218 3516 10220
rect 3572 10218 3596 10220
rect 3652 10218 3676 10220
rect 3732 10218 3756 10220
rect 3812 10218 3824 10220
rect 3504 10166 3510 10218
rect 3572 10166 3574 10218
rect 3754 10166 3756 10218
rect 3818 10166 3824 10218
rect 3504 10164 3516 10166
rect 3572 10164 3596 10166
rect 3652 10164 3676 10166
rect 3732 10164 3756 10166
rect 3812 10164 3824 10166
rect 3504 10144 3824 10164
rect 4204 10122 4232 10942
rect 4296 10666 4324 12030
rect 4480 11958 4508 12166
rect 4572 12026 4600 13050
rect 4664 12230 4692 13118
rect 4928 12768 4980 12774
rect 4928 12710 4980 12716
rect 4836 12700 4888 12706
rect 4836 12642 4888 12648
rect 4744 12632 4796 12638
rect 4744 12574 4796 12580
rect 4756 12230 4784 12574
rect 4652 12224 4704 12230
rect 4652 12166 4704 12172
rect 4744 12224 4796 12230
rect 4744 12166 4796 12172
rect 4848 12076 4876 12642
rect 4664 12048 4876 12076
rect 4560 12020 4612 12026
rect 4560 11962 4612 11968
rect 4468 11952 4520 11958
rect 4468 11894 4520 11900
rect 4480 11754 4508 11894
rect 4468 11748 4520 11754
rect 4468 11690 4520 11696
rect 4376 11408 4428 11414
rect 4376 11350 4428 11356
rect 4388 11210 4416 11350
rect 4480 11210 4508 11690
rect 4572 11618 4600 11962
rect 4664 11958 4692 12048
rect 4940 11958 4968 12710
rect 5216 12638 5244 14575
rect 5400 14134 5428 14836
rect 5388 14128 5440 14134
rect 5388 14070 5440 14076
rect 5296 13108 5348 13114
rect 5296 13050 5348 13056
rect 5204 12632 5256 12638
rect 5204 12574 5256 12580
rect 5216 12298 5244 12574
rect 5204 12292 5256 12298
rect 5204 12234 5256 12240
rect 4652 11952 4704 11958
rect 4652 11894 4704 11900
rect 4928 11952 4980 11958
rect 4928 11894 4980 11900
rect 4560 11612 4612 11618
rect 4560 11554 4612 11560
rect 4376 11204 4428 11210
rect 4376 11146 4428 11152
rect 4468 11204 4520 11210
rect 4468 11146 4520 11152
rect 4284 10660 4336 10666
rect 4388 10648 4416 11146
rect 4664 11142 4692 11894
rect 4940 11550 4968 11894
rect 4744 11544 4796 11550
rect 4744 11486 4796 11492
rect 4928 11544 4980 11550
rect 4928 11486 4980 11492
rect 4652 11136 4704 11142
rect 4652 11078 4704 11084
rect 4756 11006 4784 11486
rect 4652 11000 4704 11006
rect 4652 10942 4704 10948
rect 4744 11000 4796 11006
rect 4744 10942 4796 10948
rect 4468 10660 4520 10666
rect 4388 10620 4468 10648
rect 4284 10602 4336 10608
rect 4468 10602 4520 10608
rect 4296 10530 4324 10602
rect 4664 10546 4692 10942
rect 4284 10524 4336 10530
rect 4468 10524 4520 10530
rect 4284 10466 4336 10472
rect 4388 10484 4468 10512
rect 4192 10116 4244 10122
rect 4192 10058 4244 10064
rect 4100 9844 4152 9850
rect 4100 9786 4152 9792
rect 3364 9436 3416 9442
rect 3364 9378 3416 9384
rect 3180 9028 3232 9034
rect 3180 8970 3232 8976
rect 3088 8960 3140 8966
rect 3088 8902 3140 8908
rect 3376 8490 3404 9378
rect 3916 9300 3968 9306
rect 3916 9242 3968 9248
rect 3504 9132 3824 9152
rect 3504 9130 3516 9132
rect 3572 9130 3596 9132
rect 3652 9130 3676 9132
rect 3732 9130 3756 9132
rect 3812 9130 3824 9132
rect 3504 9078 3510 9130
rect 3572 9078 3574 9130
rect 3754 9078 3756 9130
rect 3818 9078 3824 9130
rect 3504 9076 3516 9078
rect 3572 9076 3596 9078
rect 3652 9076 3676 9078
rect 3732 9076 3756 9078
rect 3812 9076 3824 9078
rect 3504 9056 3824 9076
rect 3928 9034 3956 9242
rect 3916 9028 3968 9034
rect 3916 8970 3968 8976
rect 3364 8484 3416 8490
rect 3364 8426 3416 8432
rect 4008 8348 4060 8354
rect 4112 8336 4140 9786
rect 4388 9782 4416 10484
rect 4468 10466 4520 10472
rect 4572 10518 4692 10546
rect 4572 9918 4600 10518
rect 4756 10462 4784 10942
rect 4940 10598 4968 11486
rect 5204 11476 5256 11482
rect 5308 11464 5336 13050
rect 5400 13046 5428 14070
rect 5388 13040 5440 13046
rect 5388 12982 5440 12988
rect 5584 11482 5612 15362
rect 5768 14814 5796 16246
rect 5940 15964 5992 15970
rect 5940 15906 5992 15912
rect 5848 15896 5900 15902
rect 5848 15838 5900 15844
rect 5860 15426 5888 15838
rect 5848 15420 5900 15426
rect 5848 15362 5900 15368
rect 5952 15018 5980 15906
rect 5940 15012 5992 15018
rect 5940 14954 5992 14960
rect 5848 14944 5900 14950
rect 5848 14886 5900 14892
rect 5756 14808 5808 14814
rect 5756 14750 5808 14756
rect 5768 14270 5796 14750
rect 5860 14678 5888 14886
rect 5848 14672 5900 14678
rect 5848 14614 5900 14620
rect 5756 14264 5808 14270
rect 5756 14206 5808 14212
rect 5756 14128 5808 14134
rect 5860 14116 5888 14614
rect 5808 14088 5888 14116
rect 5756 14070 5808 14076
rect 5664 13856 5716 13862
rect 5664 13798 5716 13804
rect 5676 13182 5704 13798
rect 5768 13182 5796 14070
rect 5848 13720 5900 13726
rect 5848 13662 5900 13668
rect 5664 13176 5716 13182
rect 5664 13118 5716 13124
rect 5756 13176 5808 13182
rect 5756 13118 5808 13124
rect 5676 13017 5704 13118
rect 5756 13040 5808 13046
rect 5662 13008 5718 13017
rect 5756 12982 5808 12988
rect 5662 12943 5718 12952
rect 5664 12156 5716 12162
rect 5664 12098 5716 12104
rect 5256 11436 5336 11464
rect 5572 11476 5624 11482
rect 5204 11418 5256 11424
rect 5572 11418 5624 11424
rect 5216 10870 5244 11418
rect 5584 11142 5612 11418
rect 5572 11136 5624 11142
rect 5572 11078 5624 11084
rect 5204 10864 5256 10870
rect 5204 10806 5256 10812
rect 4928 10592 4980 10598
rect 4928 10534 4980 10540
rect 4744 10456 4796 10462
rect 4744 10398 4796 10404
rect 4652 10388 4704 10394
rect 4652 10330 4704 10336
rect 4664 10122 4692 10330
rect 4652 10116 4704 10122
rect 4652 10058 4704 10064
rect 4756 10002 4784 10398
rect 4664 9974 4784 10002
rect 4560 9912 4612 9918
rect 4560 9854 4612 9860
rect 4376 9776 4428 9782
rect 4296 9736 4376 9764
rect 4192 9436 4244 9442
rect 4192 9378 4244 9384
rect 4204 8898 4232 9378
rect 4296 9238 4324 9736
rect 4376 9718 4428 9724
rect 4560 9436 4612 9442
rect 4560 9378 4612 9384
rect 4376 9300 4428 9306
rect 4376 9242 4428 9248
rect 4284 9232 4336 9238
rect 4284 9174 4336 9180
rect 4296 9034 4324 9174
rect 4284 9028 4336 9034
rect 4284 8970 4336 8976
rect 4192 8892 4244 8898
rect 4192 8834 4244 8840
rect 4204 8762 4232 8834
rect 4388 8830 4416 9242
rect 4572 8966 4600 9378
rect 4560 8960 4612 8966
rect 4560 8902 4612 8908
rect 4376 8824 4428 8830
rect 4376 8766 4428 8772
rect 4192 8756 4244 8762
rect 4192 8698 4244 8704
rect 4204 8354 4232 8698
rect 4664 8490 4692 9974
rect 5216 9510 5244 10806
rect 5676 10598 5704 12098
rect 5768 11618 5796 12982
rect 5756 11612 5808 11618
rect 5756 11554 5808 11560
rect 5664 10592 5716 10598
rect 5664 10534 5716 10540
rect 5296 10524 5348 10530
rect 5296 10466 5348 10472
rect 5308 10122 5336 10466
rect 5676 10122 5704 10534
rect 5296 10116 5348 10122
rect 5296 10058 5348 10064
rect 5664 10116 5716 10122
rect 5664 10058 5716 10064
rect 5204 9504 5256 9510
rect 5204 9446 5256 9452
rect 5112 9368 5164 9374
rect 5216 9356 5244 9446
rect 5164 9328 5244 9356
rect 5112 9310 5164 9316
rect 4928 9232 4980 9238
rect 4928 9174 4980 9180
rect 4940 9034 4968 9174
rect 4928 9028 4980 9034
rect 4928 8970 4980 8976
rect 4744 8688 4796 8694
rect 4744 8630 4796 8636
rect 4652 8484 4704 8490
rect 4652 8426 4704 8432
rect 4376 8416 4428 8422
rect 4376 8358 4428 8364
rect 4060 8308 4140 8336
rect 4008 8290 4060 8296
rect 3504 8044 3824 8064
rect 3504 8042 3516 8044
rect 3572 8042 3596 8044
rect 3652 8042 3676 8044
rect 3732 8042 3756 8044
rect 3812 8042 3824 8044
rect 3504 7990 3510 8042
rect 3572 7990 3574 8042
rect 3754 7990 3756 8042
rect 3818 7990 3824 8042
rect 3504 7988 3516 7990
rect 3572 7988 3596 7990
rect 3652 7988 3676 7990
rect 3732 7988 3756 7990
rect 3812 7988 3824 7990
rect 3504 7968 3824 7988
rect 3364 7192 3416 7198
rect 3364 7134 3416 7140
rect 2996 6580 3048 6586
rect 2996 6522 3048 6528
rect 3008 5634 3036 6522
rect 3376 6314 3404 7134
rect 3504 6956 3824 6976
rect 3504 6954 3516 6956
rect 3572 6954 3596 6956
rect 3652 6954 3676 6956
rect 3732 6954 3756 6956
rect 3812 6954 3824 6956
rect 3504 6902 3510 6954
rect 3572 6902 3574 6954
rect 3754 6902 3756 6954
rect 3818 6902 3824 6954
rect 3504 6900 3516 6902
rect 3572 6900 3596 6902
rect 3652 6900 3676 6902
rect 3732 6900 3756 6902
rect 3812 6900 3824 6902
rect 3504 6880 3824 6900
rect 3364 6308 3416 6314
rect 3364 6250 3416 6256
rect 3272 6172 3324 6178
rect 3272 6114 3324 6120
rect 3284 5770 3312 6114
rect 3272 5764 3324 5770
rect 3272 5706 3324 5712
rect 2996 5628 3048 5634
rect 2996 5570 3048 5576
rect 3272 5492 3324 5498
rect 3272 5434 3324 5440
rect 2640 4526 2760 4554
rect 2732 4070 2760 4526
rect 3284 4070 3312 5434
rect 3376 5226 3404 6250
rect 4112 5956 4140 8308
rect 4192 8348 4244 8354
rect 4192 8290 4244 8296
rect 4204 7946 4232 8290
rect 4388 7946 4416 8358
rect 4756 8354 4784 8630
rect 5308 8490 5336 10058
rect 5296 8484 5348 8490
rect 5296 8426 5348 8432
rect 4744 8348 4796 8354
rect 4744 8290 4796 8296
rect 5756 8348 5808 8354
rect 5756 8290 5808 8296
rect 5768 7946 5796 8290
rect 4192 7940 4244 7946
rect 4192 7882 4244 7888
rect 4376 7940 4428 7946
rect 4376 7882 4428 7888
rect 5756 7940 5808 7946
rect 5756 7882 5808 7888
rect 5860 7266 5888 13662
rect 5940 12020 5992 12026
rect 5940 11962 5992 11968
rect 5952 11686 5980 11962
rect 5940 11680 5992 11686
rect 5940 11622 5992 11628
rect 5952 11210 5980 11622
rect 5940 11204 5992 11210
rect 5940 11146 5992 11152
rect 5848 7260 5900 7266
rect 5848 7202 5900 7208
rect 5860 6858 5888 7202
rect 5848 6852 5900 6858
rect 5848 6794 5900 6800
rect 6044 6654 6072 21686
rect 6216 20656 6268 20662
rect 6216 20598 6268 20604
rect 6228 20118 6256 20598
rect 6216 20112 6268 20118
rect 6216 20054 6268 20060
rect 6228 19914 6256 20054
rect 6216 19908 6268 19914
rect 6216 19850 6268 19856
rect 6228 19302 6256 19850
rect 6216 19296 6268 19302
rect 6216 19238 6268 19244
rect 6320 18690 6348 27315
rect 6492 26776 6544 26782
rect 6492 26718 6544 26724
rect 6400 26232 6452 26238
rect 6400 26174 6452 26180
rect 6412 25762 6440 26174
rect 6504 26102 6532 26718
rect 6676 26708 6728 26714
rect 6676 26650 6728 26656
rect 6688 26442 6716 26650
rect 7688 26640 7740 26646
rect 7688 26582 7740 26588
rect 6676 26436 6728 26442
rect 6676 26378 6728 26384
rect 6492 26096 6544 26102
rect 6492 26038 6544 26044
rect 6400 25756 6452 25762
rect 6400 25698 6452 25704
rect 6412 24674 6440 25698
rect 6504 25558 6532 26038
rect 6492 25552 6544 25558
rect 6492 25494 6544 25500
rect 6688 25150 6716 26378
rect 7700 26238 7728 26582
rect 7320 26232 7372 26238
rect 7320 26174 7372 26180
rect 7688 26232 7740 26238
rect 7688 26174 7740 26180
rect 7332 26102 7360 26174
rect 7412 26164 7464 26170
rect 7412 26106 7464 26112
rect 7320 26096 7372 26102
rect 7320 26038 7372 26044
rect 7424 25898 7452 26106
rect 7412 25892 7464 25898
rect 7412 25834 7464 25840
rect 6768 25756 6820 25762
rect 6768 25698 6820 25704
rect 6780 25354 6808 25698
rect 6768 25348 6820 25354
rect 6768 25290 6820 25296
rect 6676 25144 6728 25150
rect 6676 25086 6728 25092
rect 7412 25144 7464 25150
rect 7412 25086 7464 25092
rect 6952 25008 7004 25014
rect 6952 24950 7004 24956
rect 6964 24810 6992 24950
rect 7424 24810 7452 25086
rect 6952 24804 7004 24810
rect 6952 24746 7004 24752
rect 7412 24804 7464 24810
rect 7412 24746 7464 24752
rect 6490 24704 6546 24713
rect 6400 24668 6452 24674
rect 6490 24639 6546 24648
rect 6400 24610 6452 24616
rect 6412 22090 6440 24610
rect 6504 24606 6532 24639
rect 6492 24600 6544 24606
rect 6492 24542 6544 24548
rect 6504 24130 6532 24542
rect 6964 24266 6992 24746
rect 6952 24260 7004 24266
rect 6952 24202 7004 24208
rect 7424 24198 7452 24746
rect 7504 24464 7556 24470
rect 7504 24406 7556 24412
rect 7516 24266 7544 24406
rect 7504 24260 7556 24266
rect 7504 24202 7556 24208
rect 7412 24192 7464 24198
rect 7412 24134 7464 24140
rect 6492 24124 6544 24130
rect 6492 24066 6544 24072
rect 7412 24056 7464 24062
rect 7412 23998 7464 24004
rect 7424 23518 7452 23998
rect 7516 23654 7544 24202
rect 7504 23648 7556 23654
rect 7504 23590 7556 23596
rect 7412 23512 7464 23518
rect 7412 23454 7464 23460
rect 7424 23042 7452 23454
rect 7516 23178 7544 23590
rect 7504 23172 7556 23178
rect 7504 23114 7556 23120
rect 7412 23036 7464 23042
rect 7412 22978 7464 22984
rect 6400 22084 6452 22090
rect 6400 22026 6452 22032
rect 7424 21954 7452 22978
rect 7412 21948 7464 21954
rect 7412 21890 7464 21896
rect 7424 21546 7452 21890
rect 7412 21540 7464 21546
rect 7412 21482 7464 21488
rect 7700 21410 7728 26174
rect 8344 25830 8372 27315
rect 10092 27311 10396 27315
rect 9068 26096 9120 26102
rect 9068 26038 9120 26044
rect 8332 25824 8384 25830
rect 8332 25766 8384 25772
rect 7780 25552 7832 25558
rect 7780 25494 7832 25500
rect 8424 25552 8476 25558
rect 8424 25494 8476 25500
rect 7792 25354 7820 25494
rect 7780 25348 7832 25354
rect 7780 25290 7832 25296
rect 8436 25014 8464 25494
rect 9080 25218 9108 26038
rect 9252 25824 9304 25830
rect 9252 25766 9304 25772
rect 9160 25688 9212 25694
rect 9160 25630 9212 25636
rect 9068 25212 9120 25218
rect 9068 25154 9120 25160
rect 9172 25082 9200 25630
rect 9264 25150 9292 25766
rect 10092 25762 10120 27311
rect 12208 26306 12236 27315
rect 12196 26300 12248 26306
rect 12196 26242 12248 26248
rect 11736 26232 11788 26238
rect 11736 26174 11788 26180
rect 11748 25830 11776 26174
rect 12196 26164 12248 26170
rect 12196 26106 12248 26112
rect 12472 26164 12524 26170
rect 12472 26106 12524 26112
rect 11736 25824 11788 25830
rect 11736 25766 11788 25772
rect 10080 25756 10132 25762
rect 10080 25698 10132 25704
rect 10264 25756 10316 25762
rect 10264 25698 10316 25704
rect 10092 25354 10120 25698
rect 10080 25348 10132 25354
rect 10080 25290 10132 25296
rect 10276 25218 10304 25698
rect 11092 25688 11144 25694
rect 11092 25630 11144 25636
rect 10448 25280 10500 25286
rect 10448 25222 10500 25228
rect 10264 25212 10316 25218
rect 10264 25154 10316 25160
rect 9252 25144 9304 25150
rect 9252 25086 9304 25092
rect 9804 25144 9856 25150
rect 9804 25086 9856 25092
rect 9160 25076 9212 25082
rect 9160 25018 9212 25024
rect 8424 25008 8476 25014
rect 8424 24950 8476 24956
rect 7964 24464 8016 24470
rect 7964 24406 8016 24412
rect 7976 23450 8004 24406
rect 8436 24062 8464 24950
rect 8424 24056 8476 24062
rect 8424 23998 8476 24004
rect 9068 23988 9120 23994
rect 9068 23930 9120 23936
rect 7964 23444 8016 23450
rect 7964 23386 8016 23392
rect 7976 22974 8004 23386
rect 9080 22974 9108 23930
rect 7964 22968 8016 22974
rect 7964 22910 8016 22916
rect 9068 22968 9120 22974
rect 9068 22910 9120 22916
rect 8884 22900 8936 22906
rect 8884 22842 8936 22848
rect 7780 22288 7832 22294
rect 7780 22230 7832 22236
rect 7792 21886 7820 22230
rect 8332 22084 8384 22090
rect 8332 22026 8384 22032
rect 8344 21886 8372 22026
rect 8700 21948 8752 21954
rect 8700 21890 8752 21896
rect 7780 21880 7832 21886
rect 7780 21822 7832 21828
rect 8332 21880 8384 21886
rect 8332 21822 8384 21828
rect 7688 21404 7740 21410
rect 7688 21346 7740 21352
rect 7044 20724 7096 20730
rect 7044 20666 7096 20672
rect 6400 20452 6452 20458
rect 6400 20394 6452 20400
rect 6412 19914 6440 20394
rect 7056 20322 7084 20666
rect 7044 20316 7096 20322
rect 7044 20258 7096 20264
rect 6860 20112 6912 20118
rect 6860 20054 6912 20060
rect 6400 19908 6452 19914
rect 6400 19850 6452 19856
rect 6872 19710 6900 20054
rect 7056 19914 7084 20258
rect 7700 20254 7728 21346
rect 7792 20458 7820 21822
rect 7780 20452 7832 20458
rect 7780 20394 7832 20400
rect 8148 20452 8200 20458
rect 8148 20394 8200 20400
rect 7688 20248 7740 20254
rect 7688 20190 7740 20196
rect 7320 20180 7372 20186
rect 7320 20122 7372 20128
rect 7332 19914 7360 20122
rect 7044 19908 7096 19914
rect 7044 19850 7096 19856
rect 7320 19908 7372 19914
rect 7320 19850 7372 19856
rect 6860 19704 6912 19710
rect 6860 19646 6912 19652
rect 6584 19636 6636 19642
rect 6584 19578 6636 19584
rect 6308 18684 6360 18690
rect 6308 18626 6360 18632
rect 6308 18480 6360 18486
rect 6308 18422 6360 18428
rect 6320 18146 6348 18422
rect 6596 18282 6624 19578
rect 7056 19302 7084 19850
rect 7136 19568 7188 19574
rect 7136 19510 7188 19516
rect 7044 19296 7096 19302
rect 7044 19238 7096 19244
rect 7056 18826 7084 19238
rect 7044 18820 7096 18826
rect 7044 18762 7096 18768
rect 7044 18684 7096 18690
rect 7044 18626 7096 18632
rect 6584 18276 6636 18282
rect 6584 18218 6636 18224
rect 6308 18140 6360 18146
rect 6308 18082 6360 18088
rect 6216 18072 6268 18078
rect 6216 18014 6268 18020
rect 6124 17460 6176 17466
rect 6124 17402 6176 17408
rect 6136 17058 6164 17402
rect 6124 17052 6176 17058
rect 6124 16994 6176 17000
rect 6228 16922 6256 18014
rect 6320 16922 6348 18082
rect 6596 17738 6624 18218
rect 6860 18072 6912 18078
rect 6860 18014 6912 18020
rect 6872 17738 6900 18014
rect 6584 17732 6636 17738
rect 6584 17674 6636 17680
rect 6860 17732 6912 17738
rect 6860 17674 6912 17680
rect 6400 17664 6452 17670
rect 6400 17606 6452 17612
rect 6412 17534 6440 17606
rect 6400 17528 6452 17534
rect 6400 17470 6452 17476
rect 6860 17460 6912 17466
rect 6860 17402 6912 17408
rect 6216 16916 6268 16922
rect 6216 16858 6268 16864
rect 6308 16916 6360 16922
rect 6308 16858 6360 16864
rect 6216 16032 6268 16038
rect 6216 15974 6268 15980
rect 6584 16032 6636 16038
rect 6584 15974 6636 15980
rect 6228 15018 6256 15974
rect 6308 15760 6360 15766
rect 6308 15702 6360 15708
rect 6320 15222 6348 15702
rect 6308 15216 6360 15222
rect 6308 15158 6360 15164
rect 6400 15216 6452 15222
rect 6400 15158 6452 15164
rect 6216 15012 6268 15018
rect 6216 14954 6268 14960
rect 6124 14876 6176 14882
rect 6124 14818 6176 14824
rect 6136 14134 6164 14818
rect 6124 14128 6176 14134
rect 6124 14070 6176 14076
rect 6216 14128 6268 14134
rect 6216 14070 6268 14076
rect 6136 13590 6164 14070
rect 6124 13584 6176 13590
rect 6124 13526 6176 13532
rect 6136 13114 6164 13526
rect 6124 13108 6176 13114
rect 6124 13050 6176 13056
rect 6228 11958 6256 14070
rect 6320 13930 6348 15158
rect 6412 14678 6440 15158
rect 6596 14950 6624 15974
rect 6676 15896 6728 15902
rect 6676 15838 6728 15844
rect 6688 15426 6716 15838
rect 6872 15426 6900 17402
rect 6952 17052 7004 17058
rect 6952 16994 7004 17000
rect 6964 16650 6992 16994
rect 6952 16644 7004 16650
rect 6952 16586 7004 16592
rect 6964 15494 6992 16586
rect 6952 15488 7004 15494
rect 6952 15430 7004 15436
rect 6676 15420 6728 15426
rect 6676 15362 6728 15368
rect 6860 15420 6912 15426
rect 6860 15362 6912 15368
rect 6676 15012 6728 15018
rect 6676 14954 6728 14960
rect 6584 14944 6636 14950
rect 6584 14886 6636 14892
rect 6492 14740 6544 14746
rect 6492 14682 6544 14688
rect 6400 14672 6452 14678
rect 6400 14614 6452 14620
rect 6504 14474 6532 14682
rect 6492 14468 6544 14474
rect 6492 14410 6544 14416
rect 6584 14400 6636 14406
rect 6584 14342 6636 14348
rect 6308 13924 6360 13930
rect 6308 13866 6360 13872
rect 6308 13312 6360 13318
rect 6308 13254 6360 13260
rect 6320 13046 6348 13254
rect 6308 13040 6360 13046
rect 6308 12982 6360 12988
rect 6492 12768 6544 12774
rect 6492 12710 6544 12716
rect 6400 12632 6452 12638
rect 6400 12574 6452 12580
rect 6308 12496 6360 12502
rect 6308 12438 6360 12444
rect 6320 12094 6348 12438
rect 6412 12298 6440 12574
rect 6504 12502 6532 12710
rect 6492 12496 6544 12502
rect 6492 12438 6544 12444
rect 6596 12298 6624 14342
rect 6688 14105 6716 14954
rect 6872 14882 6900 15362
rect 6860 14876 6912 14882
rect 6860 14818 6912 14824
rect 6952 14808 7004 14814
rect 6952 14750 7004 14756
rect 6768 14740 6820 14746
rect 6768 14682 6820 14688
rect 6674 14096 6730 14105
rect 6674 14031 6730 14040
rect 6688 13386 6716 14031
rect 6676 13380 6728 13386
rect 6676 13322 6728 13328
rect 6688 13046 6716 13322
rect 6676 13040 6728 13046
rect 6676 12982 6728 12988
rect 6400 12292 6452 12298
rect 6400 12234 6452 12240
rect 6584 12292 6636 12298
rect 6584 12234 6636 12240
rect 6308 12088 6360 12094
rect 6308 12030 6360 12036
rect 6216 11952 6268 11958
rect 6216 11894 6268 11900
rect 6400 11612 6452 11618
rect 6400 11554 6452 11560
rect 6308 11408 6360 11414
rect 6308 11350 6360 11356
rect 6124 9912 6176 9918
rect 6124 9854 6176 9860
rect 6136 8150 6164 9854
rect 6216 8892 6268 8898
rect 6216 8834 6268 8840
rect 6228 8762 6256 8834
rect 6216 8756 6268 8762
rect 6216 8698 6268 8704
rect 6320 8694 6348 11350
rect 6412 11142 6440 11554
rect 6688 11550 6716 12982
rect 6780 11668 6808 14682
rect 6860 14672 6912 14678
rect 6860 14614 6912 14620
rect 6872 14474 6900 14614
rect 6964 14474 6992 14750
rect 6860 14468 6912 14474
rect 6860 14410 6912 14416
rect 6952 14468 7004 14474
rect 6952 14410 7004 14416
rect 6860 13788 6912 13794
rect 6860 13730 6912 13736
rect 6872 13386 6900 13730
rect 6860 13380 6912 13386
rect 6860 13322 6912 13328
rect 6860 13108 6912 13114
rect 6860 13050 6912 13056
rect 6872 13017 6900 13050
rect 6858 13008 6914 13017
rect 6858 12943 6914 12952
rect 6860 11680 6912 11686
rect 6780 11640 6860 11668
rect 6860 11622 6912 11628
rect 6676 11544 6728 11550
rect 6676 11486 6728 11492
rect 6688 11210 6716 11486
rect 6768 11476 6820 11482
rect 6768 11418 6820 11424
rect 6676 11204 6728 11210
rect 6676 11146 6728 11152
rect 6400 11136 6452 11142
rect 6400 11078 6452 11084
rect 6492 9844 6544 9850
rect 6492 9786 6544 9792
rect 6400 9504 6452 9510
rect 6400 9446 6452 9452
rect 6308 8688 6360 8694
rect 6308 8630 6360 8636
rect 6412 8422 6440 9446
rect 6504 8762 6532 9786
rect 6688 9442 6716 11146
rect 6780 10122 6808 11418
rect 6768 10116 6820 10122
rect 6768 10058 6820 10064
rect 6676 9436 6728 9442
rect 6676 9378 6728 9384
rect 6952 9436 7004 9442
rect 6952 9378 7004 9384
rect 6688 9306 6716 9378
rect 6768 9368 6820 9374
rect 6768 9310 6820 9316
rect 6676 9300 6728 9306
rect 6676 9242 6728 9248
rect 6584 9232 6636 9238
rect 6584 9174 6636 9180
rect 6492 8756 6544 8762
rect 6492 8698 6544 8704
rect 6400 8416 6452 8422
rect 6400 8358 6452 8364
rect 6124 8144 6176 8150
rect 6124 8086 6176 8092
rect 6136 7946 6164 8086
rect 6124 7940 6176 7946
rect 6124 7882 6176 7888
rect 6596 7334 6624 9174
rect 6688 8694 6716 9242
rect 6780 8966 6808 9310
rect 6964 9034 6992 9378
rect 6952 9028 7004 9034
rect 6952 8970 7004 8976
rect 6768 8960 6820 8966
rect 6768 8902 6820 8908
rect 6860 8756 6912 8762
rect 6860 8698 6912 8704
rect 6676 8688 6728 8694
rect 6676 8630 6728 8636
rect 6688 8422 6716 8630
rect 6872 8490 6900 8698
rect 6860 8484 6912 8490
rect 6860 8426 6912 8432
rect 6676 8416 6728 8422
rect 6676 8358 6728 8364
rect 6584 7328 6636 7334
rect 6504 7288 6584 7316
rect 6504 6790 6532 7288
rect 6584 7270 6636 7276
rect 6676 7260 6728 7266
rect 6676 7202 6728 7208
rect 6584 7124 6636 7130
rect 6584 7066 6636 7072
rect 6492 6784 6544 6790
rect 6492 6726 6544 6732
rect 6032 6648 6084 6654
rect 6032 6590 6084 6596
rect 5664 6172 5716 6178
rect 5664 6114 5716 6120
rect 4836 6104 4888 6110
rect 4836 6046 4888 6052
rect 5388 6104 5440 6110
rect 5388 6046 5440 6052
rect 4192 5968 4244 5974
rect 4112 5928 4192 5956
rect 4192 5910 4244 5916
rect 3504 5868 3824 5888
rect 3504 5866 3516 5868
rect 3572 5866 3596 5868
rect 3652 5866 3676 5868
rect 3732 5866 3756 5868
rect 3812 5866 3824 5868
rect 3504 5814 3510 5866
rect 3572 5814 3574 5866
rect 3754 5814 3756 5866
rect 3818 5814 3824 5866
rect 3504 5812 3516 5814
rect 3572 5812 3596 5814
rect 3652 5812 3676 5814
rect 3732 5812 3756 5814
rect 3812 5812 3824 5814
rect 3504 5792 3824 5812
rect 4204 5566 4232 5910
rect 4848 5770 4876 6046
rect 5400 5770 5428 6046
rect 5676 5770 5704 6114
rect 6044 5770 6072 6590
rect 6596 6586 6624 7066
rect 6688 6858 6716 7202
rect 6676 6852 6728 6858
rect 6676 6794 6728 6800
rect 6584 6580 6636 6586
rect 6584 6522 6636 6528
rect 6596 6246 6624 6522
rect 6584 6240 6636 6246
rect 6584 6182 6636 6188
rect 6400 6172 6452 6178
rect 6400 6114 6452 6120
rect 6412 5770 6440 6114
rect 4836 5764 4888 5770
rect 4836 5706 4888 5712
rect 5388 5764 5440 5770
rect 5388 5706 5440 5712
rect 5664 5764 5716 5770
rect 5664 5706 5716 5712
rect 6032 5764 6084 5770
rect 6032 5706 6084 5712
rect 6400 5764 6452 5770
rect 6400 5706 6452 5712
rect 4744 5696 4796 5702
rect 4744 5638 4796 5644
rect 4468 5628 4520 5634
rect 4468 5570 4520 5576
rect 4192 5560 4244 5566
rect 4192 5502 4244 5508
rect 4008 5492 4060 5498
rect 4008 5434 4060 5440
rect 3364 5220 3416 5226
rect 3364 5162 3416 5168
rect 3504 4780 3824 4800
rect 3504 4778 3516 4780
rect 3572 4778 3596 4780
rect 3652 4778 3676 4780
rect 3732 4778 3756 4780
rect 3812 4778 3824 4780
rect 3504 4726 3510 4778
rect 3572 4726 3574 4778
rect 3754 4726 3756 4778
rect 3818 4726 3824 4778
rect 3504 4724 3516 4726
rect 3572 4724 3596 4726
rect 3652 4724 3676 4726
rect 3732 4724 3756 4726
rect 3812 4724 3824 4726
rect 3504 4704 3824 4724
rect 4020 4410 4048 5434
rect 4480 5430 4508 5570
rect 4756 5566 4784 5638
rect 4744 5560 4796 5566
rect 4744 5502 4796 5508
rect 4468 5424 4520 5430
rect 4468 5366 4520 5372
rect 4480 5226 4508 5366
rect 4468 5220 4520 5226
rect 4468 5162 4520 5168
rect 4480 4682 4508 5162
rect 5400 5158 5428 5706
rect 5388 5152 5440 5158
rect 5388 5094 5440 5100
rect 5676 4954 5704 5706
rect 6044 5090 6072 5706
rect 6492 5696 6544 5702
rect 6492 5638 6544 5644
rect 6124 5628 6176 5634
rect 6124 5570 6176 5576
rect 6032 5084 6084 5090
rect 6032 5026 6084 5032
rect 5664 4948 5716 4954
rect 5664 4890 5716 4896
rect 6044 4682 6072 5026
rect 4468 4676 4520 4682
rect 4468 4618 4520 4624
rect 6032 4676 6084 4682
rect 6032 4618 6084 4624
rect 6136 4546 6164 5570
rect 6308 5560 6360 5566
rect 6308 5502 6360 5508
rect 6124 4540 6176 4546
rect 6124 4482 6176 4488
rect 4008 4404 4060 4410
rect 4008 4346 4060 4352
rect 2720 4064 2772 4070
rect 2720 4006 2772 4012
rect 3272 4064 3324 4070
rect 3272 4006 3324 4012
rect 3284 3594 3312 4006
rect 3364 3928 3416 3934
rect 3364 3870 3416 3876
rect 3272 3588 3324 3594
rect 3272 3530 3324 3536
rect 3376 3390 3404 3870
rect 3916 3860 3968 3866
rect 3916 3802 3968 3808
rect 3504 3692 3824 3712
rect 3504 3690 3516 3692
rect 3572 3690 3596 3692
rect 3652 3690 3676 3692
rect 3732 3690 3756 3692
rect 3812 3690 3824 3692
rect 3504 3638 3510 3690
rect 3572 3638 3574 3690
rect 3754 3638 3756 3690
rect 3818 3638 3824 3690
rect 3504 3636 3516 3638
rect 3572 3636 3596 3638
rect 3652 3636 3676 3638
rect 3732 3636 3756 3638
rect 3812 3636 3824 3638
rect 3504 3616 3824 3636
rect 3928 3594 3956 3802
rect 4020 3594 4048 4346
rect 3916 3588 3968 3594
rect 3916 3530 3968 3536
rect 4008 3588 4060 3594
rect 4008 3530 4060 3536
rect 6136 3390 6164 4482
rect 6216 4336 6268 4342
rect 6216 4278 6268 4284
rect 3364 3384 3416 3390
rect 3364 3326 3416 3332
rect 6124 3384 6176 3390
rect 6124 3326 6176 3332
rect 3272 3248 3324 3254
rect 3376 3236 3404 3326
rect 6228 3254 6256 4278
rect 3324 3208 3404 3236
rect 5112 3248 5164 3254
rect 3272 3190 3324 3196
rect 5112 3190 5164 3196
rect 6216 3248 6268 3254
rect 6216 3190 6268 3196
rect 3088 2160 3140 2166
rect 3088 2102 3140 2108
rect 2536 1820 2588 1826
rect 2536 1762 2588 1768
rect 2168 1752 2220 1758
rect 2168 1694 2220 1700
rect 2352 1752 2404 1758
rect 2352 1694 2404 1700
rect 2364 1418 2392 1694
rect 2076 1412 2128 1418
rect 2352 1412 2404 1418
rect 2076 1354 2128 1360
rect 2272 1372 2352 1400
rect 1616 1140 1668 1146
rect 1616 1082 1668 1088
rect 1628 874 1656 1082
rect 1340 868 1392 874
rect 1340 810 1392 816
rect 1616 868 1668 874
rect 1616 810 1668 816
rect 2272 420 2300 1372
rect 2352 1354 2404 1360
rect 3100 1146 3128 2102
rect 3284 1418 3312 3190
rect 5124 2914 5152 3190
rect 5112 2908 5164 2914
rect 5112 2850 5164 2856
rect 4744 2704 4796 2710
rect 4744 2646 4796 2652
rect 3504 2604 3824 2624
rect 3504 2602 3516 2604
rect 3572 2602 3596 2604
rect 3652 2602 3676 2604
rect 3732 2602 3756 2604
rect 3812 2602 3824 2604
rect 3504 2550 3510 2602
rect 3572 2550 3574 2602
rect 3754 2550 3756 2602
rect 3818 2550 3824 2602
rect 3504 2548 3516 2550
rect 3572 2548 3596 2550
rect 3652 2548 3676 2550
rect 3732 2548 3756 2550
rect 3812 2548 3824 2550
rect 3504 2528 3824 2548
rect 4756 2166 4784 2646
rect 5124 2506 5152 2850
rect 5112 2500 5164 2506
rect 5112 2442 5164 2448
rect 4744 2160 4796 2166
rect 4744 2102 4796 2108
rect 6216 2160 6268 2166
rect 6216 2102 6268 2108
rect 6228 1894 6256 2102
rect 4192 1888 4244 1894
rect 4192 1830 4244 1836
rect 6216 1888 6268 1894
rect 6216 1830 6268 1836
rect 3364 1820 3416 1826
rect 3364 1762 3416 1768
rect 3272 1412 3324 1418
rect 3272 1354 3324 1360
rect 3088 1140 3140 1146
rect 3088 1082 3140 1088
rect 3376 874 3404 1762
rect 3916 1752 3968 1758
rect 3916 1694 3968 1700
rect 3504 1516 3824 1536
rect 3504 1514 3516 1516
rect 3572 1514 3596 1516
rect 3652 1514 3676 1516
rect 3732 1514 3756 1516
rect 3812 1514 3824 1516
rect 3504 1462 3510 1514
rect 3572 1462 3574 1514
rect 3754 1462 3756 1514
rect 3818 1462 3824 1514
rect 3504 1460 3516 1462
rect 3572 1460 3596 1462
rect 3652 1460 3676 1462
rect 3732 1460 3756 1462
rect 3812 1460 3824 1462
rect 3504 1440 3824 1460
rect 3928 1214 3956 1694
rect 4204 1350 4232 1830
rect 5848 1820 5900 1826
rect 5848 1762 5900 1768
rect 4284 1752 4336 1758
rect 4284 1694 4336 1700
rect 4192 1344 4244 1350
rect 4192 1286 4244 1292
rect 3916 1208 3968 1214
rect 3836 1156 3916 1162
rect 3836 1150 3968 1156
rect 3836 1134 3956 1150
rect 3836 874 3864 1134
rect 4296 1078 4324 1694
rect 5860 1214 5888 1762
rect 5848 1208 5900 1214
rect 5848 1150 5900 1156
rect 3916 1072 3968 1078
rect 3916 1014 3968 1020
rect 4284 1072 4336 1078
rect 4284 1014 4336 1020
rect 3928 874 3956 1014
rect 3364 868 3416 874
rect 3364 810 3416 816
rect 3824 868 3876 874
rect 3824 810 3876 816
rect 3916 868 3968 874
rect 3916 810 3968 816
rect 3504 428 3824 448
rect 3504 426 3516 428
rect 3572 426 3596 428
rect 3652 426 3676 428
rect 3732 426 3756 428
rect 3812 426 3824 428
rect 376 0 516 420
rect 2216 0 2356 420
rect 3504 374 3510 426
rect 3572 374 3574 426
rect 3754 374 3756 426
rect 3818 374 3824 426
rect 4296 420 4324 1014
rect 6228 874 6256 1830
rect 6216 868 6268 874
rect 6216 810 6268 816
rect 6320 420 6348 5502
rect 6504 5226 6532 5638
rect 6492 5220 6544 5226
rect 6492 5162 6544 5168
rect 6504 4682 6532 5162
rect 6952 5152 7004 5158
rect 6952 5094 7004 5100
rect 6964 4682 6992 5094
rect 6492 4676 6544 4682
rect 6492 4618 6544 4624
rect 6952 4676 7004 4682
rect 6952 4618 7004 4624
rect 7056 3769 7084 18626
rect 7148 17534 7176 19510
rect 7332 17738 7360 19850
rect 7700 19370 7728 20190
rect 7872 20112 7924 20118
rect 7872 20054 7924 20060
rect 7884 19778 7912 20054
rect 8160 19778 8188 20394
rect 7872 19772 7924 19778
rect 7872 19714 7924 19720
rect 8148 19772 8200 19778
rect 8148 19714 8200 19720
rect 8056 19704 8108 19710
rect 8056 19646 8108 19652
rect 7688 19364 7740 19370
rect 7688 19306 7740 19312
rect 7596 19228 7648 19234
rect 7596 19170 7648 19176
rect 7504 19160 7556 19166
rect 7504 19102 7556 19108
rect 7516 18758 7544 19102
rect 7504 18752 7556 18758
rect 7504 18694 7556 18700
rect 7504 18616 7556 18622
rect 7504 18558 7556 18564
rect 7412 18140 7464 18146
rect 7412 18082 7464 18088
rect 7320 17732 7372 17738
rect 7320 17674 7372 17680
rect 7136 17528 7188 17534
rect 7136 17470 7188 17476
rect 7424 17398 7452 18082
rect 7516 18078 7544 18558
rect 7504 18072 7556 18078
rect 7504 18014 7556 18020
rect 7608 17942 7636 19170
rect 8068 18758 8096 19646
rect 8344 18758 8372 21822
rect 8056 18752 8108 18758
rect 8056 18694 8108 18700
rect 8332 18752 8384 18758
rect 8332 18694 8384 18700
rect 8068 18282 8096 18694
rect 8056 18276 8108 18282
rect 8056 18218 8108 18224
rect 7596 17936 7648 17942
rect 7596 17878 7648 17884
rect 7412 17392 7464 17398
rect 7412 17334 7464 17340
rect 7228 16848 7280 16854
rect 7228 16790 7280 16796
rect 7240 16582 7268 16790
rect 7228 16576 7280 16582
rect 7228 16518 7280 16524
rect 7240 16310 7268 16518
rect 7228 16304 7280 16310
rect 7228 16246 7280 16252
rect 7136 15420 7188 15426
rect 7136 15362 7188 15368
rect 7148 14270 7176 15362
rect 7240 14678 7268 16246
rect 7320 15216 7372 15222
rect 7320 15158 7372 15164
rect 7228 14672 7280 14678
rect 7228 14614 7280 14620
rect 7136 14264 7188 14270
rect 7136 14206 7188 14212
rect 7136 13584 7188 13590
rect 7136 13526 7188 13532
rect 7148 12745 7176 13526
rect 7228 13176 7280 13182
rect 7228 13118 7280 13124
rect 7134 12736 7190 12745
rect 7134 12671 7190 12680
rect 7148 12026 7176 12671
rect 7240 12502 7268 13118
rect 7332 12842 7360 15158
rect 7424 14814 7452 17334
rect 7412 14808 7464 14814
rect 7412 14750 7464 14756
rect 7504 14400 7556 14406
rect 7504 14342 7556 14348
rect 7412 13856 7464 13862
rect 7412 13798 7464 13804
rect 7424 13386 7452 13798
rect 7412 13380 7464 13386
rect 7412 13322 7464 13328
rect 7516 13114 7544 14342
rect 7504 13108 7556 13114
rect 7504 13050 7556 13056
rect 7320 12836 7372 12842
rect 7608 12824 7636 17878
rect 8056 17528 8108 17534
rect 8056 17470 8108 17476
rect 7964 17392 8016 17398
rect 7964 17334 8016 17340
rect 7976 16990 8004 17334
rect 7964 16984 8016 16990
rect 7964 16926 8016 16932
rect 7780 15760 7832 15766
rect 7780 15702 7832 15708
rect 7792 15494 7820 15702
rect 7976 15494 8004 16926
rect 7780 15488 7832 15494
rect 7780 15430 7832 15436
rect 7964 15488 8016 15494
rect 7964 15430 8016 15436
rect 7792 14678 7820 15430
rect 8068 15426 8096 17470
rect 8608 16848 8660 16854
rect 8608 16790 8660 16796
rect 8620 16310 8648 16790
rect 8240 16304 8292 16310
rect 8240 16246 8292 16252
rect 8608 16304 8660 16310
rect 8608 16246 8660 16252
rect 8252 15902 8280 16246
rect 8620 15970 8648 16246
rect 8608 15964 8660 15970
rect 8608 15906 8660 15912
rect 8240 15896 8292 15902
rect 8240 15838 8292 15844
rect 8056 15420 8108 15426
rect 8056 15362 8108 15368
rect 7872 15284 7924 15290
rect 7872 15226 7924 15232
rect 7884 15193 7912 15226
rect 7870 15184 7926 15193
rect 7870 15119 7926 15128
rect 8712 15018 8740 21890
rect 8792 18072 8844 18078
rect 8792 18014 8844 18020
rect 8700 15012 8752 15018
rect 8700 14954 8752 14960
rect 8424 14876 8476 14882
rect 8424 14818 8476 14824
rect 7780 14672 7832 14678
rect 7780 14614 7832 14620
rect 8436 14474 8464 14818
rect 8516 14808 8568 14814
rect 8516 14750 8568 14756
rect 8424 14468 8476 14474
rect 8424 14410 8476 14416
rect 8056 14332 8108 14338
rect 8056 14274 8108 14280
rect 7688 14196 7740 14202
rect 7688 14138 7740 14144
rect 7700 13182 7728 14138
rect 8068 14134 8096 14274
rect 8056 14128 8108 14134
rect 7976 14088 8056 14116
rect 7976 13726 8004 14088
rect 8056 14070 8108 14076
rect 8056 13856 8108 13862
rect 8056 13798 8108 13804
rect 7964 13720 8016 13726
rect 7964 13662 8016 13668
rect 7780 13380 7832 13386
rect 7780 13322 7832 13328
rect 7688 13176 7740 13182
rect 7688 13118 7740 13124
rect 7700 12842 7728 13118
rect 7320 12778 7372 12784
rect 7424 12796 7636 12824
rect 7688 12836 7740 12842
rect 7228 12496 7280 12502
rect 7228 12438 7280 12444
rect 7136 12020 7188 12026
rect 7136 11962 7188 11968
rect 7424 11618 7452 12796
rect 7688 12778 7740 12784
rect 7792 12706 7820 13322
rect 7872 13040 7924 13046
rect 7872 12982 7924 12988
rect 7504 12700 7556 12706
rect 7504 12642 7556 12648
rect 7780 12700 7832 12706
rect 7780 12642 7832 12648
rect 7516 12298 7544 12642
rect 7504 12292 7556 12298
rect 7504 12234 7556 12240
rect 7792 12230 7820 12642
rect 7884 12638 7912 12982
rect 7976 12774 8004 13662
rect 7964 12768 8016 12774
rect 7964 12710 8016 12716
rect 7872 12632 7924 12638
rect 7872 12574 7924 12580
rect 7964 12564 8016 12570
rect 7964 12506 8016 12512
rect 7780 12224 7832 12230
rect 7780 12166 7832 12172
rect 7504 12088 7556 12094
rect 7504 12030 7556 12036
rect 7516 11754 7544 12030
rect 7688 11952 7740 11958
rect 7688 11894 7740 11900
rect 7700 11754 7728 11894
rect 7504 11748 7556 11754
rect 7504 11690 7556 11696
rect 7688 11748 7740 11754
rect 7688 11690 7740 11696
rect 7412 11612 7464 11618
rect 7412 11554 7464 11560
rect 7228 10864 7280 10870
rect 7228 10806 7280 10812
rect 7136 10116 7188 10122
rect 7136 10058 7188 10064
rect 7148 9374 7176 10058
rect 7240 9986 7268 10806
rect 7228 9980 7280 9986
rect 7228 9922 7280 9928
rect 7424 9578 7452 11554
rect 7792 11210 7820 12166
rect 7872 11680 7924 11686
rect 7872 11622 7924 11628
rect 7780 11204 7832 11210
rect 7780 11146 7832 11152
rect 7792 10666 7820 11146
rect 7884 11006 7912 11622
rect 7872 11000 7924 11006
rect 7872 10942 7924 10948
rect 7780 10660 7832 10666
rect 7780 10602 7832 10608
rect 7412 9572 7464 9578
rect 7412 9514 7464 9520
rect 7136 9368 7188 9374
rect 7136 9310 7188 9316
rect 7884 9238 7912 10942
rect 7872 9232 7924 9238
rect 7872 9174 7924 9180
rect 7320 6648 7372 6654
rect 7320 6590 7372 6596
rect 7228 6512 7280 6518
rect 7228 6454 7280 6460
rect 7136 6172 7188 6178
rect 7136 6114 7188 6120
rect 7148 5702 7176 6114
rect 7136 5696 7188 5702
rect 7136 5638 7188 5644
rect 7240 5634 7268 6454
rect 7332 6178 7360 6590
rect 7320 6172 7372 6178
rect 7320 6114 7372 6120
rect 7228 5628 7280 5634
rect 7228 5570 7280 5576
rect 7976 4554 8004 12506
rect 8068 12502 8096 13798
rect 8148 13584 8200 13590
rect 8148 13526 8200 13532
rect 8160 13386 8188 13526
rect 8148 13380 8200 13386
rect 8148 13322 8200 13328
rect 8056 12496 8108 12502
rect 8056 12438 8108 12444
rect 8160 12298 8188 13322
rect 8332 13312 8384 13318
rect 8332 13254 8384 13260
rect 8238 12736 8294 12745
rect 8238 12671 8294 12680
rect 8252 12638 8280 12671
rect 8240 12632 8292 12638
rect 8240 12574 8292 12580
rect 8148 12292 8200 12298
rect 8148 12234 8200 12240
rect 8240 12292 8292 12298
rect 8240 12234 8292 12240
rect 8252 12026 8280 12234
rect 8240 12020 8292 12026
rect 8240 11962 8292 11968
rect 8252 11414 8280 11962
rect 8344 11958 8372 13254
rect 8436 12842 8464 14410
rect 8424 12836 8476 12842
rect 8424 12778 8476 12784
rect 8424 12632 8476 12638
rect 8424 12574 8476 12580
rect 8332 11952 8384 11958
rect 8332 11894 8384 11900
rect 8240 11408 8292 11414
rect 8240 11350 8292 11356
rect 8344 10598 8372 11894
rect 8332 10592 8384 10598
rect 8332 10534 8384 10540
rect 8240 10388 8292 10394
rect 8240 10330 8292 10336
rect 8252 10054 8280 10330
rect 8240 10048 8292 10054
rect 8240 9990 8292 9996
rect 8240 9776 8292 9782
rect 8240 9718 8292 9724
rect 8252 8898 8280 9718
rect 8240 8892 8292 8898
rect 8240 8834 8292 8840
rect 8436 8354 8464 12574
rect 8528 10666 8556 14750
rect 8804 14678 8832 18014
rect 8608 14672 8660 14678
rect 8608 14614 8660 14620
rect 8792 14672 8844 14678
rect 8792 14614 8844 14620
rect 8620 14474 8648 14614
rect 8608 14468 8660 14474
rect 8608 14410 8660 14416
rect 8896 14214 8924 22842
rect 8976 19160 9028 19166
rect 8976 19102 9028 19108
rect 8988 16650 9016 19102
rect 9172 18826 9200 25018
rect 9264 24606 9292 25086
rect 9252 24600 9304 24606
rect 9252 24542 9304 24548
rect 9816 24470 9844 25086
rect 10460 24742 10488 25222
rect 11104 25014 11132 25630
rect 11748 25150 11776 25766
rect 12208 25150 12236 26106
rect 12380 25756 12432 25762
rect 12380 25698 12432 25704
rect 11736 25144 11788 25150
rect 11736 25086 11788 25092
rect 12196 25144 12248 25150
rect 12196 25086 12248 25092
rect 11092 25008 11144 25014
rect 11092 24950 11144 24956
rect 10448 24736 10500 24742
rect 10448 24678 10500 24684
rect 9988 24600 10040 24606
rect 9988 24542 10040 24548
rect 9804 24464 9856 24470
rect 9804 24406 9856 24412
rect 9816 23110 9844 24406
rect 10000 24266 10028 24542
rect 9988 24260 10040 24266
rect 9988 24202 10040 24208
rect 10460 24198 10488 24678
rect 10448 24192 10500 24198
rect 10448 24134 10500 24140
rect 9804 23104 9856 23110
rect 9804 23046 9856 23052
rect 11000 22900 11052 22906
rect 11000 22842 11052 22848
rect 11012 22498 11040 22842
rect 11000 22492 11052 22498
rect 11000 22434 11052 22440
rect 10816 22288 10868 22294
rect 10816 22230 10868 22236
rect 10828 21954 10856 22230
rect 11012 22022 11040 22434
rect 11000 22016 11052 22022
rect 11000 21958 11052 21964
rect 10816 21948 10868 21954
rect 10816 21890 10868 21896
rect 11012 21546 11040 21958
rect 11000 21540 11052 21546
rect 11000 21482 11052 21488
rect 9252 21404 9304 21410
rect 9252 21346 9304 21352
rect 9436 21404 9488 21410
rect 9436 21346 9488 21352
rect 9264 21002 9292 21346
rect 9252 20996 9304 21002
rect 9252 20938 9304 20944
rect 9448 20712 9476 21346
rect 9528 21200 9580 21206
rect 9528 21142 9580 21148
rect 9540 21002 9568 21142
rect 9528 20996 9580 21002
rect 9528 20938 9580 20944
rect 10172 20860 10224 20866
rect 10172 20802 10224 20808
rect 9528 20724 9580 20730
rect 9448 20684 9528 20712
rect 9528 20666 9580 20672
rect 9436 20316 9488 20322
rect 9436 20258 9488 20264
rect 9344 20248 9396 20254
rect 9344 20190 9396 20196
rect 9356 19642 9384 20190
rect 9448 19914 9476 20258
rect 9436 19908 9488 19914
rect 9436 19850 9488 19856
rect 9344 19636 9396 19642
rect 9344 19578 9396 19584
rect 9160 18820 9212 18826
rect 9160 18762 9212 18768
rect 9068 18616 9120 18622
rect 9068 18558 9120 18564
rect 8976 16644 9028 16650
rect 8976 16586 9028 16592
rect 8988 16378 9016 16586
rect 9080 16514 9108 18558
rect 9172 18486 9200 18762
rect 9160 18480 9212 18486
rect 9212 18440 9292 18468
rect 9160 18422 9212 18428
rect 9160 18140 9212 18146
rect 9160 18082 9212 18088
rect 9172 17466 9200 18082
rect 9264 17534 9292 18440
rect 9356 17942 9384 19578
rect 9540 18690 9568 20666
rect 9988 19228 10040 19234
rect 9988 19170 10040 19176
rect 9528 18684 9580 18690
rect 9528 18626 9580 18632
rect 10000 18486 10028 19170
rect 10184 19098 10212 20802
rect 11104 20458 11132 24950
rect 11748 24810 11776 25086
rect 12208 24810 12236 25086
rect 12392 25014 12420 25698
rect 12380 25008 12432 25014
rect 12380 24950 12432 24956
rect 11736 24804 11788 24810
rect 11736 24746 11788 24752
rect 12196 24804 12248 24810
rect 12196 24746 12248 24752
rect 11368 24736 11420 24742
rect 11368 24678 11420 24684
rect 11380 24198 11408 24678
rect 11460 24464 11512 24470
rect 11460 24406 11512 24412
rect 11472 24266 11500 24406
rect 11460 24260 11512 24266
rect 11460 24202 11512 24208
rect 11368 24192 11420 24198
rect 11368 24134 11420 24140
rect 12392 23874 12420 24950
rect 12484 24810 12512 26106
rect 14232 25694 14260 27315
rect 14864 26164 14916 26170
rect 14864 26106 14916 26112
rect 14876 25830 14904 26106
rect 14864 25824 14916 25830
rect 14864 25766 14916 25772
rect 15876 25824 15928 25830
rect 15876 25766 15928 25772
rect 12564 25688 12616 25694
rect 12564 25630 12616 25636
rect 14220 25688 14272 25694
rect 14220 25630 14272 25636
rect 14404 25688 14456 25694
rect 14404 25630 14456 25636
rect 12576 25354 12604 25630
rect 12564 25348 12616 25354
rect 12564 25290 12616 25296
rect 14416 25082 14444 25630
rect 14876 25354 14904 25766
rect 15232 25688 15284 25694
rect 15232 25630 15284 25636
rect 14864 25348 14916 25354
rect 14864 25290 14916 25296
rect 15244 25286 15272 25630
rect 15888 25354 15916 25766
rect 16152 25688 16204 25694
rect 16152 25630 16204 25636
rect 15876 25348 15928 25354
rect 15876 25290 15928 25296
rect 15232 25280 15284 25286
rect 15232 25222 15284 25228
rect 14956 25144 15008 25150
rect 14956 25086 15008 25092
rect 12564 25076 12616 25082
rect 12564 25018 12616 25024
rect 14404 25076 14456 25082
rect 14404 25018 14456 25024
rect 12472 24804 12524 24810
rect 12472 24746 12524 24752
rect 12484 24266 12512 24746
rect 12576 24674 12604 25018
rect 12564 24668 12616 24674
rect 12564 24610 12616 24616
rect 12576 24266 12604 24610
rect 12472 24260 12524 24266
rect 12472 24202 12524 24208
rect 12564 24260 12616 24266
rect 12564 24202 12616 24208
rect 14416 24062 14444 25018
rect 14968 24674 14996 25086
rect 14956 24668 15008 24674
rect 14956 24610 15008 24616
rect 14404 24056 14456 24062
rect 14404 23998 14456 24004
rect 12392 23846 12512 23874
rect 12484 23654 12512 23846
rect 14968 23722 14996 24610
rect 15140 24600 15192 24606
rect 15140 24542 15192 24548
rect 15152 24130 15180 24542
rect 15140 24124 15192 24130
rect 15140 24066 15192 24072
rect 15152 23994 15180 24066
rect 15140 23988 15192 23994
rect 15140 23930 15192 23936
rect 15152 23722 15180 23930
rect 14956 23716 15008 23722
rect 14956 23658 15008 23664
rect 15140 23716 15192 23722
rect 15140 23658 15192 23664
rect 12472 23648 12524 23654
rect 12472 23590 12524 23596
rect 12484 23525 12512 23590
rect 13392 23580 13444 23586
rect 13392 23522 13444 23528
rect 15968 23580 16020 23586
rect 15968 23522 16020 23528
rect 12288 23512 12340 23518
rect 12288 23454 12340 23460
rect 12564 23512 12616 23518
rect 12564 23454 12616 23460
rect 11828 23036 11880 23042
rect 11828 22978 11880 22984
rect 11368 22492 11420 22498
rect 11368 22434 11420 22440
rect 11380 22090 11408 22434
rect 11368 22084 11420 22090
rect 11368 22026 11420 22032
rect 11736 21880 11788 21886
rect 11736 21822 11788 21828
rect 11092 20452 11144 20458
rect 11092 20394 11144 20400
rect 10264 20384 10316 20390
rect 10264 20326 10316 20332
rect 10276 19914 10304 20326
rect 10264 19908 10316 19914
rect 10264 19850 10316 19856
rect 11092 19228 11144 19234
rect 11092 19170 11144 19176
rect 10816 19160 10868 19166
rect 10816 19102 10868 19108
rect 11000 19160 11052 19166
rect 11000 19102 11052 19108
rect 10172 19092 10224 19098
rect 10172 19034 10224 19040
rect 9988 18480 10040 18486
rect 9988 18422 10040 18428
rect 10000 18185 10028 18422
rect 10184 18282 10212 19034
rect 10828 18486 10856 19102
rect 11012 18826 11040 19102
rect 11000 18820 11052 18826
rect 11000 18762 11052 18768
rect 11000 18548 11052 18554
rect 11104 18536 11132 19170
rect 11052 18508 11132 18536
rect 11000 18490 11052 18496
rect 10816 18480 10868 18486
rect 10816 18422 10868 18428
rect 10172 18276 10224 18282
rect 10172 18218 10224 18224
rect 9986 18176 10042 18185
rect 9436 18140 9488 18146
rect 9986 18111 10042 18120
rect 9436 18082 9488 18088
rect 9344 17936 9396 17942
rect 9344 17878 9396 17884
rect 9252 17528 9304 17534
rect 9252 17470 9304 17476
rect 9160 17460 9212 17466
rect 9160 17402 9212 17408
rect 9356 17194 9384 17878
rect 9448 17398 9476 18082
rect 10828 17942 10856 18422
rect 11012 18146 11040 18490
rect 11000 18140 11052 18146
rect 11000 18082 11052 18088
rect 10816 17936 10868 17942
rect 10816 17878 10868 17884
rect 9804 17732 9856 17738
rect 9804 17674 9856 17680
rect 9436 17392 9488 17398
rect 9436 17334 9488 17340
rect 9344 17188 9396 17194
rect 9344 17130 9396 17136
rect 9068 16508 9120 16514
rect 9068 16450 9120 16456
rect 8976 16372 9028 16378
rect 8976 16314 9028 16320
rect 9080 16106 9108 16450
rect 9344 16372 9396 16378
rect 9344 16314 9396 16320
rect 9356 16106 9384 16314
rect 9068 16100 9120 16106
rect 9068 16042 9120 16048
rect 9344 16100 9396 16106
rect 9344 16042 9396 16048
rect 9160 15896 9212 15902
rect 9160 15838 9212 15844
rect 9172 15222 9200 15838
rect 9356 15494 9384 16042
rect 9344 15488 9396 15494
rect 9344 15430 9396 15436
rect 9160 15216 9212 15222
rect 9160 15158 9212 15164
rect 8976 14876 9028 14882
rect 8976 14818 9028 14824
rect 9068 14876 9120 14882
rect 9068 14818 9120 14824
rect 8988 14474 9016 14818
rect 8976 14468 9028 14474
rect 8976 14410 9028 14416
rect 9080 14406 9108 14818
rect 9068 14400 9120 14406
rect 9068 14342 9120 14348
rect 8896 14186 9016 14214
rect 8608 13652 8660 13658
rect 8608 13594 8660 13600
rect 8620 13182 8648 13594
rect 8884 13312 8936 13318
rect 8884 13254 8936 13260
rect 8608 13176 8660 13182
rect 8608 13118 8660 13124
rect 8792 13176 8844 13182
rect 8792 13118 8844 13124
rect 8620 11550 8648 13118
rect 8804 12026 8832 13118
rect 8896 13046 8924 13254
rect 8884 13040 8936 13046
rect 8884 12982 8936 12988
rect 8792 12020 8844 12026
rect 8792 11962 8844 11968
rect 8804 11754 8832 11962
rect 8792 11748 8844 11754
rect 8792 11690 8844 11696
rect 8608 11544 8660 11550
rect 8608 11486 8660 11492
rect 8620 11006 8648 11486
rect 8896 11074 8924 12982
rect 8988 11464 9016 14186
rect 9172 13658 9200 15158
rect 9356 14814 9384 15430
rect 9344 14808 9396 14814
rect 9344 14750 9396 14756
rect 9448 14678 9476 17334
rect 9816 16990 9844 17674
rect 10828 17534 10856 17878
rect 9896 17528 9948 17534
rect 9896 17470 9948 17476
rect 10816 17528 10868 17534
rect 10816 17470 10868 17476
rect 9804 16984 9856 16990
rect 9804 16926 9856 16932
rect 9528 16032 9580 16038
rect 9528 15974 9580 15980
rect 9540 15494 9568 15974
rect 9712 15964 9764 15970
rect 9712 15906 9764 15912
rect 9620 15828 9672 15834
rect 9620 15770 9672 15776
rect 9632 15562 9660 15770
rect 9620 15556 9672 15562
rect 9620 15498 9672 15504
rect 9528 15488 9580 15494
rect 9528 15430 9580 15436
rect 9344 14672 9396 14678
rect 9344 14614 9396 14620
rect 9436 14672 9488 14678
rect 9436 14614 9488 14620
rect 9356 14474 9384 14614
rect 9540 14474 9568 15430
rect 9724 15222 9752 15906
rect 9804 15896 9856 15902
rect 9804 15838 9856 15844
rect 9816 15562 9844 15838
rect 9804 15556 9856 15562
rect 9804 15498 9856 15504
rect 9712 15216 9764 15222
rect 9712 15158 9764 15164
rect 9620 15012 9672 15018
rect 9620 14954 9672 14960
rect 9344 14468 9396 14474
rect 9344 14410 9396 14416
rect 9528 14468 9580 14474
rect 9528 14410 9580 14416
rect 9528 14264 9580 14270
rect 9528 14206 9580 14212
rect 9344 14128 9396 14134
rect 9344 14070 9396 14076
rect 9160 13652 9212 13658
rect 9160 13594 9212 13600
rect 9252 13584 9304 13590
rect 9252 13526 9304 13532
rect 9264 13182 9292 13526
rect 9252 13176 9304 13182
rect 9252 13118 9304 13124
rect 9356 11618 9384 14070
rect 9540 13969 9568 14206
rect 9526 13960 9582 13969
rect 9526 13895 9582 13904
rect 9540 13726 9568 13895
rect 9528 13720 9580 13726
rect 9528 13662 9580 13668
rect 9436 12700 9488 12706
rect 9436 12642 9488 12648
rect 9344 11612 9396 11618
rect 9344 11554 9396 11560
rect 8988 11436 9200 11464
rect 8884 11068 8936 11074
rect 8884 11010 8936 11016
rect 8608 11000 8660 11006
rect 8608 10942 8660 10948
rect 8516 10660 8568 10666
rect 8516 10602 8568 10608
rect 8528 10122 8556 10602
rect 8516 10116 8568 10122
rect 8516 10058 8568 10064
rect 8620 9850 8648 10942
rect 8700 10932 8752 10938
rect 8700 10874 8752 10880
rect 8712 10462 8740 10874
rect 9068 10864 9120 10870
rect 9068 10806 9120 10812
rect 9080 10598 9108 10806
rect 8792 10592 8844 10598
rect 8792 10534 8844 10540
rect 9068 10592 9120 10598
rect 9068 10534 9120 10540
rect 8700 10456 8752 10462
rect 8700 10398 8752 10404
rect 8712 9918 8740 10398
rect 8804 10054 8832 10534
rect 9080 10122 9108 10534
rect 9068 10116 9120 10122
rect 9068 10058 9120 10064
rect 8792 10048 8844 10054
rect 8792 9990 8844 9996
rect 9068 9980 9120 9986
rect 9068 9922 9120 9928
rect 8700 9912 8752 9918
rect 8700 9854 8752 9860
rect 8884 9912 8936 9918
rect 8884 9854 8936 9860
rect 8608 9844 8660 9850
rect 8608 9786 8660 9792
rect 8896 9782 8924 9854
rect 8516 9776 8568 9782
rect 8516 9718 8568 9724
rect 8884 9776 8936 9782
rect 8884 9718 8936 9724
rect 8528 8762 8556 9718
rect 8608 9300 8660 9306
rect 8608 9242 8660 9248
rect 8516 8756 8568 8762
rect 8516 8698 8568 8704
rect 8424 8348 8476 8354
rect 8424 8290 8476 8296
rect 8436 7334 8464 8290
rect 8424 7328 8476 7334
rect 8424 7270 8476 7276
rect 8620 6858 8648 9242
rect 8896 8966 8924 9718
rect 9080 9442 9108 9922
rect 9068 9436 9120 9442
rect 9068 9378 9120 9384
rect 9080 9034 9108 9378
rect 9068 9028 9120 9034
rect 9068 8970 9120 8976
rect 8884 8960 8936 8966
rect 8884 8902 8936 8908
rect 8896 7266 8924 8902
rect 9068 8892 9120 8898
rect 9068 8834 9120 8840
rect 9080 8490 9108 8834
rect 9068 8484 9120 8490
rect 9068 8426 9120 8432
rect 8976 8348 9028 8354
rect 8976 8290 9028 8296
rect 8988 7878 9016 8290
rect 9080 8286 9108 8426
rect 9068 8280 9120 8286
rect 9068 8222 9120 8228
rect 9080 7946 9108 8222
rect 9068 7940 9120 7946
rect 9068 7882 9120 7888
rect 8976 7872 9028 7878
rect 8976 7814 9028 7820
rect 8884 7260 8936 7266
rect 8884 7202 8936 7208
rect 8896 6858 8924 7202
rect 8608 6852 8660 6858
rect 8608 6794 8660 6800
rect 8884 6852 8936 6858
rect 8884 6794 8936 6800
rect 8620 6654 8648 6794
rect 8608 6648 8660 6654
rect 8608 6590 8660 6596
rect 8620 5226 8648 6590
rect 8976 6172 9028 6178
rect 8976 6114 9028 6120
rect 8700 5968 8752 5974
rect 8700 5910 8752 5916
rect 8712 5566 8740 5910
rect 8988 5634 9016 6114
rect 8976 5628 9028 5634
rect 8976 5570 9028 5576
rect 8700 5560 8752 5566
rect 8700 5502 8752 5508
rect 8608 5220 8660 5226
rect 8608 5162 8660 5168
rect 7976 4526 8188 4554
rect 7042 3760 7098 3769
rect 7042 3695 7098 3704
rect 6676 2908 6728 2914
rect 6676 2850 6728 2856
rect 6688 2506 6716 2850
rect 7504 2840 7556 2846
rect 7504 2782 7556 2788
rect 7136 2704 7188 2710
rect 7136 2646 7188 2652
rect 6676 2500 6728 2506
rect 6676 2442 6728 2448
rect 6688 2302 6716 2442
rect 7148 2438 7176 2646
rect 7136 2432 7188 2438
rect 7136 2374 7188 2380
rect 6676 2296 6728 2302
rect 6676 2238 6728 2244
rect 7148 1894 7176 2374
rect 7516 1962 7544 2782
rect 7780 2296 7832 2302
rect 7780 2238 7832 2244
rect 7504 1956 7556 1962
rect 7504 1898 7556 1904
rect 7136 1888 7188 1894
rect 7136 1830 7188 1836
rect 6584 1820 6636 1826
rect 6584 1762 6636 1768
rect 6596 1146 6624 1762
rect 7516 1282 7544 1898
rect 7792 1826 7820 2238
rect 8160 1826 8188 4526
rect 8712 4410 8740 5502
rect 8988 5498 9016 5570
rect 8976 5492 9028 5498
rect 8976 5434 9028 5440
rect 8988 5226 9016 5434
rect 8976 5220 9028 5226
rect 8976 5162 9028 5168
rect 9068 5084 9120 5090
rect 9068 5026 9120 5032
rect 8700 4404 8752 4410
rect 8700 4346 8752 4352
rect 8712 3594 8740 4346
rect 9080 4342 9108 5026
rect 9068 4336 9120 4342
rect 9068 4278 9120 4284
rect 9172 4002 9200 11436
rect 9356 10938 9384 11554
rect 9448 11142 9476 12642
rect 9540 12638 9568 13662
rect 9528 12632 9580 12638
rect 9528 12574 9580 12580
rect 9528 12496 9580 12502
rect 9528 12438 9580 12444
rect 9540 11686 9568 12438
rect 9528 11680 9580 11686
rect 9528 11622 9580 11628
rect 9436 11136 9488 11142
rect 9436 11078 9488 11084
rect 9540 11006 9568 11622
rect 9632 11142 9660 14954
rect 9724 13930 9752 15158
rect 9804 14672 9856 14678
rect 9804 14614 9856 14620
rect 9712 13924 9764 13930
rect 9712 13866 9764 13872
rect 9816 13318 9844 14614
rect 9804 13312 9856 13318
rect 9804 13254 9856 13260
rect 9816 13182 9844 13254
rect 9804 13176 9856 13182
rect 9804 13118 9856 13124
rect 9712 13040 9764 13046
rect 9712 12982 9764 12988
rect 9724 12842 9752 12982
rect 9712 12836 9764 12842
rect 9712 12778 9764 12784
rect 9712 11544 9764 11550
rect 9712 11486 9764 11492
rect 9620 11136 9672 11142
rect 9620 11078 9672 11084
rect 9724 11074 9752 11486
rect 9712 11068 9764 11074
rect 9712 11010 9764 11016
rect 9528 11000 9580 11006
rect 9528 10942 9580 10948
rect 9344 10932 9396 10938
rect 9344 10874 9396 10880
rect 9436 10592 9488 10598
rect 9436 10534 9488 10540
rect 9252 10524 9304 10530
rect 9252 10466 9304 10472
rect 9264 9918 9292 10466
rect 9252 9912 9304 9918
rect 9252 9854 9304 9860
rect 9344 9844 9396 9850
rect 9344 9786 9396 9792
rect 9356 9578 9384 9786
rect 9448 9782 9476 10534
rect 9540 10394 9568 10942
rect 9528 10388 9580 10394
rect 9528 10330 9580 10336
rect 9436 9776 9488 9782
rect 9436 9718 9488 9724
rect 9344 9572 9396 9578
rect 9344 9514 9396 9520
rect 9344 9300 9396 9306
rect 9344 9242 9396 9248
rect 9252 9232 9304 9238
rect 9252 9174 9304 9180
rect 9264 9034 9292 9174
rect 9356 9034 9384 9242
rect 9252 9028 9304 9034
rect 9252 8970 9304 8976
rect 9344 9028 9396 9034
rect 9344 8970 9396 8976
rect 9908 7402 9936 17470
rect 9988 17460 10040 17466
rect 9988 17402 10040 17408
rect 10000 15902 10028 17402
rect 11012 17398 11040 18082
rect 11000 17392 11052 17398
rect 11000 17334 11052 17340
rect 10264 17052 10316 17058
rect 10264 16994 10316 17000
rect 10276 16310 10304 16994
rect 10908 16984 10960 16990
rect 10908 16926 10960 16932
rect 10920 16310 10948 16926
rect 11552 16916 11604 16922
rect 11552 16858 11604 16864
rect 11184 16508 11236 16514
rect 11184 16450 11236 16456
rect 11196 16310 11224 16450
rect 10264 16304 10316 16310
rect 10264 16246 10316 16252
rect 10908 16304 10960 16310
rect 10908 16246 10960 16252
rect 11184 16304 11236 16310
rect 11184 16246 11236 16252
rect 11460 16304 11512 16310
rect 11460 16246 11512 16252
rect 9988 15896 10040 15902
rect 9988 15838 10040 15844
rect 9988 14468 10040 14474
rect 9988 14410 10040 14416
rect 10000 14270 10028 14410
rect 10080 14400 10132 14406
rect 10080 14342 10132 14348
rect 10172 14400 10224 14406
rect 10172 14342 10224 14348
rect 9988 14264 10040 14270
rect 9988 14206 10040 14212
rect 10092 13930 10120 14342
rect 10184 14105 10212 14342
rect 10170 14096 10226 14105
rect 10170 14031 10226 14040
rect 10080 13924 10132 13930
rect 10080 13866 10132 13872
rect 9988 13856 10040 13862
rect 9988 13798 10040 13804
rect 10000 13726 10028 13798
rect 10080 13788 10132 13794
rect 10080 13730 10132 13736
rect 9988 13720 10040 13726
rect 9988 13662 10040 13668
rect 10000 13182 10028 13662
rect 10092 13386 10120 13730
rect 10080 13380 10132 13386
rect 10080 13322 10132 13328
rect 9988 13176 10040 13182
rect 9988 13118 10040 13124
rect 10000 12298 10028 13118
rect 9988 12292 10040 12298
rect 9988 12234 10040 12240
rect 10184 11754 10212 14031
rect 10172 11748 10224 11754
rect 10172 11690 10224 11696
rect 10184 11618 10212 11690
rect 10172 11612 10224 11618
rect 10172 11554 10224 11560
rect 10184 11210 10212 11554
rect 10172 11204 10224 11210
rect 10172 11146 10224 11152
rect 10184 11074 10212 11146
rect 10172 11068 10224 11074
rect 10172 11010 10224 11016
rect 9896 7396 9948 7402
rect 9896 7338 9948 7344
rect 9620 7260 9672 7266
rect 9620 7202 9672 7208
rect 9896 7260 9948 7266
rect 9896 7202 9948 7208
rect 9528 7192 9580 7198
rect 9528 7134 9580 7140
rect 9252 7124 9304 7130
rect 9252 7066 9304 7072
rect 9264 6858 9292 7066
rect 9540 6858 9568 7134
rect 9252 6852 9304 6858
rect 9252 6794 9304 6800
rect 9528 6852 9580 6858
rect 9528 6794 9580 6800
rect 9540 5770 9568 6794
rect 9632 6790 9660 7202
rect 9620 6784 9672 6790
rect 9620 6726 9672 6732
rect 9908 6654 9936 7202
rect 10080 7192 10132 7198
rect 10080 7134 10132 7140
rect 10092 6722 10120 7134
rect 10080 6716 10132 6722
rect 10132 6676 10212 6704
rect 10080 6658 10132 6664
rect 9896 6648 9948 6654
rect 9896 6590 9948 6596
rect 9804 6580 9856 6586
rect 9804 6522 9856 6528
rect 9816 6110 9844 6522
rect 9804 6104 9856 6110
rect 9804 6046 9856 6052
rect 9528 5764 9580 5770
rect 9528 5706 9580 5712
rect 9436 5492 9488 5498
rect 9436 5434 9488 5440
rect 9448 5158 9476 5434
rect 9816 5226 9844 6046
rect 9804 5220 9856 5226
rect 9804 5162 9856 5168
rect 9436 5152 9488 5158
rect 9436 5094 9488 5100
rect 9448 4682 9476 5094
rect 9436 4676 9488 4682
rect 9436 4618 9488 4624
rect 10184 4546 10212 6676
rect 10172 4540 10224 4546
rect 10172 4482 10224 4488
rect 9160 3996 9212 4002
rect 9080 3956 9160 3984
rect 8700 3588 8752 3594
rect 8700 3530 8752 3536
rect 9080 3526 9108 3956
rect 9160 3938 9212 3944
rect 9160 3792 9212 3798
rect 9160 3734 9212 3740
rect 9068 3520 9120 3526
rect 9068 3462 9120 3468
rect 9080 3050 9108 3462
rect 9172 3390 9200 3734
rect 9160 3384 9212 3390
rect 9160 3326 9212 3332
rect 9068 3044 9120 3050
rect 9068 2986 9120 2992
rect 9804 2160 9856 2166
rect 9804 2102 9856 2108
rect 9816 1894 9844 2102
rect 8884 1888 8936 1894
rect 8884 1830 8936 1836
rect 9804 1888 9856 1894
rect 9804 1830 9856 1836
rect 7780 1820 7832 1826
rect 7780 1762 7832 1768
rect 8148 1820 8200 1826
rect 8148 1762 8200 1768
rect 7596 1616 7648 1622
rect 7596 1558 7648 1564
rect 7608 1418 7636 1558
rect 7596 1412 7648 1418
rect 7792 1400 7820 1762
rect 8896 1418 8924 1830
rect 10184 1826 10212 4482
rect 10276 2914 10304 16246
rect 10724 14808 10776 14814
rect 10724 14750 10776 14756
rect 10632 14672 10684 14678
rect 10632 14614 10684 14620
rect 10448 14264 10500 14270
rect 10644 14241 10672 14614
rect 10736 14474 10764 14750
rect 10724 14468 10776 14474
rect 10724 14410 10776 14416
rect 10736 14270 10764 14410
rect 10920 14270 10948 16246
rect 10724 14264 10776 14270
rect 10448 14206 10500 14212
rect 10630 14232 10686 14241
rect 10356 14196 10408 14202
rect 10356 14138 10408 14144
rect 10368 13862 10396 14138
rect 10356 13856 10408 13862
rect 10356 13798 10408 13804
rect 10368 13046 10396 13798
rect 10460 13794 10488 14206
rect 10724 14206 10776 14212
rect 10908 14264 10960 14270
rect 10908 14206 10960 14212
rect 10630 14167 10686 14176
rect 10644 14105 10672 14167
rect 10630 14096 10686 14105
rect 10630 14031 10686 14040
rect 10540 13856 10592 13862
rect 10540 13798 10592 13804
rect 10448 13788 10500 13794
rect 10448 13730 10500 13736
rect 10552 13386 10580 13798
rect 10540 13380 10592 13386
rect 10540 13322 10592 13328
rect 10356 13040 10408 13046
rect 10356 12982 10408 12988
rect 10368 9986 10396 12982
rect 11000 12700 11052 12706
rect 11000 12642 11052 12648
rect 10816 12632 10868 12638
rect 10816 12574 10868 12580
rect 10828 11958 10856 12574
rect 11012 12230 11040 12642
rect 11000 12224 11052 12230
rect 11000 12166 11052 12172
rect 10816 11952 10868 11958
rect 10816 11894 10868 11900
rect 10828 11754 10856 11894
rect 10816 11748 10868 11754
rect 10816 11690 10868 11696
rect 10828 11210 10856 11690
rect 11196 11414 11224 16246
rect 11472 16038 11500 16246
rect 11460 16032 11512 16038
rect 11460 15974 11512 15980
rect 11368 15964 11420 15970
rect 11368 15906 11420 15912
rect 11380 15562 11408 15906
rect 11564 15766 11592 16858
rect 11748 16378 11776 21822
rect 11840 21410 11868 22978
rect 12012 22968 12064 22974
rect 12012 22910 12064 22916
rect 12024 22838 12052 22910
rect 12300 22838 12328 23454
rect 12576 22974 12604 23454
rect 13404 23178 13432 23522
rect 13392 23172 13444 23178
rect 13392 23114 13444 23120
rect 12564 22968 12616 22974
rect 12564 22910 12616 22916
rect 13484 22968 13536 22974
rect 13484 22910 13536 22916
rect 15876 22968 15928 22974
rect 15876 22910 15928 22916
rect 13116 22900 13168 22906
rect 13116 22842 13168 22848
rect 12012 22832 12064 22838
rect 12012 22774 12064 22780
rect 12288 22832 12340 22838
rect 12288 22774 12340 22780
rect 12024 22498 12052 22774
rect 12012 22492 12064 22498
rect 12012 22434 12064 22440
rect 11920 21472 11972 21478
rect 11920 21414 11972 21420
rect 11828 21404 11880 21410
rect 11828 21346 11880 21352
rect 11840 20662 11868 21346
rect 11932 20730 11960 21414
rect 12104 21336 12156 21342
rect 12104 21278 12156 21284
rect 12116 20934 12144 21278
rect 12196 21268 12248 21274
rect 12196 21210 12248 21216
rect 12208 21002 12236 21210
rect 12196 20996 12248 21002
rect 12196 20938 12248 20944
rect 12104 20928 12156 20934
rect 12104 20870 12156 20876
rect 11920 20724 11972 20730
rect 11920 20666 11972 20672
rect 11828 20656 11880 20662
rect 11828 20598 11880 20604
rect 11840 19234 11868 20598
rect 11828 19228 11880 19234
rect 11828 19170 11880 19176
rect 11828 16440 11880 16446
rect 11828 16382 11880 16388
rect 11736 16372 11788 16378
rect 11736 16314 11788 16320
rect 11840 15834 11868 16382
rect 11828 15828 11880 15834
rect 11828 15770 11880 15776
rect 11552 15760 11604 15766
rect 11552 15702 11604 15708
rect 11564 15562 11592 15702
rect 11368 15556 11420 15562
rect 11368 15498 11420 15504
rect 11552 15556 11604 15562
rect 11552 15498 11604 15504
rect 11380 14474 11408 15498
rect 11644 14876 11696 14882
rect 11644 14818 11696 14824
rect 11552 14740 11604 14746
rect 11552 14682 11604 14688
rect 11368 14468 11420 14474
rect 11368 14410 11420 14416
rect 11564 14406 11592 14682
rect 11552 14400 11604 14406
rect 11552 14342 11604 14348
rect 11276 14332 11328 14338
rect 11276 14274 11328 14280
rect 11460 14332 11512 14338
rect 11460 14274 11512 14280
rect 11288 13794 11316 14274
rect 11276 13788 11328 13794
rect 11276 13730 11328 13736
rect 11288 13318 11316 13730
rect 11472 13658 11500 14274
rect 11552 14264 11604 14270
rect 11552 14206 11604 14212
rect 11656 14214 11684 14818
rect 11736 14672 11788 14678
rect 11788 14632 11868 14660
rect 11736 14614 11788 14620
rect 11460 13652 11512 13658
rect 11460 13594 11512 13600
rect 11276 13312 11328 13318
rect 11276 13254 11328 13260
rect 11564 13182 11592 14206
rect 11656 14202 11776 14214
rect 11656 14196 11788 14202
rect 11656 14186 11736 14196
rect 11736 14138 11788 14144
rect 11644 13584 11696 13590
rect 11644 13526 11696 13532
rect 11552 13176 11604 13182
rect 11552 13118 11604 13124
rect 11656 13114 11684 13526
rect 11644 13108 11696 13114
rect 11644 13050 11696 13056
rect 11460 12700 11512 12706
rect 11460 12642 11512 12648
rect 11276 12564 11328 12570
rect 11276 12506 11328 12512
rect 11288 11958 11316 12506
rect 11472 12298 11500 12642
rect 11460 12292 11512 12298
rect 11460 12234 11512 12240
rect 11460 12088 11512 12094
rect 11460 12030 11512 12036
rect 11276 11952 11328 11958
rect 11276 11894 11328 11900
rect 11184 11408 11236 11414
rect 11184 11350 11236 11356
rect 10816 11204 10868 11210
rect 10816 11146 10868 11152
rect 11288 11006 11316 11894
rect 11276 11000 11328 11006
rect 11276 10942 11328 10948
rect 11184 10932 11236 10938
rect 11184 10874 11236 10880
rect 10356 9980 10408 9986
rect 10356 9922 10408 9928
rect 11196 9442 11224 10874
rect 11184 9436 11236 9442
rect 11184 9378 11236 9384
rect 11092 9368 11144 9374
rect 11092 9310 11144 9316
rect 11104 9034 11132 9310
rect 11092 9028 11144 9034
rect 11092 8970 11144 8976
rect 11196 8898 11224 9378
rect 11288 9238 11316 10942
rect 11472 10122 11500 12030
rect 11644 11408 11696 11414
rect 11644 11350 11696 11356
rect 11460 10116 11512 10122
rect 11460 10058 11512 10064
rect 11276 9232 11328 9238
rect 11276 9174 11328 9180
rect 11184 8892 11236 8898
rect 11184 8834 11236 8840
rect 11196 7266 11224 8834
rect 11288 8830 11316 9174
rect 11460 9028 11512 9034
rect 11460 8970 11512 8976
rect 11276 8824 11328 8830
rect 11276 8766 11328 8772
rect 11368 8756 11420 8762
rect 11368 8698 11420 8704
rect 11380 8422 11408 8698
rect 11368 8416 11420 8422
rect 11368 8358 11420 8364
rect 11380 7606 11408 8358
rect 11472 8354 11500 8970
rect 11460 8348 11512 8354
rect 11460 8290 11512 8296
rect 11472 7946 11500 8290
rect 11460 7940 11512 7946
rect 11460 7882 11512 7888
rect 11368 7600 11420 7606
rect 11368 7542 11420 7548
rect 11184 7260 11236 7266
rect 11184 7202 11236 7208
rect 10356 6852 10408 6858
rect 10356 6794 10408 6800
rect 10368 6518 10396 6794
rect 11196 6790 11224 7202
rect 11380 7062 11408 7542
rect 11368 7056 11420 7062
rect 11368 6998 11420 7004
rect 11184 6784 11236 6790
rect 11184 6726 11236 6732
rect 10724 6648 10776 6654
rect 10724 6590 10776 6596
rect 10356 6512 10408 6518
rect 10356 6454 10408 6460
rect 10368 6314 10396 6454
rect 10356 6308 10408 6314
rect 10356 6250 10408 6256
rect 10368 5158 10396 6250
rect 10736 6178 10764 6590
rect 11196 6314 11224 6726
rect 11380 6518 11408 6998
rect 11368 6512 11420 6518
rect 11368 6454 11420 6460
rect 11184 6308 11236 6314
rect 11184 6250 11236 6256
rect 10724 6172 10776 6178
rect 10724 6114 10776 6120
rect 10736 5634 10764 6114
rect 10724 5628 10776 5634
rect 10724 5570 10776 5576
rect 10736 5226 10764 5570
rect 11380 5566 11408 6454
rect 11368 5560 11420 5566
rect 11368 5502 11420 5508
rect 11184 5492 11236 5498
rect 11184 5434 11236 5440
rect 10724 5220 10776 5226
rect 10724 5162 10776 5168
rect 11196 5158 11224 5434
rect 10356 5152 10408 5158
rect 10356 5094 10408 5100
rect 11184 5152 11236 5158
rect 11184 5094 11236 5100
rect 10908 5016 10960 5022
rect 10908 4958 10960 4964
rect 10920 4410 10948 4958
rect 11196 4682 11224 5094
rect 11184 4676 11236 4682
rect 11184 4618 11236 4624
rect 10908 4404 10960 4410
rect 10908 4346 10960 4352
rect 11368 3248 11420 3254
rect 11368 3190 11420 3196
rect 10264 2908 10316 2914
rect 10264 2850 10316 2856
rect 10816 2704 10868 2710
rect 10816 2646 10868 2652
rect 10828 2234 10856 2646
rect 11276 2296 11328 2302
rect 11380 2284 11408 3190
rect 11328 2256 11408 2284
rect 11276 2238 11328 2244
rect 10816 2228 10868 2234
rect 10816 2170 10868 2176
rect 10828 1962 10856 2170
rect 10908 2160 10960 2166
rect 10908 2102 10960 2108
rect 10816 1956 10868 1962
rect 10816 1898 10868 1904
rect 9712 1820 9764 1826
rect 9712 1762 9764 1768
rect 9896 1820 9948 1826
rect 9896 1762 9948 1768
rect 10172 1820 10224 1826
rect 10172 1762 10224 1768
rect 9724 1418 9752 1762
rect 7872 1412 7924 1418
rect 7792 1372 7872 1400
rect 7596 1354 7648 1360
rect 7872 1354 7924 1360
rect 8884 1412 8936 1418
rect 8884 1354 8936 1360
rect 9712 1412 9764 1418
rect 9712 1354 9764 1360
rect 9908 1282 9936 1762
rect 10920 1758 10948 2102
rect 11380 1894 11408 2256
rect 11368 1888 11420 1894
rect 11368 1830 11420 1836
rect 9988 1752 10040 1758
rect 9988 1694 10040 1700
rect 10908 1752 10960 1758
rect 10908 1694 10960 1700
rect 7504 1276 7556 1282
rect 7504 1218 7556 1224
rect 8332 1276 8384 1282
rect 8332 1218 8384 1224
rect 9896 1276 9948 1282
rect 9896 1218 9948 1224
rect 6584 1140 6636 1146
rect 6584 1082 6636 1088
rect 8344 420 8372 1218
rect 9908 1078 9936 1218
rect 10000 1214 10028 1694
rect 10920 1418 10948 1694
rect 10908 1412 10960 1418
rect 10908 1354 10960 1360
rect 11380 1282 11408 1830
rect 11460 1752 11512 1758
rect 11460 1694 11512 1700
rect 11472 1418 11500 1694
rect 11460 1412 11512 1418
rect 11460 1354 11512 1360
rect 11368 1276 11420 1282
rect 11368 1218 11420 1224
rect 9988 1208 10040 1214
rect 9988 1150 10040 1156
rect 9896 1072 9948 1078
rect 9896 1014 9948 1020
rect 10000 423 10028 1150
rect 11656 602 11684 11350
rect 11748 11074 11776 14138
rect 11840 14134 11868 14632
rect 11828 14128 11880 14134
rect 11828 14070 11880 14076
rect 11840 13658 11868 14070
rect 11828 13652 11880 13658
rect 11828 13594 11880 13600
rect 11736 11068 11788 11074
rect 11736 11010 11788 11016
rect 11932 9356 11960 20666
rect 12012 18616 12064 18622
rect 12012 18558 12064 18564
rect 12024 15018 12052 18558
rect 12196 18480 12248 18486
rect 12196 18422 12248 18428
rect 12208 17398 12236 18422
rect 12196 17392 12248 17398
rect 12196 17334 12248 17340
rect 12208 17058 12236 17334
rect 12196 17052 12248 17058
rect 12196 16994 12248 17000
rect 12104 16372 12156 16378
rect 12104 16314 12156 16320
rect 12116 16106 12144 16314
rect 12104 16100 12156 16106
rect 12104 16042 12156 16048
rect 12208 16038 12236 16994
rect 12196 16032 12248 16038
rect 12196 15974 12248 15980
rect 12012 15012 12064 15018
rect 12012 14954 12064 14960
rect 12196 14808 12248 14814
rect 12196 14750 12248 14756
rect 12104 14468 12156 14474
rect 12104 14410 12156 14416
rect 12012 14400 12064 14406
rect 12012 14342 12064 14348
rect 12024 13726 12052 14342
rect 12116 13930 12144 14410
rect 12208 14241 12236 14750
rect 12194 14232 12250 14241
rect 12194 14167 12250 14176
rect 12104 13924 12156 13930
rect 12104 13866 12156 13872
rect 12012 13720 12064 13726
rect 12012 13662 12064 13668
rect 12196 13108 12248 13114
rect 12196 13050 12248 13056
rect 12208 12842 12236 13050
rect 12196 12836 12248 12842
rect 12196 12778 12248 12784
rect 12300 12230 12328 22774
rect 12748 22492 12800 22498
rect 12748 22434 12800 22440
rect 12760 22022 12788 22434
rect 13128 22090 13156 22842
rect 13496 22430 13524 22910
rect 13484 22424 13536 22430
rect 13484 22366 13536 22372
rect 13116 22084 13168 22090
rect 13116 22026 13168 22032
rect 12748 22016 12800 22022
rect 12748 21958 12800 21964
rect 13496 21954 13524 22366
rect 15416 22288 15468 22294
rect 15416 22230 15468 22236
rect 15428 22022 15456 22230
rect 15416 22016 15468 22022
rect 15416 21958 15468 21964
rect 13484 21948 13536 21954
rect 13484 21890 13536 21896
rect 13300 21404 13352 21410
rect 13300 21346 13352 21352
rect 13312 21002 13340 21346
rect 13300 20996 13352 21002
rect 13300 20938 13352 20944
rect 13312 20662 13340 20938
rect 13300 20656 13352 20662
rect 13300 20598 13352 20604
rect 13496 20322 13524 21890
rect 13576 21200 13628 21206
rect 13576 21142 13628 21148
rect 13588 20798 13616 21142
rect 13576 20792 13628 20798
rect 13576 20734 13628 20740
rect 13588 20390 13616 20734
rect 13760 20724 13812 20730
rect 13760 20666 13812 20672
rect 13576 20384 13628 20390
rect 13576 20326 13628 20332
rect 13484 20316 13536 20322
rect 13484 20258 13536 20264
rect 13496 19914 13524 20258
rect 13668 20180 13720 20186
rect 13668 20122 13720 20128
rect 13484 19908 13536 19914
rect 13484 19850 13536 19856
rect 13680 19574 13708 20122
rect 13668 19568 13720 19574
rect 13668 19510 13720 19516
rect 13574 19264 13630 19273
rect 12932 19228 12984 19234
rect 12932 19170 12984 19176
rect 13484 19228 13536 19234
rect 13574 19199 13630 19208
rect 13484 19170 13536 19176
rect 12748 19160 12800 19166
rect 12748 19102 12800 19108
rect 12760 18622 12788 19102
rect 12748 18616 12800 18622
rect 12748 18558 12800 18564
rect 12944 18486 12972 19170
rect 13116 18616 13168 18622
rect 13116 18558 13168 18564
rect 12932 18480 12984 18486
rect 12932 18422 12984 18428
rect 12944 18010 12972 18422
rect 13128 18146 13156 18558
rect 13496 18554 13524 19170
rect 13588 19166 13616 19199
rect 13576 19160 13628 19166
rect 13576 19102 13628 19108
rect 13588 18826 13616 19102
rect 13576 18820 13628 18826
rect 13576 18762 13628 18768
rect 13484 18548 13536 18554
rect 13484 18490 13536 18496
rect 13116 18140 13168 18146
rect 13116 18082 13168 18088
rect 12932 18004 12984 18010
rect 12932 17946 12984 17952
rect 12378 17768 12434 17777
rect 13128 17738 13156 18082
rect 13668 18072 13720 18078
rect 13668 18014 13720 18020
rect 12378 17703 12434 17712
rect 13116 17732 13168 17738
rect 12392 16990 12420 17703
rect 13116 17674 13168 17680
rect 13680 17670 13708 18014
rect 13668 17664 13720 17670
rect 13668 17606 13720 17612
rect 12380 16984 12432 16990
rect 12380 16926 12432 16932
rect 12392 16650 12420 16926
rect 12380 16644 12432 16650
rect 12380 16586 12432 16592
rect 13116 16440 13168 16446
rect 13116 16382 13168 16388
rect 13128 16038 13156 16382
rect 13116 16032 13168 16038
rect 13116 15974 13168 15980
rect 12656 15216 12708 15222
rect 12656 15158 12708 15164
rect 12668 14950 12696 15158
rect 12656 14944 12708 14950
rect 12656 14886 12708 14892
rect 12932 14740 12984 14746
rect 12932 14682 12984 14688
rect 12944 14474 12972 14682
rect 12932 14468 12984 14474
rect 12932 14410 12984 14416
rect 12840 14196 12892 14202
rect 12840 14138 12892 14144
rect 12852 14105 12880 14138
rect 12838 14096 12894 14105
rect 12838 14031 12894 14040
rect 12288 12224 12340 12230
rect 12288 12166 12340 12172
rect 12852 11736 12880 14031
rect 13128 13114 13156 15974
rect 13392 15896 13444 15902
rect 13392 15838 13444 15844
rect 13668 15896 13720 15902
rect 13668 15838 13720 15844
rect 13404 15358 13432 15838
rect 13576 15828 13628 15834
rect 13576 15770 13628 15776
rect 13588 15494 13616 15770
rect 13576 15488 13628 15494
rect 13576 15430 13628 15436
rect 13392 15352 13444 15358
rect 13392 15294 13444 15300
rect 13404 15222 13432 15294
rect 13392 15216 13444 15222
rect 13392 15158 13444 15164
rect 13300 13584 13352 13590
rect 13300 13526 13352 13532
rect 13312 13182 13340 13526
rect 13404 13250 13432 15158
rect 13588 14950 13616 15430
rect 13680 15018 13708 15838
rect 13668 15012 13720 15018
rect 13668 14954 13720 14960
rect 13576 14944 13628 14950
rect 13576 14886 13628 14892
rect 13588 14474 13616 14886
rect 13576 14468 13628 14474
rect 13576 14410 13628 14416
rect 13588 14270 13616 14410
rect 13576 14264 13628 14270
rect 13576 14206 13628 14212
rect 13392 13244 13444 13250
rect 13392 13186 13444 13192
rect 13300 13176 13352 13182
rect 13300 13118 13352 13124
rect 13116 13108 13168 13114
rect 13116 13050 13168 13056
rect 13404 12842 13432 13186
rect 13392 12836 13444 12842
rect 13392 12778 13444 12784
rect 12852 11708 12972 11736
rect 12840 11612 12892 11618
rect 12840 11554 12892 11560
rect 12852 11074 12880 11554
rect 12944 11482 12972 11708
rect 13300 11680 13352 11686
rect 13300 11622 13352 11628
rect 12932 11476 12984 11482
rect 12932 11418 12984 11424
rect 13312 11414 13340 11622
rect 13024 11408 13076 11414
rect 13024 11350 13076 11356
rect 13208 11408 13260 11414
rect 13208 11350 13260 11356
rect 13300 11408 13352 11414
rect 13300 11350 13352 11356
rect 12840 11068 12892 11074
rect 12840 11010 12892 11016
rect 12564 11000 12616 11006
rect 12564 10942 12616 10948
rect 12288 10864 12340 10870
rect 12288 10806 12340 10812
rect 12300 10530 12328 10806
rect 12288 10524 12340 10530
rect 12288 10466 12340 10472
rect 12300 9986 12328 10466
rect 12288 9980 12340 9986
rect 12288 9922 12340 9928
rect 12012 9912 12064 9918
rect 12012 9854 12064 9860
rect 11840 9328 11960 9356
rect 11840 2914 11868 9328
rect 12024 8422 12052 9854
rect 12576 9578 12604 10942
rect 13036 10870 13064 11350
rect 13220 11006 13248 11350
rect 13312 11006 13340 11350
rect 13484 11136 13536 11142
rect 13484 11078 13536 11084
rect 13208 11000 13260 11006
rect 13208 10942 13260 10948
rect 13300 11000 13352 11006
rect 13300 10942 13352 10948
rect 13024 10864 13076 10870
rect 13024 10806 13076 10812
rect 12748 10524 12800 10530
rect 12748 10466 12800 10472
rect 12760 10122 12788 10466
rect 13116 10388 13168 10394
rect 13116 10330 13168 10336
rect 13128 10122 13156 10330
rect 12748 10116 12800 10122
rect 12748 10058 12800 10064
rect 13116 10116 13168 10122
rect 13116 10058 13168 10064
rect 12564 9572 12616 9578
rect 12564 9514 12616 9520
rect 12472 9436 12524 9442
rect 12472 9378 12524 9384
rect 12484 8966 12512 9378
rect 12576 9034 12604 9514
rect 13312 9442 13340 10942
rect 13392 9912 13444 9918
rect 13392 9854 13444 9860
rect 13404 9782 13432 9854
rect 13392 9776 13444 9782
rect 13392 9718 13444 9724
rect 13300 9436 13352 9442
rect 13300 9378 13352 9384
rect 12564 9028 12616 9034
rect 12564 8970 12616 8976
rect 13404 8966 13432 9718
rect 12472 8960 12524 8966
rect 12472 8902 12524 8908
rect 13392 8960 13444 8966
rect 13392 8902 13444 8908
rect 13116 8824 13168 8830
rect 13116 8766 13168 8772
rect 13024 8756 13076 8762
rect 13024 8698 13076 8704
rect 12012 8416 12064 8422
rect 12012 8358 12064 8364
rect 12024 7946 12052 8358
rect 12932 8144 12984 8150
rect 12932 8086 12984 8092
rect 12012 7940 12064 7946
rect 12012 7882 12064 7888
rect 12944 7810 12972 8086
rect 12932 7804 12984 7810
rect 12932 7746 12984 7752
rect 13036 7742 13064 8698
rect 13128 8218 13156 8766
rect 13404 8490 13432 8902
rect 13392 8484 13444 8490
rect 13392 8426 13444 8432
rect 13116 8212 13168 8218
rect 13116 8154 13168 8160
rect 13024 7736 13076 7742
rect 13024 7678 13076 7684
rect 12564 7668 12616 7674
rect 12564 7610 12616 7616
rect 12576 7334 12604 7610
rect 13036 7402 13064 7678
rect 13024 7396 13076 7402
rect 13024 7338 13076 7344
rect 12564 7328 12616 7334
rect 12564 7270 12616 7276
rect 12576 6858 12604 7270
rect 12840 7260 12892 7266
rect 12840 7202 12892 7208
rect 12748 7192 12800 7198
rect 12748 7134 12800 7140
rect 12564 6852 12616 6858
rect 12564 6794 12616 6800
rect 12760 6518 12788 7134
rect 12852 6654 12880 7202
rect 13128 7062 13156 8154
rect 13392 7940 13444 7946
rect 13392 7882 13444 7888
rect 13404 7742 13432 7882
rect 13496 7810 13524 11078
rect 13484 7804 13536 7810
rect 13484 7746 13536 7752
rect 13392 7736 13444 7742
rect 13392 7678 13444 7684
rect 13116 7056 13168 7062
rect 13116 6998 13168 7004
rect 13128 6858 13156 6998
rect 13116 6852 13168 6858
rect 13116 6794 13168 6800
rect 12840 6648 12892 6654
rect 12840 6590 12892 6596
rect 12748 6512 12800 6518
rect 12748 6454 12800 6460
rect 12840 6308 12892 6314
rect 12840 6250 12892 6256
rect 12288 6240 12340 6246
rect 12288 6182 12340 6188
rect 11920 5152 11972 5158
rect 11920 5094 11972 5100
rect 11932 4546 11960 5094
rect 11920 4540 11972 4546
rect 11920 4482 11972 4488
rect 11828 2908 11880 2914
rect 11828 2850 11880 2856
rect 11840 2506 11868 2850
rect 11828 2500 11880 2506
rect 11828 2442 11880 2448
rect 12196 1956 12248 1962
rect 12196 1898 12248 1904
rect 11828 1616 11880 1622
rect 11828 1558 11880 1564
rect 11840 1350 11868 1558
rect 12208 1418 12236 1898
rect 12300 1826 12328 6182
rect 12380 6036 12432 6042
rect 12380 5978 12432 5984
rect 12392 5566 12420 5978
rect 12852 5566 12880 6250
rect 12380 5560 12432 5566
rect 12380 5502 12432 5508
rect 12748 5560 12800 5566
rect 12748 5502 12800 5508
rect 12840 5560 12892 5566
rect 12840 5502 12892 5508
rect 12392 4478 12420 5502
rect 12760 4682 12788 5502
rect 12852 5158 12880 5502
rect 13668 5424 13720 5430
rect 13668 5366 13720 5372
rect 13680 5226 13708 5366
rect 13668 5220 13720 5226
rect 13668 5162 13720 5168
rect 12840 5152 12892 5158
rect 12840 5094 12892 5100
rect 12748 4676 12800 4682
rect 12748 4618 12800 4624
rect 12852 4614 12880 5094
rect 12840 4608 12892 4614
rect 12840 4550 12892 4556
rect 12380 4472 12432 4478
rect 12380 4414 12432 4420
rect 12380 4336 12432 4342
rect 12380 4278 12432 4284
rect 12392 3390 12420 4278
rect 12380 3384 12432 3390
rect 12380 3326 12432 3332
rect 12472 3316 12524 3322
rect 12472 3258 12524 3264
rect 12484 2370 12512 3258
rect 13208 2908 13260 2914
rect 13208 2850 13260 2856
rect 12472 2364 12524 2370
rect 12472 2306 12524 2312
rect 13220 1962 13248 2850
rect 13300 2840 13352 2846
rect 13300 2782 13352 2788
rect 13312 2302 13340 2782
rect 13772 2438 13800 20666
rect 15428 20390 15456 21958
rect 15888 21886 15916 22910
rect 15980 22838 16008 23522
rect 16164 22974 16192 25630
rect 16256 23654 16284 27315
rect 17716 26368 17768 26374
rect 17716 26310 17768 26316
rect 17728 26238 17756 26310
rect 16520 26232 16572 26238
rect 16520 26174 16572 26180
rect 17716 26232 17768 26238
rect 17716 26174 17768 26180
rect 16532 25286 16560 26174
rect 17900 26096 17952 26102
rect 17900 26038 17952 26044
rect 17624 25688 17676 25694
rect 17624 25630 17676 25636
rect 16796 25552 16848 25558
rect 16796 25494 16848 25500
rect 16808 25354 16836 25494
rect 16796 25348 16848 25354
rect 16796 25290 16848 25296
rect 16520 25280 16572 25286
rect 16520 25222 16572 25228
rect 17636 25218 17664 25630
rect 17716 25620 17768 25626
rect 17716 25562 17768 25568
rect 17624 25212 17676 25218
rect 17624 25154 17676 25160
rect 17348 25144 17400 25150
rect 17348 25086 17400 25092
rect 17360 24470 17388 25086
rect 16428 24464 16480 24470
rect 16428 24406 16480 24412
rect 17348 24464 17400 24470
rect 17348 24406 17400 24412
rect 16440 24130 16468 24406
rect 16428 24124 16480 24130
rect 16428 24066 16480 24072
rect 16244 23648 16296 23654
rect 16244 23590 16296 23596
rect 16440 23586 16468 24066
rect 16520 23920 16572 23926
rect 16520 23862 16572 23868
rect 16888 23920 16940 23926
rect 16888 23862 16940 23868
rect 16428 23580 16480 23586
rect 16428 23522 16480 23528
rect 16152 22968 16204 22974
rect 16152 22910 16204 22916
rect 16428 22900 16480 22906
rect 16428 22842 16480 22848
rect 15968 22832 16020 22838
rect 15968 22774 16020 22780
rect 15980 21954 16008 22774
rect 16336 22492 16388 22498
rect 16336 22434 16388 22440
rect 16348 22090 16376 22434
rect 16440 22430 16468 22842
rect 16428 22424 16480 22430
rect 16428 22366 16480 22372
rect 16336 22084 16388 22090
rect 16336 22026 16388 22032
rect 15968 21948 16020 21954
rect 15968 21890 16020 21896
rect 15876 21880 15928 21886
rect 15876 21822 15928 21828
rect 15888 21546 15916 21822
rect 15968 21744 16020 21750
rect 15968 21686 16020 21692
rect 15876 21540 15928 21546
rect 15876 21482 15928 21488
rect 15416 20384 15468 20390
rect 15416 20326 15468 20332
rect 15428 19914 15456 20326
rect 15416 19908 15468 19914
rect 15416 19850 15468 19856
rect 14128 19568 14180 19574
rect 14128 19510 14180 19516
rect 13852 19024 13904 19030
rect 13852 18966 13904 18972
rect 13864 18622 13892 18966
rect 13852 18616 13904 18622
rect 13852 18558 13904 18564
rect 13864 18214 13892 18558
rect 14140 18554 14168 19510
rect 15784 18752 15836 18758
rect 15784 18694 15836 18700
rect 15508 18616 15560 18622
rect 15508 18558 15560 18564
rect 14128 18548 14180 18554
rect 14128 18490 14180 18496
rect 13852 18208 13904 18214
rect 13852 18150 13904 18156
rect 13864 17738 13892 18150
rect 14140 17942 14168 18490
rect 14128 17936 14180 17942
rect 14128 17878 14180 17884
rect 13852 17732 13904 17738
rect 13852 17674 13904 17680
rect 13864 17466 13892 17674
rect 14140 17534 14168 17878
rect 15138 17632 15194 17641
rect 15138 17567 15194 17576
rect 14128 17528 14180 17534
rect 14128 17470 14180 17476
rect 13852 17460 13904 17466
rect 13852 17402 13904 17408
rect 14140 15426 14168 17470
rect 14588 17460 14640 17466
rect 14588 17402 14640 17408
rect 14600 17194 14628 17402
rect 14588 17188 14640 17194
rect 14588 17130 14640 17136
rect 14600 16650 14628 17130
rect 15152 17058 15180 17567
rect 15140 17052 15192 17058
rect 15140 16994 15192 17000
rect 14680 16848 14732 16854
rect 14680 16790 14732 16796
rect 14692 16650 14720 16790
rect 15152 16650 15180 16994
rect 15416 16848 15468 16854
rect 15416 16790 15468 16796
rect 14588 16644 14640 16650
rect 14588 16586 14640 16592
rect 14680 16644 14732 16650
rect 14680 16586 14732 16592
rect 15140 16644 15192 16650
rect 15140 16586 15192 16592
rect 14692 15902 14720 16586
rect 15152 16446 15180 16586
rect 15428 16514 15456 16790
rect 15416 16508 15468 16514
rect 15416 16450 15468 16456
rect 15140 16440 15192 16446
rect 15140 16382 15192 16388
rect 15324 16372 15376 16378
rect 15324 16314 15376 16320
rect 14680 15896 14732 15902
rect 14680 15838 14732 15844
rect 15232 15896 15284 15902
rect 15232 15838 15284 15844
rect 15244 15562 15272 15838
rect 15336 15766 15364 16314
rect 15324 15760 15376 15766
rect 15324 15702 15376 15708
rect 15232 15556 15284 15562
rect 15232 15498 15284 15504
rect 15336 15426 15364 15702
rect 15428 15562 15456 16450
rect 15416 15556 15468 15562
rect 15416 15498 15468 15504
rect 14128 15420 14180 15426
rect 14128 15362 14180 15368
rect 15324 15420 15376 15426
rect 15324 15362 15376 15368
rect 14036 14128 14088 14134
rect 14036 14070 14088 14076
rect 13944 13720 13996 13726
rect 13944 13662 13996 13668
rect 13956 11414 13984 13662
rect 13944 11408 13996 11414
rect 13944 11350 13996 11356
rect 13956 11210 13984 11350
rect 13944 11204 13996 11210
rect 13944 11146 13996 11152
rect 13852 10524 13904 10530
rect 13852 10466 13904 10472
rect 13864 10122 13892 10466
rect 13852 10116 13904 10122
rect 13852 10058 13904 10064
rect 13864 9374 13892 10058
rect 13852 9368 13904 9374
rect 13852 9310 13904 9316
rect 14048 2914 14076 14070
rect 15520 12706 15548 18558
rect 15796 18214 15824 18694
rect 15876 18548 15928 18554
rect 15876 18490 15928 18496
rect 15784 18208 15836 18214
rect 15784 18150 15836 18156
rect 15796 17602 15824 18150
rect 15888 17738 15916 18490
rect 15980 17942 16008 21686
rect 16348 19098 16376 22026
rect 16440 22022 16468 22366
rect 16532 22362 16560 23862
rect 16704 23376 16756 23382
rect 16704 23318 16756 23324
rect 16716 23178 16744 23318
rect 16704 23172 16756 23178
rect 16704 23114 16756 23120
rect 16716 22430 16744 23114
rect 16900 22498 16928 23862
rect 16888 22492 16940 22498
rect 16888 22434 16940 22440
rect 16704 22424 16756 22430
rect 16704 22366 16756 22372
rect 16520 22356 16572 22362
rect 16520 22298 16572 22304
rect 16532 22090 16560 22298
rect 16520 22084 16572 22090
rect 16520 22026 16572 22032
rect 16428 22016 16480 22022
rect 16428 21958 16480 21964
rect 16440 21410 16468 21958
rect 16716 21886 16744 22366
rect 16704 21880 16756 21886
rect 16704 21822 16756 21828
rect 16716 21410 16744 21822
rect 16900 21546 16928 22434
rect 17164 21812 17216 21818
rect 17164 21754 17216 21760
rect 16888 21540 16940 21546
rect 16888 21482 16940 21488
rect 17176 21410 17204 21754
rect 17360 21750 17388 24406
rect 17728 22566 17756 25562
rect 17912 24470 17940 26038
rect 17992 25212 18044 25218
rect 17992 25154 18044 25160
rect 18004 24606 18032 25154
rect 17992 24600 18044 24606
rect 17992 24542 18044 24548
rect 17900 24464 17952 24470
rect 17900 24406 17952 24412
rect 18004 23926 18032 24542
rect 17992 23920 18044 23926
rect 17992 23862 18044 23868
rect 18084 23580 18136 23586
rect 18084 23522 18136 23528
rect 18096 22974 18124 23522
rect 18084 22968 18136 22974
rect 18084 22910 18136 22916
rect 17716 22560 17768 22566
rect 17716 22502 17768 22508
rect 17348 21744 17400 21750
rect 17348 21686 17400 21692
rect 16428 21404 16480 21410
rect 16428 21346 16480 21352
rect 16704 21404 16756 21410
rect 16704 21346 16756 21352
rect 17164 21404 17216 21410
rect 17164 21346 17216 21352
rect 16440 21002 16468 21346
rect 16428 20996 16480 21002
rect 16428 20938 16480 20944
rect 16716 20866 16744 21346
rect 16796 21336 16848 21342
rect 16796 21278 16848 21284
rect 16704 20860 16756 20866
rect 16704 20802 16756 20808
rect 16808 20662 16836 21278
rect 16980 21268 17032 21274
rect 16980 21210 17032 21216
rect 16992 20934 17020 21210
rect 17176 21002 17204 21346
rect 18280 21206 18308 27315
rect 18864 27084 19184 27104
rect 18864 27082 18876 27084
rect 18932 27082 18956 27084
rect 19012 27082 19036 27084
rect 19092 27082 19116 27084
rect 19172 27082 19184 27084
rect 18864 27030 18870 27082
rect 18932 27030 18934 27082
rect 19114 27030 19116 27082
rect 19178 27030 19184 27082
rect 18864 27028 18876 27030
rect 18932 27028 18956 27030
rect 19012 27028 19036 27030
rect 19092 27028 19116 27030
rect 19172 27028 19184 27030
rect 18864 27008 19184 27028
rect 19280 26300 19332 26306
rect 19280 26242 19332 26248
rect 18360 26096 18412 26102
rect 18360 26038 18412 26044
rect 18372 25762 18400 26038
rect 18864 25996 19184 26016
rect 18864 25994 18876 25996
rect 18932 25994 18956 25996
rect 19012 25994 19036 25996
rect 19092 25994 19116 25996
rect 19172 25994 19184 25996
rect 18864 25942 18870 25994
rect 18932 25942 18934 25994
rect 19114 25942 19116 25994
rect 19178 25942 19184 25994
rect 18864 25940 18876 25942
rect 18932 25940 18956 25942
rect 19012 25940 19036 25942
rect 19092 25940 19116 25942
rect 19172 25940 19184 25942
rect 18864 25920 19184 25940
rect 18360 25756 18412 25762
rect 18360 25698 18412 25704
rect 18372 25082 18400 25698
rect 19004 25688 19056 25694
rect 19004 25630 19056 25636
rect 19016 25558 19044 25630
rect 19004 25552 19056 25558
rect 19004 25494 19056 25500
rect 19016 25082 19044 25494
rect 18360 25076 18412 25082
rect 18360 25018 18412 25024
rect 19004 25076 19056 25082
rect 19004 25018 19056 25024
rect 18864 24908 19184 24928
rect 18864 24906 18876 24908
rect 18932 24906 18956 24908
rect 19012 24906 19036 24908
rect 19092 24906 19116 24908
rect 19172 24906 19184 24908
rect 18864 24854 18870 24906
rect 18932 24854 18934 24906
rect 19114 24854 19116 24906
rect 19178 24854 19184 24906
rect 18864 24852 18876 24854
rect 18932 24852 18956 24854
rect 19012 24852 19036 24854
rect 19092 24852 19116 24854
rect 19172 24852 19184 24854
rect 18864 24832 19184 24852
rect 18452 24668 18504 24674
rect 18452 24610 18504 24616
rect 18820 24668 18872 24674
rect 18820 24610 18872 24616
rect 18464 24266 18492 24610
rect 18728 24600 18780 24606
rect 18728 24542 18780 24548
rect 18544 24464 18596 24470
rect 18544 24406 18596 24412
rect 18556 24266 18584 24406
rect 18452 24260 18504 24266
rect 18452 24202 18504 24208
rect 18544 24260 18596 24266
rect 18544 24202 18596 24208
rect 18464 23874 18492 24202
rect 18740 24198 18768 24542
rect 18728 24192 18780 24198
rect 18728 24134 18780 24140
rect 18372 23846 18492 23874
rect 18372 23722 18400 23846
rect 18360 23716 18412 23722
rect 18360 23658 18412 23664
rect 18372 23178 18400 23658
rect 18636 23580 18688 23586
rect 18636 23522 18688 23528
rect 18360 23172 18412 23178
rect 18360 23114 18412 23120
rect 18648 22974 18676 23522
rect 18740 23178 18768 24134
rect 18832 24130 18860 24610
rect 18820 24124 18872 24130
rect 18820 24066 18872 24072
rect 18864 23820 19184 23840
rect 18864 23818 18876 23820
rect 18932 23818 18956 23820
rect 19012 23818 19036 23820
rect 19092 23818 19116 23820
rect 19172 23818 19184 23820
rect 18864 23766 18870 23818
rect 18932 23766 18934 23818
rect 19114 23766 19116 23818
rect 19178 23766 19184 23818
rect 18864 23764 18876 23766
rect 18932 23764 18956 23766
rect 19012 23764 19036 23766
rect 19092 23764 19116 23766
rect 19172 23764 19184 23766
rect 18864 23744 19184 23764
rect 18728 23172 18780 23178
rect 18728 23114 18780 23120
rect 18544 22968 18596 22974
rect 18544 22910 18596 22916
rect 18636 22968 18688 22974
rect 18636 22910 18688 22916
rect 18556 22634 18584 22910
rect 18864 22732 19184 22752
rect 18864 22730 18876 22732
rect 18932 22730 18956 22732
rect 19012 22730 19036 22732
rect 19092 22730 19116 22732
rect 19172 22730 19184 22732
rect 18864 22678 18870 22730
rect 18932 22678 18934 22730
rect 19114 22678 19116 22730
rect 19178 22678 19184 22730
rect 18864 22676 18876 22678
rect 18932 22676 18956 22678
rect 19012 22676 19036 22678
rect 19092 22676 19116 22678
rect 19172 22676 19184 22678
rect 18864 22656 19184 22676
rect 18544 22628 18596 22634
rect 18544 22570 18596 22576
rect 19096 22288 19148 22294
rect 19096 22230 19148 22236
rect 19108 22090 19136 22230
rect 19096 22084 19148 22090
rect 19096 22026 19148 22032
rect 19108 21886 19136 22026
rect 19096 21880 19148 21886
rect 19096 21822 19148 21828
rect 18864 21644 19184 21664
rect 18864 21642 18876 21644
rect 18932 21642 18956 21644
rect 19012 21642 19036 21644
rect 19092 21642 19116 21644
rect 19172 21642 19184 21644
rect 18864 21590 18870 21642
rect 18932 21590 18934 21642
rect 19114 21590 19116 21642
rect 19178 21590 19184 21642
rect 18864 21588 18876 21590
rect 18932 21588 18956 21590
rect 19012 21588 19036 21590
rect 19092 21588 19116 21590
rect 19172 21588 19184 21590
rect 18864 21568 19184 21588
rect 18268 21200 18320 21206
rect 18268 21142 18320 21148
rect 17164 20996 17216 21002
rect 17164 20938 17216 20944
rect 16980 20928 17032 20934
rect 16980 20870 17032 20876
rect 16796 20656 16848 20662
rect 16796 20598 16848 20604
rect 16428 20384 16480 20390
rect 16428 20326 16480 20332
rect 16440 19914 16468 20326
rect 16808 20322 16836 20598
rect 16796 20316 16848 20322
rect 16796 20258 16848 20264
rect 16428 19908 16480 19914
rect 16428 19850 16480 19856
rect 16336 19092 16388 19098
rect 16336 19034 16388 19040
rect 16244 18548 16296 18554
rect 16244 18490 16296 18496
rect 16256 18214 16284 18490
rect 16244 18208 16296 18214
rect 16244 18150 16296 18156
rect 15968 17936 16020 17942
rect 15968 17878 16020 17884
rect 15876 17732 15928 17738
rect 15876 17674 15928 17680
rect 15784 17596 15836 17602
rect 15784 17538 15836 17544
rect 15980 17398 16008 17878
rect 15968 17392 16020 17398
rect 15968 17334 16020 17340
rect 15876 15556 15928 15562
rect 15876 15498 15928 15504
rect 15784 15488 15836 15494
rect 15784 15430 15836 15436
rect 15796 15290 15824 15430
rect 15784 15284 15836 15290
rect 15784 15226 15836 15232
rect 15888 15018 15916 15498
rect 15876 15012 15928 15018
rect 15876 14954 15928 14960
rect 15980 14214 16008 17334
rect 16440 17058 16468 19850
rect 16808 19846 16836 20258
rect 16992 19846 17020 20870
rect 18360 20656 18412 20662
rect 18360 20598 18412 20604
rect 17992 20316 18044 20322
rect 17992 20258 18044 20264
rect 16796 19840 16848 19846
rect 16796 19782 16848 19788
rect 16980 19840 17032 19846
rect 16980 19782 17032 19788
rect 17900 19092 17952 19098
rect 17900 19034 17952 19040
rect 17912 18622 17940 19034
rect 18004 19030 18032 20258
rect 18084 19772 18136 19778
rect 18084 19714 18136 19720
rect 17992 19024 18044 19030
rect 17992 18966 18044 18972
rect 18004 18758 18032 18966
rect 17992 18752 18044 18758
rect 17992 18694 18044 18700
rect 18096 18622 18124 19714
rect 18176 19568 18228 19574
rect 18176 19510 18228 19516
rect 18188 19166 18216 19510
rect 18176 19160 18228 19166
rect 18176 19102 18228 19108
rect 18188 18826 18216 19102
rect 18176 18820 18228 18826
rect 18176 18762 18228 18768
rect 17900 18616 17952 18622
rect 17900 18558 17952 18564
rect 18084 18616 18136 18622
rect 18084 18558 18136 18564
rect 16428 17052 16480 17058
rect 16428 16994 16480 17000
rect 16440 16514 16468 16994
rect 16704 16984 16756 16990
rect 16704 16926 16756 16932
rect 16428 16508 16480 16514
rect 16428 16450 16480 16456
rect 16440 16106 16468 16450
rect 16716 16310 16744 16926
rect 17808 16848 17860 16854
rect 17808 16790 17860 16796
rect 17820 16582 17848 16790
rect 17808 16576 17860 16582
rect 17808 16518 17860 16524
rect 17164 16440 17216 16446
rect 17164 16382 17216 16388
rect 16704 16304 16756 16310
rect 16704 16246 16756 16252
rect 16428 16100 16480 16106
rect 16428 16042 16480 16048
rect 16440 14882 16468 16042
rect 16612 15964 16664 15970
rect 16612 15906 16664 15912
rect 16624 15426 16652 15906
rect 16716 15902 16744 16246
rect 16980 15964 17032 15970
rect 16980 15906 17032 15912
rect 17072 15964 17124 15970
rect 17072 15906 17124 15912
rect 16704 15896 16756 15902
rect 16704 15838 16756 15844
rect 16888 15760 16940 15766
rect 16888 15702 16940 15708
rect 16900 15562 16928 15702
rect 16888 15556 16940 15562
rect 16888 15498 16940 15504
rect 16612 15420 16664 15426
rect 16612 15362 16664 15368
rect 16428 14876 16480 14882
rect 16428 14818 16480 14824
rect 16152 14808 16204 14814
rect 16152 14750 16204 14756
rect 16164 14474 16192 14750
rect 16152 14468 16204 14474
rect 16152 14410 16204 14416
rect 16440 14406 16468 14818
rect 16624 14814 16652 15362
rect 16900 14950 16928 15498
rect 16992 15358 17020 15906
rect 17084 15494 17112 15906
rect 17072 15488 17124 15494
rect 17072 15430 17124 15436
rect 16980 15352 17032 15358
rect 16980 15294 17032 15300
rect 16888 14944 16940 14950
rect 16888 14886 16940 14892
rect 17176 14882 17204 16382
rect 17820 15970 17848 16518
rect 17912 16106 17940 18558
rect 18096 18078 18124 18558
rect 18188 18282 18216 18762
rect 18372 18622 18400 20598
rect 18864 20556 19184 20576
rect 18864 20554 18876 20556
rect 18932 20554 18956 20556
rect 19012 20554 19036 20556
rect 19092 20554 19116 20556
rect 19172 20554 19184 20556
rect 18864 20502 18870 20554
rect 18932 20502 18934 20554
rect 19114 20502 19116 20554
rect 19178 20502 19184 20554
rect 18864 20500 18876 20502
rect 18932 20500 18956 20502
rect 19012 20500 19036 20502
rect 19092 20500 19116 20502
rect 19172 20500 19184 20502
rect 18864 20480 19184 20500
rect 18728 19704 18780 19710
rect 18728 19646 18780 19652
rect 18740 19234 18768 19646
rect 18864 19468 19184 19488
rect 18864 19466 18876 19468
rect 18932 19466 18956 19468
rect 19012 19466 19036 19468
rect 19092 19466 19116 19468
rect 19172 19466 19184 19468
rect 18864 19414 18870 19466
rect 18932 19414 18934 19466
rect 19114 19414 19116 19466
rect 19178 19414 19184 19466
rect 18864 19412 18876 19414
rect 18932 19412 18956 19414
rect 19012 19412 19036 19414
rect 19092 19412 19116 19414
rect 19172 19412 19184 19414
rect 18864 19392 19184 19412
rect 18544 19228 18596 19234
rect 18544 19170 18596 19176
rect 18728 19228 18780 19234
rect 18728 19170 18780 19176
rect 18360 18616 18412 18622
rect 18360 18558 18412 18564
rect 18556 18486 18584 19170
rect 18740 18690 18768 19170
rect 19292 19098 19320 26242
rect 19648 25756 19700 25762
rect 19648 25698 19700 25704
rect 19464 25620 19516 25626
rect 19464 25562 19516 25568
rect 19476 25354 19504 25562
rect 19464 25348 19516 25354
rect 19464 25290 19516 25296
rect 19660 25014 19688 25698
rect 19648 25008 19700 25014
rect 19648 24950 19700 24956
rect 19660 24674 19688 24950
rect 19648 24668 19700 24674
rect 19648 24610 19700 24616
rect 20200 22492 20252 22498
rect 20200 22434 20252 22440
rect 19372 21812 19424 21818
rect 19372 21754 19424 21760
rect 19384 21002 19412 21754
rect 20108 21744 20160 21750
rect 20108 21686 20160 21692
rect 20120 21206 20148 21686
rect 20212 21478 20240 22434
rect 20200 21472 20252 21478
rect 20200 21414 20252 21420
rect 20108 21200 20160 21206
rect 20108 21142 20160 21148
rect 19372 20996 19424 21002
rect 19372 20938 19424 20944
rect 20120 20322 20148 21142
rect 20304 20730 20332 27315
rect 20476 26164 20528 26170
rect 20476 26106 20528 26112
rect 21856 26164 21908 26170
rect 21856 26106 21908 26112
rect 20488 25558 20516 26106
rect 20568 26096 20620 26102
rect 20568 26038 20620 26044
rect 20476 25552 20528 25558
rect 20476 25494 20528 25500
rect 20488 25150 20516 25494
rect 20476 25144 20528 25150
rect 20476 25086 20528 25092
rect 20488 24198 20516 25086
rect 20580 25082 20608 26038
rect 21868 25830 21896 26106
rect 21856 25824 21908 25830
rect 21856 25766 21908 25772
rect 20844 25688 20896 25694
rect 20844 25630 20896 25636
rect 21120 25688 21172 25694
rect 21120 25630 21172 25636
rect 20660 25620 20712 25626
rect 20660 25562 20712 25568
rect 20672 25150 20700 25562
rect 20660 25144 20712 25150
rect 20660 25086 20712 25092
rect 20568 25076 20620 25082
rect 20568 25018 20620 25024
rect 20580 24606 20608 25018
rect 20856 24810 20884 25630
rect 21132 25286 21160 25630
rect 21868 25336 21896 25766
rect 21948 25348 22000 25354
rect 21868 25308 21948 25336
rect 21948 25290 22000 25296
rect 21120 25280 21172 25286
rect 21120 25222 21172 25228
rect 20844 24804 20896 24810
rect 20844 24746 20896 24752
rect 21488 24668 21540 24674
rect 21488 24610 21540 24616
rect 20568 24600 20620 24606
rect 20568 24542 20620 24548
rect 20476 24192 20528 24198
rect 20476 24134 20528 24140
rect 20488 23994 20516 24134
rect 20476 23988 20528 23994
rect 20476 23930 20528 23936
rect 20580 23586 20608 24542
rect 20752 24532 20804 24538
rect 20752 24474 20804 24480
rect 20660 24464 20712 24470
rect 20660 24406 20712 24412
rect 20672 24198 20700 24406
rect 20660 24192 20712 24198
rect 20660 24134 20712 24140
rect 20672 23874 20700 24134
rect 20764 24130 20792 24474
rect 21028 24464 21080 24470
rect 21028 24406 21080 24412
rect 21396 24464 21448 24470
rect 21396 24406 21448 24412
rect 20752 24124 20804 24130
rect 20752 24066 20804 24072
rect 21040 24062 21068 24406
rect 21028 24056 21080 24062
rect 21028 23998 21080 24004
rect 21408 23926 21436 24406
rect 21500 24266 21528 24610
rect 21488 24260 21540 24266
rect 21488 24202 21540 24208
rect 21396 23920 21448 23926
rect 20672 23846 20792 23874
rect 21396 23862 21448 23868
rect 20568 23580 20620 23586
rect 20568 23522 20620 23528
rect 20660 23580 20712 23586
rect 20660 23522 20712 23528
rect 20672 23178 20700 23522
rect 20660 23172 20712 23178
rect 20660 23114 20712 23120
rect 20476 22424 20528 22430
rect 20476 22366 20528 22372
rect 20488 21886 20516 22366
rect 20476 21880 20528 21886
rect 20476 21822 20528 21828
rect 20488 21546 20516 21822
rect 20476 21540 20528 21546
rect 20476 21482 20528 21488
rect 20764 21290 20792 23846
rect 20936 23512 20988 23518
rect 20936 23454 20988 23460
rect 20844 23376 20896 23382
rect 20844 23318 20896 23324
rect 20856 22838 20884 23318
rect 20948 23178 20976 23454
rect 20936 23172 20988 23178
rect 20936 23114 20988 23120
rect 20844 22832 20896 22838
rect 20844 22774 20896 22780
rect 20856 22498 20884 22774
rect 20844 22492 20896 22498
rect 20844 22434 20896 22440
rect 21408 21460 21436 23862
rect 21500 23722 21528 24202
rect 21488 23716 21540 23722
rect 21488 23658 21540 23664
rect 21672 22900 21724 22906
rect 21672 22842 21724 22848
rect 21408 21432 21528 21460
rect 21304 21404 21356 21410
rect 21356 21364 21436 21392
rect 21304 21346 21356 21352
rect 21212 21336 21264 21342
rect 20764 21262 20884 21290
rect 21212 21278 21264 21284
rect 20752 21200 20804 21206
rect 20752 21142 20804 21148
rect 20764 20798 20792 21142
rect 20752 20792 20804 20798
rect 20752 20734 20804 20740
rect 20292 20724 20344 20730
rect 20292 20666 20344 20672
rect 20108 20316 20160 20322
rect 20108 20258 20160 20264
rect 19372 19636 19424 19642
rect 19372 19578 19424 19584
rect 19384 19234 19412 19578
rect 20120 19370 20148 20258
rect 20856 19914 20884 21262
rect 21224 20662 21252 21278
rect 21408 20662 21436 21364
rect 21212 20656 21264 20662
rect 21212 20598 21264 20604
rect 21396 20656 21448 20662
rect 21396 20598 21448 20604
rect 20936 20112 20988 20118
rect 20936 20054 20988 20060
rect 20660 19908 20712 19914
rect 20660 19850 20712 19856
rect 20844 19908 20896 19914
rect 20844 19850 20896 19856
rect 20476 19772 20528 19778
rect 20476 19714 20528 19720
rect 20292 19704 20344 19710
rect 20292 19646 20344 19652
rect 20108 19364 20160 19370
rect 20108 19306 20160 19312
rect 19372 19228 19424 19234
rect 19372 19170 19424 19176
rect 19280 19092 19332 19098
rect 19280 19034 19332 19040
rect 19924 19092 19976 19098
rect 19924 19034 19976 19040
rect 19280 18752 19332 18758
rect 19280 18694 19332 18700
rect 18728 18684 18780 18690
rect 18728 18626 18780 18632
rect 18544 18480 18596 18486
rect 18544 18422 18596 18428
rect 18176 18276 18228 18282
rect 18176 18218 18228 18224
rect 18084 18072 18136 18078
rect 18084 18014 18136 18020
rect 18556 16446 18584 18422
rect 18740 18214 18768 18626
rect 18864 18380 19184 18400
rect 18864 18378 18876 18380
rect 18932 18378 18956 18380
rect 19012 18378 19036 18380
rect 19092 18378 19116 18380
rect 19172 18378 19184 18380
rect 18864 18326 18870 18378
rect 18932 18326 18934 18378
rect 19114 18326 19116 18378
rect 19178 18326 19184 18378
rect 18864 18324 18876 18326
rect 18932 18324 18956 18326
rect 19012 18324 19036 18326
rect 19092 18324 19116 18326
rect 19172 18324 19184 18326
rect 18864 18304 19184 18324
rect 18728 18208 18780 18214
rect 18728 18150 18780 18156
rect 18636 18140 18688 18146
rect 18636 18082 18688 18088
rect 18648 17670 18676 18082
rect 18740 17738 18768 18150
rect 18728 17732 18780 17738
rect 18728 17674 18780 17680
rect 18636 17664 18688 17670
rect 18636 17606 18688 17612
rect 18864 17292 19184 17312
rect 18864 17290 18876 17292
rect 18932 17290 18956 17292
rect 19012 17290 19036 17292
rect 19092 17290 19116 17292
rect 19172 17290 19184 17292
rect 18864 17238 18870 17290
rect 18932 17238 18934 17290
rect 19114 17238 19116 17290
rect 19178 17238 19184 17290
rect 18864 17236 18876 17238
rect 18932 17236 18956 17238
rect 19012 17236 19036 17238
rect 19092 17236 19116 17238
rect 19172 17236 19184 17238
rect 18864 17216 19184 17236
rect 19292 16446 19320 18694
rect 18544 16440 18596 16446
rect 18544 16382 18596 16388
rect 19280 16440 19332 16446
rect 19280 16382 19332 16388
rect 19372 16304 19424 16310
rect 19372 16246 19424 16252
rect 18864 16204 19184 16224
rect 18864 16202 18876 16204
rect 18932 16202 18956 16204
rect 19012 16202 19036 16204
rect 19092 16202 19116 16204
rect 19172 16202 19184 16204
rect 18864 16150 18870 16202
rect 18932 16150 18934 16202
rect 19114 16150 19116 16202
rect 19178 16150 19184 16202
rect 18864 16148 18876 16150
rect 18932 16148 18956 16150
rect 19012 16148 19036 16150
rect 19092 16148 19116 16150
rect 19172 16148 19184 16150
rect 18864 16128 19184 16148
rect 17900 16100 17952 16106
rect 17900 16042 17952 16048
rect 17808 15964 17860 15970
rect 17808 15906 17860 15912
rect 18864 15116 19184 15136
rect 18864 15114 18876 15116
rect 18932 15114 18956 15116
rect 19012 15114 19036 15116
rect 19092 15114 19116 15116
rect 19172 15114 19184 15116
rect 18864 15062 18870 15114
rect 18932 15062 18934 15114
rect 19114 15062 19116 15114
rect 19178 15062 19184 15114
rect 18864 15060 18876 15062
rect 18932 15060 18956 15062
rect 19012 15060 19036 15062
rect 19092 15060 19116 15062
rect 19172 15060 19184 15062
rect 18864 15040 19184 15060
rect 17164 14876 17216 14882
rect 17164 14818 17216 14824
rect 17992 14876 18044 14882
rect 17992 14818 18044 14824
rect 16612 14808 16664 14814
rect 16612 14750 16664 14756
rect 16624 14406 16652 14750
rect 16428 14400 16480 14406
rect 16428 14342 16480 14348
rect 16612 14400 16664 14406
rect 16612 14342 16664 14348
rect 15888 14186 16008 14214
rect 17176 14202 17204 14818
rect 17440 14672 17492 14678
rect 17440 14614 17492 14620
rect 17452 14474 17480 14614
rect 17440 14468 17492 14474
rect 17440 14410 17492 14416
rect 17164 14196 17216 14202
rect 15784 13652 15836 13658
rect 15784 13594 15836 13600
rect 15796 13386 15824 13594
rect 15784 13380 15836 13386
rect 15784 13322 15836 13328
rect 15508 12700 15560 12706
rect 15508 12642 15560 12648
rect 15416 12632 15468 12638
rect 15416 12574 15468 12580
rect 14312 12496 14364 12502
rect 14312 12438 14364 12444
rect 14324 12162 14352 12438
rect 14312 12156 14364 12162
rect 14312 12098 14364 12104
rect 14496 12020 14548 12026
rect 14496 11962 14548 11968
rect 15324 12020 15376 12026
rect 15428 12008 15456 12574
rect 15376 11980 15456 12008
rect 15324 11962 15376 11968
rect 14128 11204 14180 11210
rect 14128 11146 14180 11152
rect 14220 11204 14272 11210
rect 14220 11146 14272 11152
rect 14140 9442 14168 11146
rect 14232 10938 14260 11146
rect 14220 10932 14272 10938
rect 14220 10874 14272 10880
rect 14220 10592 14272 10598
rect 14220 10534 14272 10540
rect 14232 9850 14260 10534
rect 14404 10320 14456 10326
rect 14404 10262 14456 10268
rect 14312 10048 14364 10054
rect 14312 9990 14364 9996
rect 14324 9850 14352 9990
rect 14220 9844 14272 9850
rect 14220 9786 14272 9792
rect 14312 9844 14364 9850
rect 14312 9786 14364 9792
rect 14128 9436 14180 9442
rect 14128 9378 14180 9384
rect 14232 8966 14260 9786
rect 14416 9510 14444 10262
rect 14508 10122 14536 11962
rect 15428 11754 15456 11980
rect 15416 11748 15468 11754
rect 15416 11690 15468 11696
rect 15520 11618 15548 12642
rect 15600 11680 15652 11686
rect 15600 11622 15652 11628
rect 15508 11612 15560 11618
rect 15508 11554 15560 11560
rect 14864 11476 14916 11482
rect 14864 11418 14916 11424
rect 14772 11408 14824 11414
rect 14772 11350 14824 11356
rect 14784 11142 14812 11350
rect 14772 11136 14824 11142
rect 14772 11078 14824 11084
rect 14784 10666 14812 11078
rect 14876 11074 14904 11418
rect 15520 11074 15548 11554
rect 14864 11068 14916 11074
rect 15508 11068 15560 11074
rect 14916 11028 14996 11056
rect 14864 11010 14916 11016
rect 14772 10660 14824 10666
rect 14772 10602 14824 10608
rect 14496 10116 14548 10122
rect 14496 10058 14548 10064
rect 14404 9504 14456 9510
rect 14404 9446 14456 9452
rect 14772 9436 14824 9442
rect 14772 9378 14824 9384
rect 14220 8960 14272 8966
rect 14220 8902 14272 8908
rect 14680 8824 14732 8830
rect 14680 8766 14732 8772
rect 14496 8756 14548 8762
rect 14496 8698 14548 8704
rect 14220 7260 14272 7266
rect 14220 7202 14272 7208
rect 14232 6518 14260 7202
rect 14508 6858 14536 8698
rect 14692 8286 14720 8766
rect 14784 8490 14812 9378
rect 14864 9232 14916 9238
rect 14864 9174 14916 9180
rect 14876 9034 14904 9174
rect 14864 9028 14916 9034
rect 14864 8970 14916 8976
rect 14772 8484 14824 8490
rect 14772 8426 14824 8432
rect 14680 8280 14732 8286
rect 14680 8222 14732 8228
rect 14772 8280 14824 8286
rect 14772 8222 14824 8228
rect 14784 7674 14812 8222
rect 14772 7668 14824 7674
rect 14772 7610 14824 7616
rect 14496 6852 14548 6858
rect 14496 6794 14548 6800
rect 14220 6512 14272 6518
rect 14220 6454 14272 6460
rect 14232 6246 14260 6454
rect 14220 6240 14272 6246
rect 14220 6182 14272 6188
rect 14588 6240 14640 6246
rect 14588 6182 14640 6188
rect 14220 5696 14272 5702
rect 14220 5638 14272 5644
rect 14232 5566 14260 5638
rect 14220 5560 14272 5566
rect 14220 5502 14272 5508
rect 14496 5492 14548 5498
rect 14496 5434 14548 5440
rect 14508 4070 14536 5434
rect 14600 5226 14628 6182
rect 14784 6178 14812 7610
rect 14864 7600 14916 7606
rect 14864 7542 14916 7548
rect 14876 6586 14904 7542
rect 14864 6580 14916 6586
rect 14864 6522 14916 6528
rect 14772 6172 14824 6178
rect 14772 6114 14824 6120
rect 14784 5702 14812 6114
rect 14772 5696 14824 5702
rect 14772 5638 14824 5644
rect 14968 5566 14996 11028
rect 15508 11010 15560 11016
rect 15612 10530 15640 11622
rect 15600 10524 15652 10530
rect 15600 10466 15652 10472
rect 15324 10456 15376 10462
rect 15324 10398 15376 10404
rect 15140 10320 15192 10326
rect 15140 10262 15192 10268
rect 15152 9918 15180 10262
rect 15140 9912 15192 9918
rect 15140 9854 15192 9860
rect 15336 9578 15364 10398
rect 15600 9912 15652 9918
rect 15600 9854 15652 9860
rect 15692 9912 15744 9918
rect 15692 9854 15744 9860
rect 15324 9572 15376 9578
rect 15324 9514 15376 9520
rect 15612 9510 15640 9854
rect 15704 9782 15732 9854
rect 15796 9782 15824 13322
rect 15888 12502 15916 14186
rect 17164 14138 17216 14144
rect 17808 14196 17860 14202
rect 17808 14138 17860 14144
rect 15968 13720 16020 13726
rect 15968 13662 16020 13668
rect 15980 13386 16008 13662
rect 17820 13386 17848 14138
rect 18004 13930 18032 14818
rect 18728 14672 18780 14678
rect 18728 14614 18780 14620
rect 18452 14332 18504 14338
rect 18452 14274 18504 14280
rect 18464 14134 18492 14274
rect 18740 14270 18768 14614
rect 18728 14264 18780 14270
rect 18728 14206 18780 14212
rect 19280 14264 19332 14270
rect 19280 14206 19332 14212
rect 18452 14128 18504 14134
rect 18452 14070 18504 14076
rect 17992 13924 18044 13930
rect 17992 13866 18044 13872
rect 18464 13726 18492 14070
rect 18864 14028 19184 14048
rect 18864 14026 18876 14028
rect 18932 14026 18956 14028
rect 19012 14026 19036 14028
rect 19092 14026 19116 14028
rect 19172 14026 19184 14028
rect 18864 13974 18870 14026
rect 18932 13974 18934 14026
rect 19114 13974 19116 14026
rect 19178 13974 19184 14026
rect 18864 13972 18876 13974
rect 18932 13972 18956 13974
rect 19012 13972 19036 13974
rect 19092 13972 19116 13974
rect 19172 13972 19184 13974
rect 18864 13952 19184 13972
rect 18544 13924 18596 13930
rect 18544 13866 18596 13872
rect 18556 13794 18584 13866
rect 18544 13788 18596 13794
rect 18544 13730 18596 13736
rect 18820 13788 18872 13794
rect 18820 13730 18872 13736
rect 18452 13720 18504 13726
rect 18452 13662 18504 13668
rect 18464 13386 18492 13662
rect 15968 13380 16020 13386
rect 15968 13322 16020 13328
rect 17808 13380 17860 13386
rect 17808 13322 17860 13328
rect 18452 13380 18504 13386
rect 18452 13322 18504 13328
rect 17256 13312 17308 13318
rect 17256 13254 17308 13260
rect 15876 12496 15928 12502
rect 15876 12438 15928 12444
rect 15888 10598 15916 12438
rect 16336 12020 16388 12026
rect 16336 11962 16388 11968
rect 16348 11686 16376 11962
rect 16336 11680 16388 11686
rect 16336 11622 16388 11628
rect 15876 10592 15928 10598
rect 15876 10534 15928 10540
rect 16980 10320 17032 10326
rect 16980 10262 17032 10268
rect 16992 10122 17020 10262
rect 16980 10116 17032 10122
rect 16980 10058 17032 10064
rect 15692 9776 15744 9782
rect 15692 9718 15744 9724
rect 15784 9776 15836 9782
rect 15784 9718 15836 9724
rect 15600 9504 15652 9510
rect 15600 9446 15652 9452
rect 16428 9436 16480 9442
rect 16428 9378 16480 9384
rect 15324 9368 15376 9374
rect 15324 9310 15376 9316
rect 15232 9232 15284 9238
rect 15232 9174 15284 9180
rect 15244 8898 15272 9174
rect 15336 9034 15364 9310
rect 16440 9034 16468 9378
rect 16520 9300 16572 9306
rect 16520 9242 16572 9248
rect 16532 9034 16560 9242
rect 15324 9028 15376 9034
rect 15324 8970 15376 8976
rect 16428 9028 16480 9034
rect 16428 8970 16480 8976
rect 16520 9028 16572 9034
rect 16520 8970 16572 8976
rect 15232 8892 15284 8898
rect 15232 8834 15284 8840
rect 15244 8336 15272 8834
rect 16440 8354 16468 8970
rect 16532 8830 16560 8970
rect 16520 8824 16572 8830
rect 16520 8766 16572 8772
rect 15324 8348 15376 8354
rect 15244 8308 15324 8336
rect 15244 7946 15272 8308
rect 15324 8290 15376 8296
rect 15600 8348 15652 8354
rect 15600 8290 15652 8296
rect 16428 8348 16480 8354
rect 16428 8290 16480 8296
rect 15232 7940 15284 7946
rect 15232 7882 15284 7888
rect 15612 7878 15640 8290
rect 15692 8280 15744 8286
rect 15692 8222 15744 8228
rect 15600 7872 15652 7878
rect 15600 7814 15652 7820
rect 15612 7402 15640 7814
rect 15704 7606 15732 8222
rect 15876 7736 15928 7742
rect 15876 7678 15928 7684
rect 15784 7668 15836 7674
rect 15784 7610 15836 7616
rect 15692 7600 15744 7606
rect 15692 7542 15744 7548
rect 15600 7396 15652 7402
rect 15600 7338 15652 7344
rect 15048 7056 15100 7062
rect 15048 6998 15100 7004
rect 15060 6314 15088 6998
rect 15612 6790 15640 7338
rect 15704 7198 15732 7542
rect 15692 7192 15744 7198
rect 15692 7134 15744 7140
rect 15600 6784 15652 6790
rect 15600 6726 15652 6732
rect 15692 6784 15744 6790
rect 15692 6726 15744 6732
rect 15704 6654 15732 6726
rect 15140 6648 15192 6654
rect 15140 6590 15192 6596
rect 15692 6648 15744 6654
rect 15692 6590 15744 6596
rect 15152 6518 15180 6590
rect 15796 6586 15824 7610
rect 15232 6580 15284 6586
rect 15232 6522 15284 6528
rect 15784 6580 15836 6586
rect 15784 6522 15836 6528
rect 15140 6512 15192 6518
rect 15140 6454 15192 6460
rect 15048 6308 15100 6314
rect 15048 6250 15100 6256
rect 14956 5560 15008 5566
rect 14956 5502 15008 5508
rect 14588 5220 14640 5226
rect 14588 5162 14640 5168
rect 14600 4886 14628 5162
rect 15060 5090 15088 6250
rect 15244 6246 15272 6522
rect 15232 6240 15284 6246
rect 15232 6182 15284 6188
rect 15232 6104 15284 6110
rect 15232 6046 15284 6052
rect 15140 5560 15192 5566
rect 15140 5502 15192 5508
rect 15152 5158 15180 5502
rect 15244 5226 15272 6046
rect 15600 5696 15652 5702
rect 15600 5638 15652 5644
rect 15612 5566 15640 5638
rect 15888 5566 15916 7678
rect 16152 7260 16204 7266
rect 16152 7202 16204 7208
rect 16164 6858 16192 7202
rect 16152 6852 16204 6858
rect 16152 6794 16204 6800
rect 16060 6716 16112 6722
rect 16060 6658 16112 6664
rect 16072 6178 16100 6658
rect 16164 6586 16192 6794
rect 16152 6580 16204 6586
rect 16152 6522 16204 6528
rect 16060 6172 16112 6178
rect 16060 6114 16112 6120
rect 15968 6104 16020 6110
rect 15968 6046 16020 6052
rect 15980 5770 16008 6046
rect 16072 5770 16100 6114
rect 16532 6110 16560 8766
rect 16520 6104 16572 6110
rect 16520 6046 16572 6052
rect 16244 5968 16296 5974
rect 16244 5910 16296 5916
rect 16256 5770 16284 5910
rect 15968 5764 16020 5770
rect 15968 5706 16020 5712
rect 16060 5764 16112 5770
rect 16060 5706 16112 5712
rect 16244 5764 16296 5770
rect 16244 5706 16296 5712
rect 15600 5560 15652 5566
rect 15600 5502 15652 5508
rect 15876 5560 15928 5566
rect 15876 5502 15928 5508
rect 15232 5220 15284 5226
rect 15232 5162 15284 5168
rect 15140 5152 15192 5158
rect 15140 5094 15192 5100
rect 15048 5084 15100 5090
rect 15048 5026 15100 5032
rect 14588 4880 14640 4886
rect 14588 4822 14640 4828
rect 15060 4614 15088 5026
rect 15152 4682 15180 5094
rect 15888 5090 15916 5502
rect 15876 5084 15928 5090
rect 15876 5026 15928 5032
rect 15888 4682 15916 5026
rect 15980 5022 16008 5706
rect 17072 5492 17124 5498
rect 17072 5434 17124 5440
rect 15968 5016 16020 5022
rect 15968 4958 16020 4964
rect 15140 4676 15192 4682
rect 15140 4618 15192 4624
rect 15876 4676 15928 4682
rect 15876 4618 15928 4624
rect 15048 4608 15100 4614
rect 15048 4550 15100 4556
rect 15980 4546 16008 4958
rect 16152 4880 16204 4886
rect 16152 4822 16204 4828
rect 16164 4682 16192 4822
rect 16152 4676 16204 4682
rect 16152 4618 16204 4624
rect 15968 4540 16020 4546
rect 15968 4482 16020 4488
rect 15508 4336 15560 4342
rect 15508 4278 15560 4284
rect 14496 4064 14548 4070
rect 14496 4006 14548 4012
rect 15232 4064 15284 4070
rect 15232 4006 15284 4012
rect 15244 3594 15272 4006
rect 15520 3934 15548 4278
rect 15968 4064 16020 4070
rect 15968 4006 16020 4012
rect 15508 3928 15560 3934
rect 15508 3870 15560 3876
rect 15876 3928 15928 3934
rect 15876 3870 15928 3876
rect 15232 3588 15284 3594
rect 15232 3530 15284 3536
rect 15520 3322 15548 3870
rect 15888 3594 15916 3870
rect 15876 3588 15928 3594
rect 15876 3530 15928 3536
rect 15980 3526 16008 4006
rect 17084 3934 17112 5434
rect 17268 4585 17296 13254
rect 17820 13182 17848 13322
rect 17808 13176 17860 13182
rect 17808 13118 17860 13124
rect 17440 13108 17492 13114
rect 17440 13050 17492 13056
rect 17452 12774 17480 13050
rect 17440 12768 17492 12774
rect 17440 12710 17492 12716
rect 17452 12298 17480 12710
rect 18556 12706 18584 13730
rect 18728 13652 18780 13658
rect 18728 13594 18780 13600
rect 18636 13584 18688 13590
rect 18636 13526 18688 13532
rect 18648 13318 18676 13526
rect 18740 13386 18768 13594
rect 18832 13386 18860 13730
rect 19292 13590 19320 14206
rect 19384 13930 19412 16246
rect 19936 14338 19964 19034
rect 20120 18622 20148 19306
rect 20108 18616 20160 18622
rect 20108 18558 20160 18564
rect 20304 18214 20332 19646
rect 20384 18616 20436 18622
rect 20384 18558 20436 18564
rect 20396 18282 20424 18558
rect 20384 18276 20436 18282
rect 20384 18218 20436 18224
rect 20292 18208 20344 18214
rect 20292 18150 20344 18156
rect 20304 17602 20332 18150
rect 20488 18146 20516 19714
rect 20476 18140 20528 18146
rect 20476 18082 20528 18088
rect 20488 17738 20516 18082
rect 20476 17732 20528 17738
rect 20476 17674 20528 17680
rect 20292 17596 20344 17602
rect 20292 17538 20344 17544
rect 20476 17120 20528 17126
rect 20476 17062 20528 17068
rect 20292 16848 20344 16854
rect 20292 16790 20344 16796
rect 20304 16310 20332 16790
rect 20488 16650 20516 17062
rect 20672 17058 20700 19850
rect 20948 19710 20976 20054
rect 20936 19704 20988 19710
rect 21224 19681 21252 20598
rect 20936 19646 20988 19652
rect 21210 19672 21266 19681
rect 21210 19607 21266 19616
rect 21408 19166 21436 20598
rect 21396 19160 21448 19166
rect 21396 19102 21448 19108
rect 21408 18826 21436 19102
rect 21396 18820 21448 18826
rect 21396 18762 21448 18768
rect 20752 18072 20804 18078
rect 20752 18014 20804 18020
rect 20764 17534 20792 18014
rect 20752 17528 20804 17534
rect 20752 17470 20804 17476
rect 21120 17528 21172 17534
rect 21120 17470 21172 17476
rect 21028 17460 21080 17466
rect 21028 17402 21080 17408
rect 20660 17052 20712 17058
rect 20660 16994 20712 17000
rect 20672 16650 20700 16994
rect 20476 16644 20528 16650
rect 20476 16586 20528 16592
rect 20660 16644 20712 16650
rect 20660 16586 20712 16592
rect 20292 16304 20344 16310
rect 20292 16246 20344 16252
rect 20672 16038 20700 16586
rect 20660 16032 20712 16038
rect 20660 15974 20712 15980
rect 20200 15896 20252 15902
rect 20200 15838 20252 15844
rect 20212 15494 20240 15838
rect 20292 15828 20344 15834
rect 20292 15770 20344 15776
rect 20304 15562 20332 15770
rect 20292 15556 20344 15562
rect 20292 15498 20344 15504
rect 20200 15488 20252 15494
rect 20200 15430 20252 15436
rect 20212 14406 20240 15430
rect 20672 15426 20700 15974
rect 21040 15970 21068 17402
rect 21132 16990 21160 17470
rect 21500 17126 21528 21432
rect 21684 21410 21712 22842
rect 21764 22288 21816 22294
rect 21764 22230 21816 22236
rect 21776 21750 21804 22230
rect 21764 21744 21816 21750
rect 21764 21686 21816 21692
rect 21672 21404 21724 21410
rect 21672 21346 21724 21352
rect 21684 20730 21712 21346
rect 21776 21342 21804 21686
rect 21764 21336 21816 21342
rect 21764 21278 21816 21284
rect 21776 21002 21804 21278
rect 21764 20996 21816 21002
rect 21764 20938 21816 20944
rect 21672 20724 21724 20730
rect 21672 20666 21724 20672
rect 22040 20724 22092 20730
rect 22040 20666 22092 20672
rect 21764 20384 21816 20390
rect 21764 20326 21816 20332
rect 21672 20112 21724 20118
rect 21672 20054 21724 20060
rect 21684 19642 21712 20054
rect 21776 19914 21804 20326
rect 22052 20118 22080 20666
rect 22132 20316 22184 20322
rect 22132 20258 22184 20264
rect 22040 20112 22092 20118
rect 22040 20054 22092 20060
rect 21764 19908 21816 19914
rect 21764 19850 21816 19856
rect 22052 19846 22080 20054
rect 22144 19914 22172 20258
rect 22132 19908 22184 19914
rect 22132 19850 22184 19856
rect 22040 19840 22092 19846
rect 22040 19782 22092 19788
rect 21856 19704 21908 19710
rect 21856 19646 21908 19652
rect 21672 19636 21724 19642
rect 21672 19578 21724 19584
rect 21868 19166 21896 19646
rect 22224 19228 22276 19234
rect 22224 19170 22276 19176
rect 21856 19160 21908 19166
rect 21856 19102 21908 19108
rect 21868 18690 21896 19102
rect 22236 18826 22264 19170
rect 22224 18820 22276 18826
rect 22224 18762 22276 18768
rect 21856 18684 21908 18690
rect 21856 18626 21908 18632
rect 22236 18554 22264 18762
rect 22224 18548 22276 18554
rect 22224 18490 22276 18496
rect 22328 17777 22356 27315
rect 24064 26640 24116 26646
rect 24064 26582 24116 26588
rect 23604 26436 23656 26442
rect 23604 26378 23656 26384
rect 23512 26096 23564 26102
rect 23512 26038 23564 26044
rect 22868 25688 22920 25694
rect 22868 25630 22920 25636
rect 22880 25354 22908 25630
rect 22868 25348 22920 25354
rect 22868 25290 22920 25296
rect 22408 25212 22460 25218
rect 22408 25154 22460 25160
rect 22420 24470 22448 25154
rect 22880 24674 22908 25290
rect 23420 25144 23472 25150
rect 23420 25086 23472 25092
rect 23236 24804 23288 24810
rect 23236 24746 23288 24752
rect 22868 24668 22920 24674
rect 22868 24610 22920 24616
rect 22408 24464 22460 24470
rect 22408 24406 22460 24412
rect 22420 24198 22448 24406
rect 22880 24266 22908 24610
rect 22868 24260 22920 24266
rect 22868 24202 22920 24208
rect 22408 24192 22460 24198
rect 22408 24134 22460 24140
rect 23248 22974 23276 24746
rect 23432 23994 23460 25086
rect 23524 25014 23552 26038
rect 23512 25008 23564 25014
rect 23512 24950 23564 24956
rect 23524 24810 23552 24950
rect 23512 24804 23564 24810
rect 23512 24746 23564 24752
rect 23616 24266 23644 26378
rect 24076 26306 24104 26582
rect 23696 26300 23748 26306
rect 23696 26242 23748 26248
rect 24064 26300 24116 26306
rect 24064 26242 24116 26248
rect 23708 26102 23736 26242
rect 23696 26096 23748 26102
rect 23696 26038 23748 26044
rect 24076 25200 24104 26242
rect 24248 25552 24300 25558
rect 24248 25494 24300 25500
rect 24156 25212 24208 25218
rect 24076 25172 24156 25200
rect 24076 24810 24104 25172
rect 24156 25154 24208 25160
rect 24260 25082 24288 25494
rect 24248 25076 24300 25082
rect 24248 25018 24300 25024
rect 24064 24804 24116 24810
rect 24064 24746 24116 24752
rect 23604 24260 23656 24266
rect 23604 24202 23656 24208
rect 24076 24062 24104 24746
rect 24064 24056 24116 24062
rect 24064 23998 24116 24004
rect 23420 23988 23472 23994
rect 23420 23930 23472 23936
rect 23236 22968 23288 22974
rect 23236 22910 23288 22916
rect 22776 22492 22828 22498
rect 22776 22434 22828 22440
rect 22408 22424 22460 22430
rect 22408 22366 22460 22372
rect 22420 22022 22448 22366
rect 22592 22288 22644 22294
rect 22592 22230 22644 22236
rect 22408 22016 22460 22022
rect 22408 21958 22460 21964
rect 22420 20390 22448 21958
rect 22604 21750 22632 22230
rect 22788 22090 22816 22434
rect 23248 22294 23276 22910
rect 23236 22288 23288 22294
rect 23236 22230 23288 22236
rect 22776 22084 22828 22090
rect 22776 22026 22828 22032
rect 23248 21954 23276 22230
rect 23236 21948 23288 21954
rect 23236 21890 23288 21896
rect 23144 21812 23196 21818
rect 23144 21754 23196 21760
rect 22592 21744 22644 21750
rect 22592 21686 22644 21692
rect 22604 21410 22632 21686
rect 23156 21478 23184 21754
rect 22776 21472 22828 21478
rect 22776 21414 22828 21420
rect 23144 21472 23196 21478
rect 23144 21414 23196 21420
rect 22592 21404 22644 21410
rect 22592 21346 22644 21352
rect 22788 21002 22816 21414
rect 23144 21336 23196 21342
rect 23144 21278 23196 21284
rect 22776 20996 22828 21002
rect 22776 20938 22828 20944
rect 23156 20662 23184 21278
rect 23144 20656 23196 20662
rect 23144 20598 23196 20604
rect 22408 20384 22460 20390
rect 22408 20326 22460 20332
rect 22420 19302 22448 20326
rect 23156 19681 23184 20598
rect 23248 20458 23276 21890
rect 23432 21342 23460 23930
rect 24156 23376 24208 23382
rect 24156 23318 24208 23324
rect 24168 23042 24196 23318
rect 24156 23036 24208 23042
rect 24156 22978 24208 22984
rect 24260 23024 24288 25018
rect 24352 24713 24380 27315
rect 26320 27320 26460 27735
rect 26320 27315 26364 27320
rect 25444 27262 25496 27268
rect 26416 27315 26460 27320
rect 26364 27262 26416 27268
rect 24432 26096 24484 26102
rect 24432 26038 24484 26044
rect 24338 24704 24394 24713
rect 24444 24674 24472 26038
rect 25350 25112 25406 25121
rect 24708 25076 24760 25082
rect 25350 25047 25406 25056
rect 24708 25018 24760 25024
rect 24338 24639 24394 24648
rect 24432 24668 24484 24674
rect 24432 24610 24484 24616
rect 24444 23926 24472 24610
rect 24720 24606 24748 25018
rect 24708 24600 24760 24606
rect 24708 24542 24760 24548
rect 24432 23920 24484 23926
rect 24484 23868 24564 23874
rect 24432 23862 24564 23868
rect 24444 23846 24564 23862
rect 24432 23036 24484 23042
rect 24260 22996 24432 23024
rect 24260 22634 24288 22996
rect 24432 22978 24484 22984
rect 24432 22900 24484 22906
rect 24432 22842 24484 22848
rect 24444 22673 24472 22842
rect 24430 22664 24486 22673
rect 24248 22628 24300 22634
rect 24430 22599 24486 22608
rect 24248 22570 24300 22576
rect 24432 22492 24484 22498
rect 24536 22480 24564 23846
rect 24720 23722 24748 24542
rect 24708 23716 24760 23722
rect 24708 23658 24760 23664
rect 24708 22900 24760 22906
rect 24708 22842 24760 22848
rect 24720 22566 24748 22842
rect 24708 22560 24760 22566
rect 24708 22502 24760 22508
rect 24484 22452 24564 22480
rect 24432 22434 24484 22440
rect 24248 22424 24300 22430
rect 24248 22366 24300 22372
rect 23880 22356 23932 22362
rect 23880 22298 23932 22304
rect 23892 21750 23920 22298
rect 24260 21954 24288 22366
rect 24248 21948 24300 21954
rect 24248 21890 24300 21896
rect 23880 21744 23932 21750
rect 23880 21686 23932 21692
rect 24444 21546 24472 22434
rect 24524 21812 24576 21818
rect 24524 21754 24576 21760
rect 24432 21540 24484 21546
rect 24432 21482 24484 21488
rect 23512 21404 23564 21410
rect 23512 21346 23564 21352
rect 23696 21404 23748 21410
rect 23696 21346 23748 21352
rect 23420 21336 23472 21342
rect 23420 21278 23472 21284
rect 23328 21268 23380 21274
rect 23328 21210 23380 21216
rect 23340 20662 23368 21210
rect 23524 21002 23552 21346
rect 23512 20996 23564 21002
rect 23512 20938 23564 20944
rect 23708 20730 23736 21346
rect 24536 20866 24564 21754
rect 24720 21546 24748 22502
rect 24708 21540 24760 21546
rect 24708 21482 24760 21488
rect 24616 21200 24668 21206
rect 24616 21142 24668 21148
rect 24524 20860 24576 20866
rect 24524 20802 24576 20808
rect 24628 20798 24656 21142
rect 24616 20792 24668 20798
rect 24616 20734 24668 20740
rect 23696 20724 23748 20730
rect 23696 20666 23748 20672
rect 24156 20724 24208 20730
rect 24156 20666 24208 20672
rect 23328 20656 23380 20662
rect 23328 20598 23380 20604
rect 23236 20452 23288 20458
rect 23236 20394 23288 20400
rect 23248 19778 23276 20394
rect 23236 19772 23288 19778
rect 23236 19714 23288 19720
rect 23142 19672 23198 19681
rect 23142 19607 23198 19616
rect 23156 19370 23184 19607
rect 23236 19568 23288 19574
rect 23236 19510 23288 19516
rect 23144 19364 23196 19370
rect 23144 19306 23196 19312
rect 22408 19296 22460 19302
rect 22408 19238 22460 19244
rect 22408 19160 22460 19166
rect 22408 19102 22460 19108
rect 22420 18758 22448 19102
rect 23248 19030 23276 19510
rect 23340 19234 23368 20598
rect 23972 19636 24024 19642
rect 23972 19578 24024 19584
rect 23788 19568 23840 19574
rect 23984 19522 24012 19578
rect 23840 19516 24012 19522
rect 23788 19510 24012 19516
rect 23800 19494 24012 19510
rect 23512 19364 23564 19370
rect 23512 19306 23564 19312
rect 23328 19228 23380 19234
rect 23328 19170 23380 19176
rect 23236 19024 23288 19030
rect 23236 18966 23288 18972
rect 22408 18752 22460 18758
rect 22408 18694 22460 18700
rect 22408 18480 22460 18486
rect 22408 18422 22460 18428
rect 22420 18282 22448 18422
rect 22408 18276 22460 18282
rect 22408 18218 22460 18224
rect 23248 18078 23276 18966
rect 23340 18282 23368 19170
rect 23524 18690 23552 19306
rect 23604 19024 23656 19030
rect 23604 18966 23656 18972
rect 23420 18684 23472 18690
rect 23420 18626 23472 18632
rect 23512 18684 23564 18690
rect 23512 18626 23564 18632
rect 23328 18276 23380 18282
rect 23328 18218 23380 18224
rect 23432 18146 23460 18626
rect 23420 18140 23472 18146
rect 23420 18082 23472 18088
rect 23236 18072 23288 18078
rect 23236 18014 23288 18020
rect 22314 17768 22370 17777
rect 23432 17738 23460 18082
rect 22314 17703 22370 17712
rect 23420 17732 23472 17738
rect 23420 17674 23472 17680
rect 23524 17618 23552 18626
rect 23616 18622 23644 18966
rect 23604 18616 23656 18622
rect 23604 18558 23656 18564
rect 23800 18214 23828 19494
rect 24064 19296 24116 19302
rect 24064 19238 24116 19244
rect 23972 18616 24024 18622
rect 23972 18558 24024 18564
rect 23788 18208 23840 18214
rect 23788 18150 23840 18156
rect 23432 17590 23552 17618
rect 21488 17120 21540 17126
rect 21488 17062 21540 17068
rect 21212 17052 21264 17058
rect 21212 16994 21264 17000
rect 21120 16984 21172 16990
rect 21120 16926 21172 16932
rect 21132 16650 21160 16926
rect 21120 16644 21172 16650
rect 21120 16586 21172 16592
rect 21224 16582 21252 16994
rect 23236 16916 23288 16922
rect 23236 16858 23288 16864
rect 23144 16848 23196 16854
rect 23144 16790 23196 16796
rect 23156 16582 23184 16790
rect 21212 16576 21264 16582
rect 21212 16518 21264 16524
rect 23144 16576 23196 16582
rect 23144 16518 23196 16524
rect 23248 16446 23276 16858
rect 23328 16508 23380 16514
rect 23328 16450 23380 16456
rect 23236 16440 23288 16446
rect 23236 16382 23288 16388
rect 21488 16304 21540 16310
rect 21488 16246 21540 16252
rect 21028 15964 21080 15970
rect 21028 15906 21080 15912
rect 21040 15562 21068 15906
rect 21500 15834 21528 16246
rect 22684 15964 22736 15970
rect 22684 15906 22736 15912
rect 21488 15828 21540 15834
rect 21488 15770 21540 15776
rect 21028 15556 21080 15562
rect 21028 15498 21080 15504
rect 20660 15420 20712 15426
rect 20660 15362 20712 15368
rect 20476 14672 20528 14678
rect 20476 14614 20528 14620
rect 20200 14400 20252 14406
rect 20200 14342 20252 14348
rect 19924 14332 19976 14338
rect 19924 14274 19976 14280
rect 19372 13924 19424 13930
rect 19372 13866 19424 13872
rect 19188 13584 19240 13590
rect 19188 13526 19240 13532
rect 19280 13584 19332 13590
rect 19280 13526 19332 13532
rect 18728 13380 18780 13386
rect 18728 13322 18780 13328
rect 18820 13380 18872 13386
rect 18820 13322 18872 13328
rect 18636 13312 18688 13318
rect 18636 13254 18688 13260
rect 19200 13182 19228 13526
rect 19292 13318 19320 13526
rect 19384 13386 19412 13866
rect 19936 13726 19964 14274
rect 20488 14270 20516 14614
rect 20568 14400 20620 14406
rect 20568 14342 20620 14348
rect 20476 14264 20528 14270
rect 20476 14206 20528 14212
rect 20488 13862 20516 14206
rect 20580 13930 20608 14342
rect 20568 13924 20620 13930
rect 20568 13866 20620 13872
rect 20476 13856 20528 13862
rect 20476 13798 20528 13804
rect 20384 13788 20436 13794
rect 20384 13730 20436 13736
rect 19924 13720 19976 13726
rect 19924 13662 19976 13668
rect 19372 13380 19424 13386
rect 19372 13322 19424 13328
rect 19280 13312 19332 13318
rect 19280 13254 19332 13260
rect 20396 13182 20424 13730
rect 20488 13386 20516 13798
rect 21500 13697 21528 15770
rect 22696 15222 22724 15906
rect 23248 15766 23276 16382
rect 23236 15760 23288 15766
rect 23236 15702 23288 15708
rect 22776 15352 22828 15358
rect 22776 15294 22828 15300
rect 22684 15216 22736 15222
rect 22684 15158 22736 15164
rect 22316 14808 22368 14814
rect 22316 14750 22368 14756
rect 21672 14332 21724 14338
rect 21672 14274 21724 14280
rect 21684 13794 21712 14274
rect 22328 13930 22356 14750
rect 22316 13924 22368 13930
rect 22316 13866 22368 13872
rect 21672 13788 21724 13794
rect 21672 13730 21724 13736
rect 22132 13788 22184 13794
rect 22132 13730 22184 13736
rect 21948 13720 22000 13726
rect 21486 13688 21542 13697
rect 21948 13662 22000 13668
rect 21486 13623 21542 13632
rect 21212 13584 21264 13590
rect 21212 13526 21264 13532
rect 20476 13380 20528 13386
rect 20476 13322 20528 13328
rect 19188 13176 19240 13182
rect 19188 13118 19240 13124
rect 20016 13176 20068 13182
rect 20016 13118 20068 13124
rect 20384 13176 20436 13182
rect 20384 13118 20436 13124
rect 18864 12940 19184 12960
rect 18864 12938 18876 12940
rect 18932 12938 18956 12940
rect 19012 12938 19036 12940
rect 19092 12938 19116 12940
rect 19172 12938 19184 12940
rect 18864 12886 18870 12938
rect 18932 12886 18934 12938
rect 19114 12886 19116 12938
rect 19178 12886 19184 12938
rect 18864 12884 18876 12886
rect 18932 12884 18956 12886
rect 19012 12884 19036 12886
rect 19092 12884 19116 12886
rect 19172 12884 19184 12886
rect 18864 12864 19184 12884
rect 17532 12700 17584 12706
rect 17532 12642 17584 12648
rect 18544 12700 18596 12706
rect 18544 12642 18596 12648
rect 17440 12292 17492 12298
rect 17440 12234 17492 12240
rect 17544 12230 17572 12642
rect 17716 12496 17768 12502
rect 17716 12438 17768 12444
rect 17728 12298 17756 12438
rect 17716 12292 17768 12298
rect 17716 12234 17768 12240
rect 17532 12224 17584 12230
rect 17532 12166 17584 12172
rect 17348 10116 17400 10122
rect 17348 10058 17400 10064
rect 17360 9782 17388 10058
rect 17348 9776 17400 9782
rect 17348 9718 17400 9724
rect 17440 9776 17492 9782
rect 17440 9718 17492 9724
rect 17452 7334 17480 9718
rect 17728 9442 17756 12234
rect 18864 11852 19184 11872
rect 18864 11850 18876 11852
rect 18932 11850 18956 11852
rect 19012 11850 19036 11852
rect 19092 11850 19116 11852
rect 19172 11850 19184 11852
rect 18864 11798 18870 11850
rect 18932 11798 18934 11850
rect 19114 11798 19116 11850
rect 19178 11798 19184 11850
rect 18864 11796 18876 11798
rect 18932 11796 18956 11798
rect 19012 11796 19036 11798
rect 19092 11796 19116 11798
rect 19172 11796 19184 11798
rect 18864 11776 19184 11796
rect 19280 11136 19332 11142
rect 19280 11078 19332 11084
rect 18728 11000 18780 11006
rect 18728 10942 18780 10948
rect 17992 10932 18044 10938
rect 17992 10874 18044 10880
rect 18004 10530 18032 10874
rect 17992 10524 18044 10530
rect 17992 10466 18044 10472
rect 18360 10524 18412 10530
rect 18360 10466 18412 10472
rect 18544 10524 18596 10530
rect 18544 10466 18596 10472
rect 18004 9782 18032 10466
rect 18084 10456 18136 10462
rect 18084 10398 18136 10404
rect 17992 9776 18044 9782
rect 17992 9718 18044 9724
rect 18096 9578 18124 10398
rect 18372 10054 18400 10466
rect 18556 10122 18584 10466
rect 18740 10326 18768 10942
rect 18864 10764 19184 10784
rect 18864 10762 18876 10764
rect 18932 10762 18956 10764
rect 19012 10762 19036 10764
rect 19092 10762 19116 10764
rect 19172 10762 19184 10764
rect 18864 10710 18870 10762
rect 18932 10710 18934 10762
rect 19114 10710 19116 10762
rect 19178 10710 19184 10762
rect 18864 10708 18876 10710
rect 18932 10708 18956 10710
rect 19012 10708 19036 10710
rect 19092 10708 19116 10710
rect 19172 10708 19184 10710
rect 18864 10688 19184 10708
rect 19292 10666 19320 11078
rect 19372 11000 19424 11006
rect 19372 10942 19424 10948
rect 19280 10660 19332 10666
rect 19280 10602 19332 10608
rect 18728 10320 18780 10326
rect 18728 10262 18780 10268
rect 19096 10320 19148 10326
rect 19096 10262 19148 10268
rect 18544 10116 18596 10122
rect 18544 10058 18596 10064
rect 18360 10048 18412 10054
rect 18360 9990 18412 9996
rect 18084 9572 18136 9578
rect 18004 9532 18084 9560
rect 17716 9436 17768 9442
rect 17716 9378 17768 9384
rect 17716 8824 17768 8830
rect 17716 8766 17768 8772
rect 17728 8354 17756 8766
rect 17716 8348 17768 8354
rect 17716 8290 17768 8296
rect 17624 7804 17676 7810
rect 17624 7746 17676 7752
rect 17636 7713 17664 7746
rect 17622 7704 17678 7713
rect 17622 7639 17678 7648
rect 17532 7600 17584 7606
rect 17532 7542 17584 7548
rect 17624 7600 17676 7606
rect 17624 7542 17676 7548
rect 17440 7328 17492 7334
rect 17440 7270 17492 7276
rect 17452 6518 17480 7270
rect 17544 7198 17572 7542
rect 17636 7266 17664 7542
rect 17728 7402 17756 8290
rect 17808 8144 17860 8150
rect 17808 8086 17860 8092
rect 17820 7946 17848 8086
rect 17808 7940 17860 7946
rect 17808 7882 17860 7888
rect 17900 7668 17952 7674
rect 17900 7610 17952 7616
rect 17716 7396 17768 7402
rect 17716 7338 17768 7344
rect 17624 7260 17676 7266
rect 17624 7202 17676 7208
rect 17532 7192 17584 7198
rect 17532 7134 17584 7140
rect 17440 6512 17492 6518
rect 17440 6454 17492 6460
rect 17624 6172 17676 6178
rect 17624 6114 17676 6120
rect 17440 6036 17492 6042
rect 17440 5978 17492 5984
rect 17452 5566 17480 5978
rect 17636 5770 17664 6114
rect 17808 6104 17860 6110
rect 17808 6046 17860 6052
rect 17624 5764 17676 5770
rect 17624 5706 17676 5712
rect 17440 5560 17492 5566
rect 17440 5502 17492 5508
rect 17820 5226 17848 6046
rect 17912 5770 17940 7610
rect 18004 6790 18032 9532
rect 18084 9514 18136 9520
rect 18268 8892 18320 8898
rect 18320 8852 18400 8880
rect 18268 8834 18320 8840
rect 18372 8762 18400 8852
rect 18452 8824 18504 8830
rect 18452 8766 18504 8772
rect 18360 8756 18412 8762
rect 18360 8698 18412 8704
rect 18268 8688 18320 8694
rect 18268 8630 18320 8636
rect 18280 8354 18308 8630
rect 18268 8348 18320 8354
rect 18268 8290 18320 8296
rect 18084 7668 18136 7674
rect 18084 7610 18136 7616
rect 18096 7402 18124 7610
rect 18084 7396 18136 7402
rect 18084 7338 18136 7344
rect 18280 7198 18308 8290
rect 18360 7804 18412 7810
rect 18360 7746 18412 7752
rect 18268 7192 18320 7198
rect 18268 7134 18320 7140
rect 18176 7124 18228 7130
rect 18176 7066 18228 7072
rect 17992 6784 18044 6790
rect 17992 6726 18044 6732
rect 18004 6194 18032 6726
rect 18004 6166 18124 6194
rect 17992 6104 18044 6110
rect 17992 6046 18044 6052
rect 17900 5764 17952 5770
rect 17900 5706 17952 5712
rect 18004 5650 18032 6046
rect 17912 5622 18032 5650
rect 18096 5956 18124 6166
rect 18188 6110 18216 7066
rect 18176 6104 18228 6110
rect 18176 6046 18228 6052
rect 18176 5968 18228 5974
rect 18096 5928 18176 5956
rect 17912 5498 17940 5622
rect 17992 5560 18044 5566
rect 17992 5502 18044 5508
rect 17900 5492 17952 5498
rect 17900 5434 17952 5440
rect 17808 5220 17860 5226
rect 17808 5162 17860 5168
rect 18004 5022 18032 5502
rect 18096 5158 18124 5928
rect 18176 5910 18228 5916
rect 18372 5634 18400 7746
rect 18464 7742 18492 8766
rect 18452 7736 18504 7742
rect 18452 7678 18504 7684
rect 18556 6654 18584 10058
rect 18740 9442 18768 10262
rect 19108 9850 19136 10262
rect 19292 9918 19320 10602
rect 19280 9912 19332 9918
rect 19280 9854 19332 9860
rect 19096 9844 19148 9850
rect 19096 9786 19148 9792
rect 18864 9676 19184 9696
rect 18864 9674 18876 9676
rect 18932 9674 18956 9676
rect 19012 9674 19036 9676
rect 19092 9674 19116 9676
rect 19172 9674 19184 9676
rect 18864 9622 18870 9674
rect 18932 9622 18934 9674
rect 19114 9622 19116 9674
rect 19178 9622 19184 9674
rect 18864 9620 18876 9622
rect 18932 9620 18956 9622
rect 19012 9620 19036 9622
rect 19092 9620 19116 9622
rect 19172 9620 19184 9622
rect 18864 9600 19184 9620
rect 19280 9504 19332 9510
rect 19280 9446 19332 9452
rect 18728 9436 18780 9442
rect 18728 9378 18780 9384
rect 18912 9436 18964 9442
rect 18912 9378 18964 9384
rect 18740 9034 18768 9378
rect 18728 9028 18780 9034
rect 18728 8970 18780 8976
rect 18924 8966 18952 9378
rect 19292 9034 19320 9446
rect 19384 9442 19412 10942
rect 19740 9912 19792 9918
rect 19740 9854 19792 9860
rect 19752 9578 19780 9854
rect 19740 9572 19792 9578
rect 19740 9514 19792 9520
rect 19372 9436 19424 9442
rect 19372 9378 19424 9384
rect 19280 9028 19332 9034
rect 19280 8970 19332 8976
rect 18912 8960 18964 8966
rect 18912 8902 18964 8908
rect 18864 8588 19184 8608
rect 18864 8586 18876 8588
rect 18932 8586 18956 8588
rect 19012 8586 19036 8588
rect 19092 8586 19116 8588
rect 19172 8586 19184 8588
rect 18864 8534 18870 8586
rect 18932 8534 18934 8586
rect 19114 8534 19116 8586
rect 19178 8534 19184 8586
rect 18864 8532 18876 8534
rect 18932 8532 18956 8534
rect 19012 8532 19036 8534
rect 19092 8532 19116 8534
rect 19172 8532 19184 8534
rect 18864 8512 19184 8532
rect 18636 8144 18688 8150
rect 18636 8086 18688 8092
rect 18820 8144 18872 8150
rect 18820 8086 18872 8092
rect 18648 7742 18676 8086
rect 18832 7810 18860 8086
rect 20028 7810 20056 13118
rect 20488 12842 20516 13322
rect 21224 13250 21252 13526
rect 21960 13386 21988 13662
rect 22144 13386 22172 13730
rect 21948 13380 22000 13386
rect 21948 13322 22000 13328
rect 22132 13380 22184 13386
rect 22132 13322 22184 13328
rect 21856 13312 21908 13318
rect 21856 13254 21908 13260
rect 21212 13244 21264 13250
rect 21212 13186 21264 13192
rect 21868 13182 21896 13254
rect 21672 13176 21724 13182
rect 21672 13118 21724 13124
rect 21856 13176 21908 13182
rect 21856 13118 21908 13124
rect 22224 13176 22276 13182
rect 22328 13164 22356 13866
rect 22276 13136 22356 13164
rect 22224 13118 22276 13124
rect 20660 13108 20712 13114
rect 20660 13050 20712 13056
rect 20672 12842 20700 13050
rect 21684 13046 21712 13118
rect 21672 13040 21724 13046
rect 21672 12982 21724 12988
rect 20476 12836 20528 12842
rect 20476 12778 20528 12784
rect 20660 12836 20712 12842
rect 20660 12778 20712 12784
rect 20488 12230 20516 12778
rect 20672 12298 20700 12778
rect 21684 12706 21712 12982
rect 21868 12706 21896 13118
rect 21948 13108 22000 13114
rect 21948 13050 22000 13056
rect 21672 12700 21724 12706
rect 21672 12642 21724 12648
rect 21856 12700 21908 12706
rect 21856 12642 21908 12648
rect 20660 12292 20712 12298
rect 20660 12234 20712 12240
rect 20476 12224 20528 12230
rect 20476 12166 20528 12172
rect 21684 12026 21712 12642
rect 21868 12162 21896 12642
rect 21960 12638 21988 13050
rect 22696 12706 22724 15158
rect 22788 14882 22816 15294
rect 23248 15222 23276 15702
rect 23236 15216 23288 15222
rect 23236 15158 23288 15164
rect 22776 14876 22828 14882
rect 22776 14818 22828 14824
rect 23052 14876 23104 14882
rect 23052 14818 23104 14824
rect 22788 14270 22816 14818
rect 22776 14264 22828 14270
rect 22776 14206 22828 14212
rect 23064 14134 23092 14818
rect 23248 14814 23276 15158
rect 23340 14882 23368 16450
rect 23432 16038 23460 17590
rect 23512 17528 23564 17534
rect 23696 17528 23748 17534
rect 23564 17488 23696 17516
rect 23512 17470 23564 17476
rect 23420 16032 23472 16038
rect 23420 15974 23472 15980
rect 23432 14950 23460 15974
rect 23420 14944 23472 14950
rect 23420 14886 23472 14892
rect 23328 14876 23380 14882
rect 23328 14818 23380 14824
rect 23236 14808 23288 14814
rect 23236 14750 23288 14756
rect 23248 14474 23276 14750
rect 23236 14468 23288 14474
rect 23236 14410 23288 14416
rect 23340 14406 23368 14818
rect 23328 14400 23380 14406
rect 23328 14342 23380 14348
rect 23052 14128 23104 14134
rect 23052 14070 23104 14076
rect 23064 13930 23092 14070
rect 23052 13924 23104 13930
rect 23052 13866 23104 13872
rect 23064 13386 23092 13866
rect 23340 13794 23368 14342
rect 23616 14338 23644 17488
rect 23696 17470 23748 17476
rect 23800 17398 23828 18150
rect 23984 17738 24012 18558
rect 24076 18486 24104 19238
rect 24168 18826 24196 20666
rect 25168 20656 25220 20662
rect 25168 20598 25220 20604
rect 24984 19568 25036 19574
rect 24984 19510 25036 19516
rect 24996 18826 25024 19510
rect 24156 18820 24208 18826
rect 24156 18762 24208 18768
rect 24984 18820 25036 18826
rect 24984 18762 25036 18768
rect 24168 18622 24196 18762
rect 25180 18622 25208 20598
rect 24156 18616 24208 18622
rect 24156 18558 24208 18564
rect 25168 18616 25220 18622
rect 25168 18558 25220 18564
rect 24064 18480 24116 18486
rect 24064 18422 24116 18428
rect 23972 17732 24024 17738
rect 23972 17674 24024 17680
rect 23788 17392 23840 17398
rect 23788 17334 23840 17340
rect 23984 16802 24012 17674
rect 24076 17534 24104 18422
rect 24168 17670 24196 18558
rect 24432 17936 24484 17942
rect 24432 17878 24484 17884
rect 24156 17664 24208 17670
rect 24156 17606 24208 17612
rect 24064 17528 24116 17534
rect 24064 17470 24116 17476
rect 23984 16774 24104 16802
rect 24076 16650 24104 16774
rect 24064 16644 24116 16650
rect 24064 16586 24116 16592
rect 23788 16508 23840 16514
rect 23788 16450 23840 16456
rect 23696 16372 23748 16378
rect 23696 16314 23748 16320
rect 23708 15018 23736 16314
rect 23800 15358 23828 16450
rect 24076 16446 24104 16586
rect 24064 16440 24116 16446
rect 24064 16382 24116 16388
rect 24064 15828 24116 15834
rect 24064 15770 24116 15776
rect 24076 15562 24104 15770
rect 24064 15556 24116 15562
rect 24064 15498 24116 15504
rect 23788 15352 23840 15358
rect 23788 15294 23840 15300
rect 23696 15012 23748 15018
rect 23696 14954 23748 14960
rect 24064 14944 24116 14950
rect 24064 14886 24116 14892
rect 23696 14876 23748 14882
rect 23696 14818 23748 14824
rect 23420 14332 23472 14338
rect 23420 14274 23472 14280
rect 23604 14332 23656 14338
rect 23604 14274 23656 14280
rect 23432 13930 23460 14274
rect 23420 13924 23472 13930
rect 23420 13866 23472 13872
rect 23328 13788 23380 13794
rect 23328 13730 23380 13736
rect 23052 13380 23104 13386
rect 23052 13322 23104 13328
rect 23340 13250 23368 13730
rect 23328 13244 23380 13250
rect 23328 13186 23380 13192
rect 23328 12768 23380 12774
rect 23328 12710 23380 12716
rect 22684 12700 22736 12706
rect 22684 12642 22736 12648
rect 21948 12632 22000 12638
rect 21948 12574 22000 12580
rect 21960 12298 21988 12574
rect 21948 12292 22000 12298
rect 21948 12234 22000 12240
rect 22696 12230 22724 12642
rect 22776 12632 22828 12638
rect 22776 12574 22828 12580
rect 22788 12298 22816 12574
rect 23340 12298 23368 12710
rect 23512 12564 23564 12570
rect 23512 12506 23564 12512
rect 23524 12298 23552 12506
rect 22776 12292 22828 12298
rect 22776 12234 22828 12240
rect 23328 12292 23380 12298
rect 23328 12234 23380 12240
rect 23512 12292 23564 12298
rect 23512 12234 23564 12240
rect 22684 12224 22736 12230
rect 22684 12166 22736 12172
rect 21856 12156 21908 12162
rect 21856 12098 21908 12104
rect 21672 12020 21724 12026
rect 21672 11962 21724 11968
rect 20936 10932 20988 10938
rect 20936 10874 20988 10880
rect 20948 10598 20976 10874
rect 22696 10666 22724 12166
rect 23708 12094 23736 14818
rect 23788 14264 23840 14270
rect 23788 14206 23840 14212
rect 23800 13930 23828 14206
rect 23788 13924 23840 13930
rect 23788 13866 23840 13872
rect 23800 13250 23828 13866
rect 23788 13244 23840 13250
rect 23788 13186 23840 13192
rect 23788 13108 23840 13114
rect 23788 13050 23840 13056
rect 23800 12638 23828 13050
rect 24076 12706 24104 14886
rect 24168 13386 24196 17606
rect 24444 17534 24472 17878
rect 24432 17528 24484 17534
rect 24432 17470 24484 17476
rect 24340 17052 24392 17058
rect 24340 16994 24392 17000
rect 24248 16440 24300 16446
rect 24248 16382 24300 16388
rect 24260 15902 24288 16382
rect 24248 15896 24300 15902
rect 24248 15838 24300 15844
rect 24260 15222 24288 15838
rect 24352 15290 24380 16994
rect 24984 16848 25036 16854
rect 24984 16790 25036 16796
rect 24996 16514 25024 16790
rect 24984 16508 25036 16514
rect 24984 16450 25036 16456
rect 24708 16304 24760 16310
rect 24708 16246 24760 16252
rect 24720 15902 24748 16246
rect 24708 15896 24760 15902
rect 24708 15838 24760 15844
rect 24340 15284 24392 15290
rect 24340 15226 24392 15232
rect 24892 15284 24944 15290
rect 24892 15226 24944 15232
rect 24248 15216 24300 15222
rect 24248 15158 24300 15164
rect 24352 14950 24380 15226
rect 24904 15018 24932 15226
rect 24892 15012 24944 15018
rect 24892 14954 24944 14960
rect 24340 14944 24392 14950
rect 24340 14886 24392 14892
rect 24904 14338 24932 14954
rect 24892 14332 24944 14338
rect 24892 14274 24944 14280
rect 24432 14264 24484 14270
rect 24432 14206 24484 14212
rect 24156 13380 24208 13386
rect 24156 13322 24208 13328
rect 24168 13182 24196 13322
rect 24156 13176 24208 13182
rect 24156 13118 24208 13124
rect 24168 12774 24196 13118
rect 24156 12768 24208 12774
rect 24156 12710 24208 12716
rect 24064 12700 24116 12706
rect 24064 12642 24116 12648
rect 23788 12632 23840 12638
rect 23788 12574 23840 12580
rect 23696 12088 23748 12094
rect 23696 12030 23748 12036
rect 23328 11748 23380 11754
rect 23328 11690 23380 11696
rect 22684 10660 22736 10666
rect 22684 10602 22736 10608
rect 23236 10660 23288 10666
rect 23236 10602 23288 10608
rect 20936 10592 20988 10598
rect 20936 10534 20988 10540
rect 20476 10456 20528 10462
rect 20476 10398 20528 10404
rect 20292 10320 20344 10326
rect 20292 10262 20344 10268
rect 20304 9986 20332 10262
rect 20488 10122 20516 10398
rect 20948 10122 20976 10534
rect 23052 10524 23104 10530
rect 23052 10466 23104 10472
rect 22224 10456 22276 10462
rect 22224 10398 22276 10404
rect 20476 10116 20528 10122
rect 20476 10058 20528 10064
rect 20936 10116 20988 10122
rect 20936 10058 20988 10064
rect 22236 9986 22264 10398
rect 20292 9980 20344 9986
rect 20292 9922 20344 9928
rect 22224 9980 22276 9986
rect 22224 9922 22276 9928
rect 20304 9578 20332 9922
rect 20476 9912 20528 9918
rect 20476 9854 20528 9860
rect 20292 9572 20344 9578
rect 20292 9514 20344 9520
rect 20488 9034 20516 9854
rect 21304 9844 21356 9850
rect 21304 9786 21356 9792
rect 20476 9028 20528 9034
rect 20476 8970 20528 8976
rect 21316 8830 21344 9786
rect 23064 9782 23092 10466
rect 23248 10122 23276 10602
rect 23340 10530 23368 11690
rect 23708 11618 23736 12030
rect 24076 11754 24104 12642
rect 24064 11748 24116 11754
rect 24064 11690 24116 11696
rect 24444 11618 24472 14206
rect 24708 12020 24760 12026
rect 24708 11962 24760 11968
rect 24616 11952 24668 11958
rect 24616 11894 24668 11900
rect 23696 11612 23748 11618
rect 24432 11612 24484 11618
rect 23748 11572 23828 11600
rect 23696 11554 23748 11560
rect 23800 10666 23828 11572
rect 24432 11554 24484 11560
rect 24444 11210 24472 11554
rect 24432 11204 24484 11210
rect 24432 11146 24484 11152
rect 24444 11074 24472 11146
rect 24432 11068 24484 11074
rect 24432 11010 24484 11016
rect 23788 10660 23840 10666
rect 23840 10620 23920 10648
rect 23788 10602 23840 10608
rect 23328 10524 23380 10530
rect 23328 10466 23380 10472
rect 23788 10524 23840 10530
rect 23788 10466 23840 10472
rect 23512 10456 23564 10462
rect 23512 10398 23564 10404
rect 23524 10122 23552 10398
rect 23236 10116 23288 10122
rect 23512 10116 23564 10122
rect 23288 10064 23460 10074
rect 23236 10058 23460 10064
rect 23512 10058 23564 10064
rect 23248 10046 23460 10058
rect 22224 9776 22276 9782
rect 22224 9718 22276 9724
rect 23052 9776 23104 9782
rect 23052 9718 23104 9724
rect 22236 9034 22264 9718
rect 23064 9510 23092 9718
rect 23052 9504 23104 9510
rect 23052 9446 23104 9452
rect 23432 9442 23460 10046
rect 23604 9776 23656 9782
rect 23604 9718 23656 9724
rect 23420 9436 23472 9442
rect 23420 9378 23472 9384
rect 23328 9368 23380 9374
rect 23328 9310 23380 9316
rect 23052 9300 23104 9306
rect 23052 9242 23104 9248
rect 22776 9232 22828 9238
rect 22776 9174 22828 9180
rect 22788 9034 22816 9174
rect 23064 9034 23092 9242
rect 21488 9028 21540 9034
rect 21488 8970 21540 8976
rect 22224 9028 22276 9034
rect 22224 8970 22276 8976
rect 22776 9028 22828 9034
rect 22776 8970 22828 8976
rect 23052 9028 23104 9034
rect 23052 8970 23104 8976
rect 21304 8824 21356 8830
rect 21304 8766 21356 8772
rect 20936 7940 20988 7946
rect 20936 7882 20988 7888
rect 18820 7804 18872 7810
rect 18820 7746 18872 7752
rect 20016 7804 20068 7810
rect 20016 7746 20068 7752
rect 18636 7736 18688 7742
rect 18636 7678 18688 7684
rect 19464 7736 19516 7742
rect 19464 7678 19516 7684
rect 19476 7606 19504 7678
rect 19464 7600 19516 7606
rect 19464 7542 19516 7548
rect 18864 7500 19184 7520
rect 18864 7498 18876 7500
rect 18932 7498 18956 7500
rect 19012 7498 19036 7500
rect 19092 7498 19116 7500
rect 19172 7498 19184 7500
rect 18864 7446 18870 7498
rect 18932 7446 18934 7498
rect 19114 7446 19116 7498
rect 19178 7446 19184 7498
rect 18864 7444 18876 7446
rect 18932 7444 18956 7446
rect 19012 7444 19036 7446
rect 19092 7444 19116 7446
rect 19172 7444 19184 7446
rect 18864 7424 19184 7444
rect 19476 7402 19504 7542
rect 19464 7396 19516 7402
rect 19464 7338 19516 7344
rect 20028 7266 20056 7746
rect 19648 7260 19700 7266
rect 19648 7202 19700 7208
rect 20016 7260 20068 7266
rect 20016 7202 20068 7208
rect 18636 7192 18688 7198
rect 18636 7134 18688 7140
rect 19280 7192 19332 7198
rect 19280 7134 19332 7140
rect 18544 6648 18596 6654
rect 18544 6590 18596 6596
rect 18648 6246 18676 7134
rect 19292 6858 19320 7134
rect 19660 7062 19688 7202
rect 19648 7056 19700 7062
rect 19648 6998 19700 7004
rect 19280 6852 19332 6858
rect 19280 6794 19332 6800
rect 18864 6412 19184 6432
rect 18864 6410 18876 6412
rect 18932 6410 18956 6412
rect 19012 6410 19036 6412
rect 19092 6410 19116 6412
rect 19172 6410 19184 6412
rect 18864 6358 18870 6410
rect 18932 6358 18934 6410
rect 19114 6358 19116 6410
rect 19178 6358 19184 6410
rect 18864 6356 18876 6358
rect 18932 6356 18956 6358
rect 19012 6356 19036 6358
rect 19092 6356 19116 6358
rect 19172 6356 19184 6358
rect 18864 6336 19184 6356
rect 18636 6240 18688 6246
rect 18636 6182 18688 6188
rect 18360 5628 18412 5634
rect 18360 5570 18412 5576
rect 18372 5226 18400 5570
rect 18864 5324 19184 5344
rect 18864 5322 18876 5324
rect 18932 5322 18956 5324
rect 19012 5322 19036 5324
rect 19092 5322 19116 5324
rect 19172 5322 19184 5324
rect 18864 5270 18870 5322
rect 18932 5270 18934 5322
rect 19114 5270 19116 5322
rect 19178 5270 19184 5322
rect 18864 5268 18876 5270
rect 18932 5268 18956 5270
rect 19012 5268 19036 5270
rect 19092 5268 19116 5270
rect 19172 5268 19184 5270
rect 18864 5248 19184 5268
rect 18360 5220 18412 5226
rect 18360 5162 18412 5168
rect 19292 5158 19320 6794
rect 19660 6518 19688 6998
rect 20028 6858 20056 7202
rect 20108 7192 20160 7198
rect 20108 7134 20160 7140
rect 20016 6852 20068 6858
rect 20016 6794 20068 6800
rect 20120 6586 20148 7134
rect 20384 7124 20436 7130
rect 20436 7084 20516 7112
rect 20384 7066 20436 7072
rect 20108 6580 20160 6586
rect 20108 6522 20160 6528
rect 19648 6512 19700 6518
rect 19648 6454 19700 6460
rect 19660 6314 19688 6454
rect 19648 6308 19700 6314
rect 19648 6250 19700 6256
rect 20292 6240 20344 6246
rect 20292 6182 20344 6188
rect 20304 5770 20332 6182
rect 20384 6172 20436 6178
rect 20384 6114 20436 6120
rect 20292 5764 20344 5770
rect 20292 5706 20344 5712
rect 20396 5634 20424 6114
rect 20488 5974 20516 7084
rect 20948 6654 20976 7882
rect 21316 7402 21344 8766
rect 21500 7946 21528 8970
rect 23340 8830 23368 9310
rect 23432 9034 23460 9378
rect 23616 9306 23644 9718
rect 23800 9578 23828 10466
rect 23892 10122 23920 10620
rect 24444 10530 24472 11010
rect 24432 10524 24484 10530
rect 24432 10466 24484 10472
rect 24064 10320 24116 10326
rect 24064 10262 24116 10268
rect 23880 10116 23932 10122
rect 23880 10058 23932 10064
rect 23788 9572 23840 9578
rect 23788 9514 23840 9520
rect 23696 9436 23748 9442
rect 23696 9378 23748 9384
rect 23604 9300 23656 9306
rect 23604 9242 23656 9248
rect 23708 9238 23736 9378
rect 23696 9232 23748 9238
rect 23696 9174 23748 9180
rect 23420 9028 23472 9034
rect 23420 8970 23472 8976
rect 23328 8824 23380 8830
rect 23328 8766 23380 8772
rect 23340 8490 23368 8766
rect 23328 8484 23380 8490
rect 23328 8426 23380 8432
rect 23432 8354 23460 8970
rect 23512 8756 23564 8762
rect 23512 8698 23564 8704
rect 23420 8348 23472 8354
rect 23420 8290 23472 8296
rect 23432 7946 23460 8290
rect 23524 8286 23552 8698
rect 23512 8280 23564 8286
rect 23512 8222 23564 8228
rect 21488 7940 21540 7946
rect 21488 7882 21540 7888
rect 23420 7940 23472 7946
rect 23420 7882 23472 7888
rect 21500 7742 21528 7882
rect 21488 7736 21540 7742
rect 21488 7678 21540 7684
rect 23524 7606 23552 8222
rect 23708 8218 23736 9174
rect 23696 8212 23748 8218
rect 23696 8154 23748 8160
rect 23708 7946 23736 8154
rect 23696 7940 23748 7946
rect 23696 7882 23748 7888
rect 23892 7742 23920 10058
rect 24076 9986 24104 10262
rect 24064 9980 24116 9986
rect 24064 9922 24116 9928
rect 24628 9458 24656 11894
rect 24720 11686 24748 11962
rect 24708 11680 24760 11686
rect 24708 11622 24760 11628
rect 24720 11210 24748 11622
rect 24708 11204 24760 11210
rect 24708 11146 24760 11152
rect 24708 10456 24760 10462
rect 24708 10398 24760 10404
rect 24720 9850 24748 10398
rect 25258 10152 25314 10161
rect 25258 10087 25314 10096
rect 24708 9844 24760 9850
rect 24708 9786 24760 9792
rect 24720 9578 24748 9786
rect 24708 9572 24760 9578
rect 24708 9514 24760 9520
rect 25076 9504 25128 9510
rect 24156 9436 24208 9442
rect 24628 9430 24748 9458
rect 25076 9446 25128 9452
rect 24156 9378 24208 9384
rect 24168 8336 24196 9378
rect 24248 8348 24300 8354
rect 24168 8308 24248 8336
rect 24248 8290 24300 8296
rect 23972 8280 24024 8286
rect 23972 8222 24024 8228
rect 23984 7946 24012 8222
rect 23972 7940 24024 7946
rect 23972 7882 24024 7888
rect 23880 7736 23932 7742
rect 23880 7678 23932 7684
rect 23512 7600 23564 7606
rect 23512 7542 23564 7548
rect 21304 7396 21356 7402
rect 21304 7338 21356 7344
rect 21212 6784 21264 6790
rect 21212 6726 21264 6732
rect 20936 6648 20988 6654
rect 20936 6590 20988 6596
rect 20948 6314 20976 6590
rect 20936 6308 20988 6314
rect 20936 6250 20988 6256
rect 20476 5968 20528 5974
rect 20476 5910 20528 5916
rect 20488 5770 20516 5910
rect 20476 5764 20528 5770
rect 20476 5706 20528 5712
rect 20384 5628 20436 5634
rect 20384 5570 20436 5576
rect 19372 5560 19424 5566
rect 19372 5502 19424 5508
rect 19832 5560 19884 5566
rect 19832 5502 19884 5508
rect 18084 5152 18136 5158
rect 18820 5152 18872 5158
rect 18084 5094 18136 5100
rect 18740 5112 18820 5140
rect 17992 5016 18044 5022
rect 17992 4958 18044 4964
rect 17254 4576 17310 4585
rect 17254 4511 17310 4520
rect 17900 4472 17952 4478
rect 17900 4414 17952 4420
rect 17072 3928 17124 3934
rect 17072 3870 17124 3876
rect 17438 3760 17494 3769
rect 17438 3695 17494 3704
rect 15968 3520 16020 3526
rect 15968 3462 16020 3468
rect 15508 3316 15560 3322
rect 15508 3258 15560 3264
rect 14036 2908 14088 2914
rect 14036 2850 14088 2856
rect 14404 2908 14456 2914
rect 14404 2850 14456 2856
rect 15968 2908 16020 2914
rect 15968 2850 16020 2856
rect 14416 2506 14444 2850
rect 14956 2840 15008 2846
rect 14956 2782 15008 2788
rect 14968 2506 14996 2782
rect 15692 2704 15744 2710
rect 15692 2646 15744 2652
rect 14404 2500 14456 2506
rect 14404 2442 14456 2448
rect 14956 2500 15008 2506
rect 14956 2442 15008 2448
rect 13760 2432 13812 2438
rect 13760 2374 13812 2380
rect 13300 2296 13352 2302
rect 13300 2238 13352 2244
rect 15508 2228 15560 2234
rect 15508 2170 15560 2176
rect 13208 1956 13260 1962
rect 13208 1898 13260 1904
rect 15520 1894 15548 2170
rect 15704 1894 15732 2646
rect 15508 1888 15560 1894
rect 15508 1830 15560 1836
rect 15692 1888 15744 1894
rect 15692 1830 15744 1836
rect 12288 1820 12340 1826
rect 12288 1762 12340 1768
rect 13392 1820 13444 1826
rect 13392 1762 13444 1768
rect 14588 1820 14640 1826
rect 14588 1762 14640 1768
rect 15232 1820 15284 1826
rect 15232 1762 15284 1768
rect 12196 1412 12248 1418
rect 12196 1354 12248 1360
rect 11828 1344 11880 1350
rect 11828 1286 11880 1292
rect 12208 1214 12236 1354
rect 12300 1350 12328 1762
rect 13024 1752 13076 1758
rect 13024 1694 13076 1700
rect 13036 1350 13064 1694
rect 12288 1344 12340 1350
rect 12288 1286 12340 1292
rect 13024 1344 13076 1350
rect 13024 1286 13076 1292
rect 12196 1208 12248 1214
rect 12196 1150 12248 1156
rect 13404 1078 13432 1762
rect 13484 1752 13536 1758
rect 13484 1694 13536 1700
rect 14404 1752 14456 1758
rect 14404 1694 14456 1700
rect 13496 1418 13524 1694
rect 13484 1412 13536 1418
rect 13484 1354 13536 1360
rect 13392 1072 13444 1078
rect 13392 1014 13444 1020
rect 11644 596 11696 602
rect 11644 538 11696 544
rect 12380 596 12432 602
rect 12380 538 12432 544
rect 10000 420 10396 423
rect 12392 420 12420 538
rect 14416 420 14444 1694
rect 14600 1214 14628 1762
rect 14588 1208 14640 1214
rect 14588 1150 14640 1156
rect 15244 1146 15272 1762
rect 15232 1140 15284 1146
rect 15232 1082 15284 1088
rect 15520 874 15548 1830
rect 15704 1622 15732 1830
rect 15692 1616 15744 1622
rect 15692 1558 15744 1564
rect 15980 1350 16008 2850
rect 17452 2506 17480 3695
rect 17912 3390 17940 4414
rect 17900 3384 17952 3390
rect 17900 3326 17952 3332
rect 18004 3322 18032 4958
rect 18740 4682 18768 5112
rect 18820 5094 18872 5100
rect 19280 5152 19332 5158
rect 19280 5094 19332 5100
rect 18912 5084 18964 5090
rect 18912 5026 18964 5032
rect 18820 4948 18872 4954
rect 18820 4890 18872 4896
rect 18832 4682 18860 4890
rect 18728 4676 18780 4682
rect 18728 4618 18780 4624
rect 18820 4676 18872 4682
rect 18820 4618 18872 4624
rect 18832 4554 18860 4618
rect 18924 4614 18952 5026
rect 19384 4682 19412 5502
rect 19372 4676 19424 4682
rect 19372 4618 19424 4624
rect 19844 4614 19872 5502
rect 21224 5158 21252 6726
rect 21316 6722 21344 7338
rect 22040 7260 22092 7266
rect 22040 7202 22092 7208
rect 21672 7056 21724 7062
rect 21672 6998 21724 7004
rect 21304 6716 21356 6722
rect 21304 6658 21356 6664
rect 21684 6654 21712 6998
rect 22052 6858 22080 7202
rect 22040 6852 22092 6858
rect 22040 6794 22092 6800
rect 23524 6722 23552 7542
rect 23892 7402 23920 7678
rect 24260 7606 24288 8290
rect 24248 7600 24300 7606
rect 24248 7542 24300 7548
rect 23880 7396 23932 7402
rect 23880 7338 23932 7344
rect 23512 6716 23564 6722
rect 23512 6658 23564 6664
rect 21672 6648 21724 6654
rect 21672 6590 21724 6596
rect 21684 6246 21712 6590
rect 22316 6580 22368 6586
rect 22316 6522 22368 6528
rect 21672 6240 21724 6246
rect 21672 6182 21724 6188
rect 22328 5974 22356 6522
rect 22500 6172 22552 6178
rect 22500 6114 22552 6120
rect 22316 5968 22368 5974
rect 22316 5910 22368 5916
rect 22328 5770 22356 5910
rect 22316 5764 22368 5770
rect 22316 5706 22368 5712
rect 22512 5430 22540 6114
rect 22592 6104 22644 6110
rect 22592 6046 22644 6052
rect 23420 6104 23472 6110
rect 23420 6046 23472 6052
rect 21304 5424 21356 5430
rect 21304 5366 21356 5372
rect 21764 5424 21816 5430
rect 21764 5366 21816 5372
rect 22500 5424 22552 5430
rect 22500 5366 22552 5372
rect 21212 5152 21264 5158
rect 21212 5094 21264 5100
rect 21028 5016 21080 5022
rect 21028 4958 21080 4964
rect 21040 4614 21068 4958
rect 18740 4546 18860 4554
rect 18912 4608 18964 4614
rect 18912 4550 18964 4556
rect 19832 4608 19884 4614
rect 19832 4550 19884 4556
rect 21028 4608 21080 4614
rect 21028 4550 21080 4556
rect 21224 4554 21252 5094
rect 21316 4682 21344 5366
rect 21776 5158 21804 5366
rect 21764 5152 21816 5158
rect 21764 5094 21816 5100
rect 22512 5022 22540 5366
rect 22500 5016 22552 5022
rect 22500 4958 22552 4964
rect 22512 4682 22540 4958
rect 21304 4676 21356 4682
rect 21304 4618 21356 4624
rect 22500 4676 22552 4682
rect 22500 4618 22552 4624
rect 18728 4540 18860 4546
rect 18780 4526 18860 4540
rect 18728 4482 18780 4488
rect 18864 4236 19184 4256
rect 18864 4234 18876 4236
rect 18932 4234 18956 4236
rect 19012 4234 19036 4236
rect 19092 4234 19116 4236
rect 19172 4234 19184 4236
rect 18864 4182 18870 4234
rect 18932 4182 18934 4234
rect 19114 4182 19116 4234
rect 19178 4182 19184 4234
rect 18864 4180 18876 4182
rect 18932 4180 18956 4182
rect 19012 4180 19036 4182
rect 19092 4180 19116 4182
rect 19172 4180 19184 4182
rect 18864 4160 19184 4180
rect 18082 3896 18138 3905
rect 18082 3831 18138 3840
rect 17992 3316 18044 3322
rect 17992 3258 18044 3264
rect 18096 2982 18124 3831
rect 21040 3594 21068 4550
rect 21224 4546 21344 4554
rect 21224 4540 21356 4546
rect 21224 4526 21304 4540
rect 21304 4482 21356 4488
rect 22500 3792 22552 3798
rect 22500 3734 22552 3740
rect 22512 3594 22540 3734
rect 21028 3588 21080 3594
rect 22500 3588 22552 3594
rect 21080 3548 21160 3576
rect 21028 3530 21080 3536
rect 18864 3148 19184 3168
rect 18864 3146 18876 3148
rect 18932 3146 18956 3148
rect 19012 3146 19036 3148
rect 19092 3146 19116 3148
rect 19172 3146 19184 3148
rect 18864 3094 18870 3146
rect 18932 3094 18934 3146
rect 19114 3094 19116 3146
rect 19178 3094 19184 3146
rect 18864 3092 18876 3094
rect 18932 3092 18956 3094
rect 19012 3092 19036 3094
rect 19092 3092 19116 3094
rect 19172 3092 19184 3094
rect 18864 3072 19184 3092
rect 18084 2976 18136 2982
rect 18084 2918 18136 2924
rect 20936 2976 20988 2982
rect 20936 2918 20988 2924
rect 17992 2840 18044 2846
rect 17992 2782 18044 2788
rect 17440 2500 17492 2506
rect 17440 2442 17492 2448
rect 16520 2296 16572 2302
rect 16520 2238 16572 2244
rect 16532 1826 16560 2238
rect 17452 2234 17480 2442
rect 17900 2296 17952 2302
rect 17900 2238 17952 2244
rect 16704 2228 16756 2234
rect 16704 2170 16756 2176
rect 17440 2228 17492 2234
rect 17440 2170 17492 2176
rect 16716 1894 16744 2170
rect 16704 1888 16756 1894
rect 17912 1865 17940 2238
rect 18004 1962 18032 2782
rect 18096 2506 18124 2918
rect 18636 2908 18688 2914
rect 18636 2850 18688 2856
rect 18176 2840 18228 2846
rect 18176 2782 18228 2788
rect 18084 2500 18136 2506
rect 18084 2442 18136 2448
rect 18188 2234 18216 2782
rect 18648 2370 18676 2850
rect 20476 2840 20528 2846
rect 20476 2782 20528 2788
rect 18636 2364 18688 2370
rect 18636 2306 18688 2312
rect 18176 2228 18228 2234
rect 18176 2170 18228 2176
rect 17992 1956 18044 1962
rect 17992 1898 18044 1904
rect 18188 1894 18216 2170
rect 18176 1888 18228 1894
rect 16704 1830 16756 1836
rect 17898 1856 17954 1865
rect 16520 1820 16572 1826
rect 16520 1762 16572 1768
rect 16336 1616 16388 1622
rect 16336 1558 16388 1564
rect 16348 1418 16376 1558
rect 16336 1412 16388 1418
rect 16532 1400 16560 1762
rect 16612 1412 16664 1418
rect 16532 1372 16612 1400
rect 16336 1354 16388 1360
rect 16612 1354 16664 1360
rect 15968 1344 16020 1350
rect 15968 1286 16020 1292
rect 16428 1208 16480 1214
rect 16428 1150 16480 1156
rect 15508 868 15560 874
rect 15508 810 15560 816
rect 16440 806 16468 1150
rect 16716 1146 16744 1830
rect 17898 1791 17954 1800
rect 18082 1856 18138 1865
rect 18176 1830 18228 1836
rect 18082 1791 18138 1800
rect 18648 1808 18676 2306
rect 19556 2296 19608 2302
rect 19556 2238 19608 2244
rect 19280 2228 19332 2234
rect 19280 2170 19332 2176
rect 18864 2060 19184 2080
rect 18864 2058 18876 2060
rect 18932 2058 18956 2060
rect 19012 2058 19036 2060
rect 19092 2058 19116 2060
rect 19172 2058 19184 2060
rect 18864 2006 18870 2058
rect 18932 2006 18934 2058
rect 19114 2006 19116 2058
rect 19178 2006 19184 2058
rect 18864 2004 18876 2006
rect 18932 2004 18956 2006
rect 19012 2004 19036 2006
rect 19092 2004 19116 2006
rect 19172 2004 19184 2006
rect 18864 1984 19184 2004
rect 18912 1820 18964 1826
rect 18096 1758 18124 1791
rect 18648 1780 18912 1808
rect 18912 1762 18964 1768
rect 18084 1752 18136 1758
rect 18084 1694 18136 1700
rect 17900 1616 17952 1622
rect 17900 1558 17952 1564
rect 16704 1140 16756 1146
rect 16704 1082 16756 1088
rect 17912 1078 17940 1558
rect 18452 1276 18504 1282
rect 18452 1218 18504 1224
rect 17900 1072 17952 1078
rect 17900 1014 17952 1020
rect 16428 800 16480 806
rect 16428 742 16480 748
rect 16440 420 16468 742
rect 18464 420 18492 1218
rect 18634 1176 18690 1185
rect 18924 1146 18952 1762
rect 19004 1752 19056 1758
rect 19004 1694 19056 1700
rect 19016 1418 19044 1694
rect 19004 1412 19056 1418
rect 19004 1354 19056 1360
rect 19292 1185 19320 2170
rect 19568 1962 19596 2238
rect 19556 1956 19608 1962
rect 19556 1898 19608 1904
rect 19464 1888 19516 1894
rect 19464 1830 19516 1836
rect 19476 1350 19504 1830
rect 20488 1758 20516 2782
rect 20752 2772 20804 2778
rect 20752 2714 20804 2720
rect 20764 2370 20792 2714
rect 20752 2364 20804 2370
rect 20752 2306 20804 2312
rect 20764 1962 20792 2306
rect 20948 2166 20976 2918
rect 21132 2370 21160 3548
rect 22500 3530 22552 3536
rect 22132 2908 22184 2914
rect 22132 2850 22184 2856
rect 22408 2908 22460 2914
rect 22408 2850 22460 2856
rect 22144 2506 22172 2850
rect 22420 2710 22448 2850
rect 22512 2846 22540 3530
rect 22500 2840 22552 2846
rect 22500 2782 22552 2788
rect 22408 2704 22460 2710
rect 22408 2646 22460 2652
rect 22132 2500 22184 2506
rect 22132 2442 22184 2448
rect 21120 2364 21172 2370
rect 21120 2306 21172 2312
rect 21028 2296 21080 2302
rect 21028 2238 21080 2244
rect 20936 2160 20988 2166
rect 20936 2102 20988 2108
rect 20752 1956 20804 1962
rect 20752 1898 20804 1904
rect 20844 1820 20896 1826
rect 20844 1762 20896 1768
rect 20476 1752 20528 1758
rect 20476 1694 20528 1700
rect 20856 1418 20884 1762
rect 20844 1412 20896 1418
rect 20844 1354 20896 1360
rect 19464 1344 19516 1350
rect 19464 1286 19516 1292
rect 20948 1282 20976 2102
rect 21040 1418 21068 2238
rect 22144 1962 22172 2442
rect 22420 2438 22448 2646
rect 22512 2506 22540 2782
rect 22500 2500 22552 2506
rect 22500 2442 22552 2448
rect 22408 2432 22460 2438
rect 22604 2386 22632 6046
rect 23432 5770 23460 6046
rect 23788 5968 23840 5974
rect 23788 5910 23840 5916
rect 23420 5764 23472 5770
rect 23420 5706 23472 5712
rect 23800 5702 23828 5910
rect 23788 5696 23840 5702
rect 23788 5638 23840 5644
rect 23892 5634 23920 7338
rect 24260 6178 24288 7542
rect 24616 6512 24668 6518
rect 24616 6454 24668 6460
rect 24628 6178 24656 6454
rect 24248 6172 24300 6178
rect 24248 6114 24300 6120
rect 24616 6172 24668 6178
rect 24616 6114 24668 6120
rect 24156 5968 24208 5974
rect 24156 5910 24208 5916
rect 24168 5634 24196 5910
rect 24260 5770 24288 6114
rect 24616 6036 24668 6042
rect 24616 5978 24668 5984
rect 24248 5764 24300 5770
rect 24248 5706 24300 5712
rect 23880 5628 23932 5634
rect 23880 5570 23932 5576
rect 24156 5628 24208 5634
rect 24156 5570 24208 5576
rect 23892 5226 23920 5570
rect 24168 5226 24196 5570
rect 24628 5498 24656 5978
rect 24616 5492 24668 5498
rect 24616 5434 24668 5440
rect 24432 5424 24484 5430
rect 24432 5366 24484 5372
rect 23880 5220 23932 5226
rect 23880 5162 23932 5168
rect 24156 5220 24208 5226
rect 24156 5162 24208 5168
rect 23892 4614 23920 5162
rect 24444 5090 24472 5366
rect 24628 5158 24656 5434
rect 24616 5152 24668 5158
rect 24616 5094 24668 5100
rect 24432 5084 24484 5090
rect 24432 5026 24484 5032
rect 24444 4682 24472 5026
rect 24628 4682 24656 5094
rect 24432 4676 24484 4682
rect 24432 4618 24484 4624
rect 24616 4676 24668 4682
rect 24616 4618 24668 4624
rect 23880 4608 23932 4614
rect 23880 4550 23932 4556
rect 23604 4132 23656 4138
rect 23604 4074 23656 4080
rect 22684 4064 22736 4070
rect 22684 4006 22736 4012
rect 22696 3254 22724 4006
rect 22776 3996 22828 4002
rect 22776 3938 22828 3944
rect 22788 3594 22816 3938
rect 22776 3588 22828 3594
rect 22776 3530 22828 3536
rect 23616 3390 23644 4074
rect 23880 3792 23932 3798
rect 23880 3734 23932 3740
rect 24340 3792 24392 3798
rect 24340 3734 24392 3740
rect 23892 3594 23920 3734
rect 23880 3588 23932 3594
rect 23880 3530 23932 3536
rect 23880 3452 23932 3458
rect 23880 3394 23932 3400
rect 23604 3384 23656 3390
rect 23604 3326 23656 3332
rect 22684 3248 22736 3254
rect 22684 3190 22736 3196
rect 23512 3248 23564 3254
rect 23512 3190 23564 3196
rect 22696 3050 22724 3190
rect 22684 3044 22736 3050
rect 22684 2986 22736 2992
rect 23524 2914 23552 3190
rect 23512 2908 23564 2914
rect 23512 2850 23564 2856
rect 22408 2374 22460 2380
rect 22512 2358 22632 2386
rect 22132 1956 22184 1962
rect 22132 1898 22184 1904
rect 21764 1752 21816 1758
rect 21764 1694 21816 1700
rect 21028 1412 21080 1418
rect 21028 1354 21080 1360
rect 21776 1350 21804 1694
rect 21764 1344 21816 1350
rect 21764 1286 21816 1292
rect 20936 1276 20988 1282
rect 20936 1218 20988 1224
rect 19278 1176 19334 1185
rect 18634 1111 18690 1120
rect 18912 1140 18964 1146
rect 18648 1078 18676 1111
rect 19278 1111 19334 1120
rect 20476 1140 20528 1146
rect 18912 1082 18964 1088
rect 20476 1082 20528 1088
rect 18636 1072 18688 1078
rect 18636 1014 18688 1020
rect 18864 972 19184 992
rect 18864 970 18876 972
rect 18932 970 18956 972
rect 19012 970 19036 972
rect 19092 970 19116 972
rect 19172 970 19184 972
rect 18864 918 18870 970
rect 18932 918 18934 970
rect 19114 918 19116 970
rect 19178 918 19184 970
rect 18864 916 18876 918
rect 18932 916 18956 918
rect 19012 916 19036 918
rect 19092 916 19116 918
rect 19172 916 19184 918
rect 18864 896 19184 916
rect 20488 420 20516 1082
rect 22512 420 22540 2358
rect 23524 2166 23552 2850
rect 23616 2506 23644 3326
rect 23892 2914 23920 3394
rect 24352 3322 24380 3734
rect 24340 3316 24392 3322
rect 24340 3258 24392 3264
rect 24156 3044 24208 3050
rect 24156 2986 24208 2992
rect 23880 2908 23932 2914
rect 23880 2850 23932 2856
rect 23604 2500 23656 2506
rect 23604 2442 23656 2448
rect 23420 2160 23472 2166
rect 23420 2102 23472 2108
rect 23512 2160 23564 2166
rect 23512 2102 23564 2108
rect 23432 2001 23460 2102
rect 23418 1992 23474 2001
rect 23052 1956 23104 1962
rect 23418 1927 23474 1936
rect 23052 1898 23104 1904
rect 23064 1418 23092 1898
rect 23236 1888 23288 1894
rect 23236 1830 23288 1836
rect 23248 1418 23276 1830
rect 23432 1826 23460 1927
rect 23524 1865 23552 2102
rect 23616 1894 23644 2442
rect 23892 2234 23920 2850
rect 24064 2704 24116 2710
rect 24064 2646 24116 2652
rect 23880 2228 23932 2234
rect 23880 2170 23932 2176
rect 23892 1962 23920 2170
rect 24076 1962 24104 2646
rect 24168 2370 24196 2986
rect 24156 2364 24208 2370
rect 24156 2306 24208 2312
rect 23880 1956 23932 1962
rect 23880 1898 23932 1904
rect 24064 1956 24116 1962
rect 24064 1898 24116 1904
rect 24168 1894 24196 2306
rect 24352 2234 24380 3258
rect 24432 2704 24484 2710
rect 24432 2646 24484 2652
rect 24444 2506 24472 2646
rect 24432 2500 24484 2506
rect 24432 2442 24484 2448
rect 24340 2228 24392 2234
rect 24340 2170 24392 2176
rect 24352 1962 24380 2170
rect 24720 1962 24748 9430
rect 24892 7668 24944 7674
rect 24892 7610 24944 7616
rect 24904 7334 24932 7610
rect 24892 7328 24944 7334
rect 24892 7270 24944 7276
rect 24904 6722 24932 7270
rect 24892 6716 24944 6722
rect 24892 6658 24944 6664
rect 25088 6654 25116 9446
rect 25168 9368 25220 9374
rect 25168 9310 25220 9316
rect 25180 8898 25208 9310
rect 25168 8892 25220 8898
rect 25168 8834 25220 8840
rect 25076 6648 25128 6654
rect 25076 6590 25128 6596
rect 25088 5430 25116 6590
rect 25076 5424 25128 5430
rect 25076 5366 25128 5372
rect 25272 3050 25300 10087
rect 25364 4138 25392 25047
rect 25456 19273 25484 27262
rect 26376 27228 26404 27262
rect 25812 19636 25864 19642
rect 25812 19578 25864 19584
rect 25442 19264 25498 19273
rect 25442 19199 25498 19208
rect 25824 17738 25852 19578
rect 26178 19400 26234 19409
rect 26178 19335 26234 19344
rect 26192 19302 26220 19335
rect 26180 19296 26232 19302
rect 26180 19238 26232 19244
rect 26088 19024 26140 19030
rect 26088 18966 26140 18972
rect 25996 18480 26048 18486
rect 26100 18468 26128 18966
rect 26192 18826 26220 19238
rect 26180 18820 26232 18826
rect 26180 18762 26232 18768
rect 26180 18480 26232 18486
rect 26100 18440 26180 18468
rect 25996 18422 26048 18428
rect 26180 18422 26232 18428
rect 25812 17732 25864 17738
rect 25812 17674 25864 17680
rect 25824 16514 25852 17674
rect 25812 16508 25864 16514
rect 25732 16468 25812 16496
rect 25732 16106 25760 16468
rect 25812 16450 25864 16456
rect 25812 16372 25864 16378
rect 25812 16314 25864 16320
rect 25720 16100 25772 16106
rect 25720 16042 25772 16048
rect 25824 15970 25852 16314
rect 25812 15964 25864 15970
rect 25812 15906 25864 15912
rect 25824 15426 25852 15906
rect 25812 15420 25864 15426
rect 25812 15362 25864 15368
rect 25824 14950 25852 15362
rect 25812 14944 25864 14950
rect 25812 14886 25864 14892
rect 26008 14270 26036 18422
rect 26192 18185 26220 18422
rect 26178 18176 26234 18185
rect 26178 18111 26234 18120
rect 26456 17052 26508 17058
rect 26456 16994 26508 17000
rect 26364 16848 26416 16854
rect 26364 16790 26416 16796
rect 26376 16689 26404 16790
rect 26362 16680 26418 16689
rect 26468 16650 26496 16994
rect 26362 16615 26418 16624
rect 26456 16644 26508 16650
rect 26376 16582 26404 16615
rect 26456 16586 26508 16592
rect 26364 16576 26416 16582
rect 26364 16518 26416 16524
rect 26272 16372 26324 16378
rect 26272 16314 26324 16320
rect 26284 15766 26312 16314
rect 26272 15760 26324 15766
rect 26272 15702 26324 15708
rect 26284 15562 26312 15702
rect 26272 15556 26324 15562
rect 26272 15498 26324 15504
rect 25996 14264 26048 14270
rect 25996 14206 26048 14212
rect 25720 13040 25772 13046
rect 25720 12982 25772 12988
rect 25732 12026 25760 12982
rect 25720 12020 25772 12026
rect 25720 11962 25772 11968
rect 25732 11754 25760 11962
rect 25720 11748 25772 11754
rect 25720 11690 25772 11696
rect 25444 9980 25496 9986
rect 25444 9922 25496 9928
rect 25456 9034 25484 9922
rect 25444 9028 25496 9034
rect 25444 8970 25496 8976
rect 25456 8830 25484 8970
rect 25444 8824 25496 8830
rect 25444 8766 25496 8772
rect 26180 8348 26232 8354
rect 26180 8290 26232 8296
rect 26192 7674 26220 8290
rect 26272 8144 26324 8150
rect 26272 8086 26324 8092
rect 26284 7946 26312 8086
rect 26272 7940 26324 7946
rect 26272 7882 26324 7888
rect 26180 7668 26232 7674
rect 26180 7610 26232 7616
rect 26192 7402 26220 7610
rect 26180 7396 26232 7402
rect 26180 7338 26232 7344
rect 25904 6172 25956 6178
rect 25904 6114 25956 6120
rect 25916 5634 25944 6114
rect 25904 5628 25956 5634
rect 25904 5570 25956 5576
rect 25352 4132 25404 4138
rect 25352 4074 25404 4080
rect 25260 3044 25312 3050
rect 25260 2986 25312 2992
rect 24892 2228 24944 2234
rect 24892 2170 24944 2176
rect 24340 1956 24392 1962
rect 24340 1898 24392 1904
rect 24708 1956 24760 1962
rect 24708 1898 24760 1904
rect 23604 1888 23656 1894
rect 23510 1856 23566 1865
rect 23420 1820 23472 1826
rect 23604 1830 23656 1836
rect 24156 1888 24208 1894
rect 24156 1830 24208 1836
rect 23510 1791 23566 1800
rect 23420 1762 23472 1768
rect 23432 1418 23460 1762
rect 24168 1418 24196 1830
rect 23052 1412 23104 1418
rect 23052 1354 23104 1360
rect 23236 1412 23288 1418
rect 23236 1354 23288 1360
rect 23420 1412 23472 1418
rect 23420 1354 23472 1360
rect 24156 1412 24208 1418
rect 24156 1354 24208 1360
rect 24904 1185 24932 2170
rect 26364 1956 26416 1962
rect 26364 1898 26416 1904
rect 26272 1820 26324 1826
rect 26272 1762 26324 1768
rect 25628 1208 25680 1214
rect 24890 1176 24946 1185
rect 25628 1150 25680 1156
rect 24890 1111 24892 1120
rect 24944 1111 24946 1120
rect 24892 1082 24944 1088
rect 24524 1072 24576 1078
rect 24524 1014 24576 1020
rect 24536 420 24564 1014
rect 24904 806 24932 1082
rect 25640 874 25668 1150
rect 26284 1078 26312 1762
rect 26376 1418 26404 1898
rect 26364 1412 26416 1418
rect 26364 1354 26416 1360
rect 26272 1072 26324 1078
rect 26272 1014 26324 1020
rect 25628 868 25680 874
rect 25628 810 25680 816
rect 24892 800 24944 806
rect 24892 742 24944 748
rect 26284 423 26312 1014
rect 26284 420 26588 423
rect 3504 372 3516 374
rect 3572 372 3596 374
rect 3652 372 3676 374
rect 3732 372 3756 374
rect 3812 372 3824 374
rect 3504 352 3824 372
rect 4240 0 4380 420
rect 6264 0 6404 420
rect 8288 0 8428 420
rect 10000 395 10452 420
rect 10312 0 10452 395
rect 12336 0 12476 420
rect 14360 0 14500 420
rect 16384 0 16524 420
rect 18408 0 18548 420
rect 20432 0 20572 420
rect 22456 0 22596 420
rect 24480 0 24620 420
rect 26284 395 26644 420
rect 26504 0 26644 395
<< via2 >>
rect 878 26960 934 27016
rect 878 20976 934 21032
rect 1430 23968 1486 24024
rect 878 17984 934 18040
rect 878 14992 934 15048
rect 694 12000 750 12056
rect 694 9008 750 9064
rect 878 6016 934 6072
rect 3516 26538 3572 26540
rect 3596 26538 3652 26540
rect 3676 26538 3732 26540
rect 3756 26538 3812 26540
rect 3516 26486 3562 26538
rect 3562 26486 3572 26538
rect 3596 26486 3626 26538
rect 3626 26486 3638 26538
rect 3638 26486 3652 26538
rect 3676 26486 3690 26538
rect 3690 26486 3702 26538
rect 3702 26486 3732 26538
rect 3756 26486 3766 26538
rect 3766 26486 3812 26538
rect 3516 26484 3572 26486
rect 3596 26484 3652 26486
rect 3676 26484 3732 26486
rect 3756 26484 3812 26486
rect 3516 25450 3572 25452
rect 3596 25450 3652 25452
rect 3676 25450 3732 25452
rect 3756 25450 3812 25452
rect 3516 25398 3562 25450
rect 3562 25398 3572 25450
rect 3596 25398 3626 25450
rect 3626 25398 3638 25450
rect 3638 25398 3652 25450
rect 3676 25398 3690 25450
rect 3690 25398 3702 25450
rect 3702 25398 3732 25450
rect 3756 25398 3766 25450
rect 3766 25398 3812 25450
rect 3516 25396 3572 25398
rect 3596 25396 3652 25398
rect 3676 25396 3732 25398
rect 3756 25396 3812 25398
rect 3516 24362 3572 24364
rect 3596 24362 3652 24364
rect 3676 24362 3732 24364
rect 3756 24362 3812 24364
rect 3516 24310 3562 24362
rect 3562 24310 3572 24362
rect 3596 24310 3626 24362
rect 3626 24310 3638 24362
rect 3638 24310 3652 24362
rect 3676 24310 3690 24362
rect 3690 24310 3702 24362
rect 3702 24310 3732 24362
rect 3756 24310 3766 24362
rect 3766 24310 3812 24362
rect 3516 24308 3572 24310
rect 3596 24308 3652 24310
rect 3676 24308 3732 24310
rect 3756 24308 3812 24310
rect 3516 23274 3572 23276
rect 3596 23274 3652 23276
rect 3676 23274 3732 23276
rect 3756 23274 3812 23276
rect 3516 23222 3562 23274
rect 3562 23222 3572 23274
rect 3596 23222 3626 23274
rect 3626 23222 3638 23274
rect 3638 23222 3652 23274
rect 3676 23222 3690 23274
rect 3690 23222 3702 23274
rect 3702 23222 3732 23274
rect 3756 23222 3766 23274
rect 3766 23222 3812 23274
rect 3516 23220 3572 23222
rect 3596 23220 3652 23222
rect 3676 23220 3732 23222
rect 3756 23220 3812 23222
rect 3516 22186 3572 22188
rect 3596 22186 3652 22188
rect 3676 22186 3732 22188
rect 3756 22186 3812 22188
rect 3516 22134 3562 22186
rect 3562 22134 3572 22186
rect 3596 22134 3626 22186
rect 3626 22134 3638 22186
rect 3638 22134 3652 22186
rect 3676 22134 3690 22186
rect 3690 22134 3702 22186
rect 3702 22134 3732 22186
rect 3756 22134 3766 22186
rect 3766 22134 3812 22186
rect 3516 22132 3572 22134
rect 3596 22132 3652 22134
rect 3676 22132 3732 22134
rect 3756 22132 3812 22134
rect 3516 21098 3572 21100
rect 3596 21098 3652 21100
rect 3676 21098 3732 21100
rect 3756 21098 3812 21100
rect 3516 21046 3562 21098
rect 3562 21046 3572 21098
rect 3596 21046 3626 21098
rect 3626 21046 3638 21098
rect 3638 21046 3652 21098
rect 3676 21046 3690 21098
rect 3690 21046 3702 21098
rect 3702 21046 3732 21098
rect 3756 21046 3766 21098
rect 3766 21046 3812 21098
rect 3516 21044 3572 21046
rect 3596 21044 3652 21046
rect 3676 21044 3732 21046
rect 3756 21044 3812 21046
rect 3516 20010 3572 20012
rect 3596 20010 3652 20012
rect 3676 20010 3732 20012
rect 3756 20010 3812 20012
rect 3516 19958 3562 20010
rect 3562 19958 3572 20010
rect 3596 19958 3626 20010
rect 3626 19958 3638 20010
rect 3638 19958 3652 20010
rect 3676 19958 3690 20010
rect 3690 19958 3702 20010
rect 3702 19958 3732 20010
rect 3756 19958 3766 20010
rect 3766 19958 3812 20010
rect 3516 19956 3572 19958
rect 3596 19956 3652 19958
rect 3676 19956 3732 19958
rect 3756 19956 3812 19958
rect 1982 15400 2038 15456
rect 1706 15128 1762 15184
rect 3516 18922 3572 18924
rect 3596 18922 3652 18924
rect 3676 18922 3732 18924
rect 3756 18922 3812 18924
rect 3516 18870 3562 18922
rect 3562 18870 3572 18922
rect 3596 18870 3626 18922
rect 3626 18870 3638 18922
rect 3638 18870 3652 18922
rect 3676 18870 3690 18922
rect 3690 18870 3702 18922
rect 3702 18870 3732 18922
rect 3756 18870 3766 18922
rect 3766 18870 3812 18922
rect 3516 18868 3572 18870
rect 3596 18868 3652 18870
rect 3676 18868 3732 18870
rect 3756 18868 3812 18870
rect 2350 17576 2406 17632
rect 3516 17834 3572 17836
rect 3596 17834 3652 17836
rect 3676 17834 3732 17836
rect 3756 17834 3812 17836
rect 3516 17782 3562 17834
rect 3562 17782 3572 17834
rect 3596 17782 3626 17834
rect 3626 17782 3638 17834
rect 3638 17782 3652 17834
rect 3676 17782 3690 17834
rect 3690 17782 3702 17834
rect 3702 17782 3732 17834
rect 3756 17782 3766 17834
rect 3766 17782 3812 17834
rect 3516 17780 3572 17782
rect 3596 17780 3652 17782
rect 3676 17780 3732 17782
rect 3756 17780 3812 17782
rect 3516 16746 3572 16748
rect 3596 16746 3652 16748
rect 3676 16746 3732 16748
rect 3756 16746 3812 16748
rect 3516 16694 3562 16746
rect 3562 16694 3572 16746
rect 3596 16694 3626 16746
rect 3626 16694 3638 16746
rect 3638 16694 3652 16746
rect 3676 16694 3690 16746
rect 3690 16694 3702 16746
rect 3702 16694 3732 16746
rect 3756 16694 3766 16746
rect 3766 16694 3812 16746
rect 3516 16692 3572 16694
rect 3596 16692 3652 16694
rect 3676 16692 3732 16694
rect 3756 16692 3812 16694
rect 1430 3840 1486 3896
rect 418 3024 474 3080
rect 418 1800 474 1856
rect 2994 15400 3050 15456
rect 3516 15658 3572 15660
rect 3596 15658 3652 15660
rect 3676 15658 3732 15660
rect 3756 15658 3812 15660
rect 3516 15606 3562 15658
rect 3562 15606 3572 15658
rect 3596 15606 3626 15658
rect 3626 15606 3638 15658
rect 3638 15606 3652 15658
rect 3676 15606 3690 15658
rect 3690 15606 3702 15658
rect 3702 15606 3732 15658
rect 3756 15606 3766 15658
rect 3766 15606 3812 15658
rect 3516 15604 3572 15606
rect 3596 15604 3652 15606
rect 3676 15604 3732 15606
rect 3756 15604 3812 15606
rect 3516 14570 3572 14572
rect 3596 14570 3652 14572
rect 3676 14570 3732 14572
rect 3756 14570 3812 14572
rect 3516 14518 3562 14570
rect 3562 14518 3572 14570
rect 3596 14518 3626 14570
rect 3626 14518 3638 14570
rect 3638 14518 3652 14570
rect 3676 14518 3690 14570
rect 3690 14518 3702 14570
rect 3702 14518 3732 14570
rect 3756 14518 3766 14570
rect 3766 14518 3812 14570
rect 3516 14516 3572 14518
rect 3596 14516 3652 14518
rect 3676 14516 3732 14518
rect 3756 14516 3812 14518
rect 3270 14176 3326 14232
rect 3516 13482 3572 13484
rect 3596 13482 3652 13484
rect 3676 13482 3732 13484
rect 3756 13482 3812 13484
rect 3516 13430 3562 13482
rect 3562 13430 3572 13482
rect 3596 13430 3626 13482
rect 3626 13430 3638 13482
rect 3638 13430 3652 13482
rect 3676 13430 3690 13482
rect 3690 13430 3702 13482
rect 3702 13430 3732 13482
rect 3756 13430 3766 13482
rect 3766 13430 3812 13482
rect 3516 13428 3572 13430
rect 3596 13428 3652 13430
rect 3676 13428 3732 13430
rect 3756 13428 3812 13430
rect 4926 14584 4982 14640
rect 5202 14584 5258 14640
rect 4282 14176 4338 14232
rect 3516 12394 3572 12396
rect 3596 12394 3652 12396
rect 3676 12394 3732 12396
rect 3756 12394 3812 12396
rect 3516 12342 3562 12394
rect 3562 12342 3572 12394
rect 3596 12342 3626 12394
rect 3626 12342 3638 12394
rect 3638 12342 3652 12394
rect 3676 12342 3690 12394
rect 3690 12342 3702 12394
rect 3702 12342 3732 12394
rect 3756 12342 3766 12394
rect 3766 12342 3812 12394
rect 3516 12340 3572 12342
rect 3596 12340 3652 12342
rect 3676 12340 3732 12342
rect 3756 12340 3812 12342
rect 3516 11306 3572 11308
rect 3596 11306 3652 11308
rect 3676 11306 3732 11308
rect 3756 11306 3812 11308
rect 3516 11254 3562 11306
rect 3562 11254 3572 11306
rect 3596 11254 3626 11306
rect 3626 11254 3638 11306
rect 3638 11254 3652 11306
rect 3676 11254 3690 11306
rect 3690 11254 3702 11306
rect 3702 11254 3732 11306
rect 3756 11254 3766 11306
rect 3766 11254 3812 11306
rect 3516 11252 3572 11254
rect 3596 11252 3652 11254
rect 3676 11252 3732 11254
rect 3756 11252 3812 11254
rect 3516 10218 3572 10220
rect 3596 10218 3652 10220
rect 3676 10218 3732 10220
rect 3756 10218 3812 10220
rect 3516 10166 3562 10218
rect 3562 10166 3572 10218
rect 3596 10166 3626 10218
rect 3626 10166 3638 10218
rect 3638 10166 3652 10218
rect 3676 10166 3690 10218
rect 3690 10166 3702 10218
rect 3702 10166 3732 10218
rect 3756 10166 3766 10218
rect 3766 10166 3812 10218
rect 3516 10164 3572 10166
rect 3596 10164 3652 10166
rect 3676 10164 3732 10166
rect 3756 10164 3812 10166
rect 3516 9130 3572 9132
rect 3596 9130 3652 9132
rect 3676 9130 3732 9132
rect 3756 9130 3812 9132
rect 3516 9078 3562 9130
rect 3562 9078 3572 9130
rect 3596 9078 3626 9130
rect 3626 9078 3638 9130
rect 3638 9078 3652 9130
rect 3676 9078 3690 9130
rect 3690 9078 3702 9130
rect 3702 9078 3732 9130
rect 3756 9078 3766 9130
rect 3766 9078 3812 9130
rect 3516 9076 3572 9078
rect 3596 9076 3652 9078
rect 3676 9076 3732 9078
rect 3756 9076 3812 9078
rect 5662 12952 5718 13008
rect 3516 8042 3572 8044
rect 3596 8042 3652 8044
rect 3676 8042 3732 8044
rect 3756 8042 3812 8044
rect 3516 7990 3562 8042
rect 3562 7990 3572 8042
rect 3596 7990 3626 8042
rect 3626 7990 3638 8042
rect 3638 7990 3652 8042
rect 3676 7990 3690 8042
rect 3690 7990 3702 8042
rect 3702 7990 3732 8042
rect 3756 7990 3766 8042
rect 3766 7990 3812 8042
rect 3516 7988 3572 7990
rect 3596 7988 3652 7990
rect 3676 7988 3732 7990
rect 3756 7988 3812 7990
rect 3516 6954 3572 6956
rect 3596 6954 3652 6956
rect 3676 6954 3732 6956
rect 3756 6954 3812 6956
rect 3516 6902 3562 6954
rect 3562 6902 3572 6954
rect 3596 6902 3626 6954
rect 3626 6902 3638 6954
rect 3638 6902 3652 6954
rect 3676 6902 3690 6954
rect 3690 6902 3702 6954
rect 3702 6902 3732 6954
rect 3756 6902 3766 6954
rect 3766 6902 3812 6954
rect 3516 6900 3572 6902
rect 3596 6900 3652 6902
rect 3676 6900 3732 6902
rect 3756 6900 3812 6902
rect 6490 24648 6546 24704
rect 6674 14040 6730 14096
rect 6858 12952 6914 13008
rect 3516 5866 3572 5868
rect 3596 5866 3652 5868
rect 3676 5866 3732 5868
rect 3756 5866 3812 5868
rect 3516 5814 3562 5866
rect 3562 5814 3572 5866
rect 3596 5814 3626 5866
rect 3626 5814 3638 5866
rect 3638 5814 3652 5866
rect 3676 5814 3690 5866
rect 3690 5814 3702 5866
rect 3702 5814 3732 5866
rect 3756 5814 3766 5866
rect 3766 5814 3812 5866
rect 3516 5812 3572 5814
rect 3596 5812 3652 5814
rect 3676 5812 3732 5814
rect 3756 5812 3812 5814
rect 3516 4778 3572 4780
rect 3596 4778 3652 4780
rect 3676 4778 3732 4780
rect 3756 4778 3812 4780
rect 3516 4726 3562 4778
rect 3562 4726 3572 4778
rect 3596 4726 3626 4778
rect 3626 4726 3638 4778
rect 3638 4726 3652 4778
rect 3676 4726 3690 4778
rect 3690 4726 3702 4778
rect 3702 4726 3732 4778
rect 3756 4726 3766 4778
rect 3766 4726 3812 4778
rect 3516 4724 3572 4726
rect 3596 4724 3652 4726
rect 3676 4724 3732 4726
rect 3756 4724 3812 4726
rect 3516 3690 3572 3692
rect 3596 3690 3652 3692
rect 3676 3690 3732 3692
rect 3756 3690 3812 3692
rect 3516 3638 3562 3690
rect 3562 3638 3572 3690
rect 3596 3638 3626 3690
rect 3626 3638 3638 3690
rect 3638 3638 3652 3690
rect 3676 3638 3690 3690
rect 3690 3638 3702 3690
rect 3702 3638 3732 3690
rect 3756 3638 3766 3690
rect 3766 3638 3812 3690
rect 3516 3636 3572 3638
rect 3596 3636 3652 3638
rect 3676 3636 3732 3638
rect 3756 3636 3812 3638
rect 3516 2602 3572 2604
rect 3596 2602 3652 2604
rect 3676 2602 3732 2604
rect 3756 2602 3812 2604
rect 3516 2550 3562 2602
rect 3562 2550 3572 2602
rect 3596 2550 3626 2602
rect 3626 2550 3638 2602
rect 3638 2550 3652 2602
rect 3676 2550 3690 2602
rect 3690 2550 3702 2602
rect 3702 2550 3732 2602
rect 3756 2550 3766 2602
rect 3766 2550 3812 2602
rect 3516 2548 3572 2550
rect 3596 2548 3652 2550
rect 3676 2548 3732 2550
rect 3756 2548 3812 2550
rect 3516 1514 3572 1516
rect 3596 1514 3652 1516
rect 3676 1514 3732 1516
rect 3756 1514 3812 1516
rect 3516 1462 3562 1514
rect 3562 1462 3572 1514
rect 3596 1462 3626 1514
rect 3626 1462 3638 1514
rect 3638 1462 3652 1514
rect 3676 1462 3690 1514
rect 3690 1462 3702 1514
rect 3702 1462 3732 1514
rect 3756 1462 3766 1514
rect 3766 1462 3812 1514
rect 3516 1460 3572 1462
rect 3596 1460 3652 1462
rect 3676 1460 3732 1462
rect 3756 1460 3812 1462
rect 3516 426 3572 428
rect 3596 426 3652 428
rect 3676 426 3732 428
rect 3756 426 3812 428
rect 3516 374 3562 426
rect 3562 374 3572 426
rect 3596 374 3626 426
rect 3626 374 3638 426
rect 3638 374 3652 426
rect 3676 374 3690 426
rect 3690 374 3702 426
rect 3702 374 3732 426
rect 3756 374 3766 426
rect 3766 374 3812 426
rect 7134 12680 7190 12736
rect 7870 15128 7926 15184
rect 8238 12680 8294 12736
rect 9986 18120 10042 18176
rect 9526 13904 9582 13960
rect 7042 3704 7098 3760
rect 10170 14040 10226 14096
rect 10630 14176 10686 14232
rect 10630 14040 10686 14096
rect 12194 14176 12250 14232
rect 13574 19208 13630 19264
rect 12378 17712 12434 17768
rect 12838 14040 12894 14096
rect 15138 17576 15194 17632
rect 18876 27082 18932 27084
rect 18956 27082 19012 27084
rect 19036 27082 19092 27084
rect 19116 27082 19172 27084
rect 18876 27030 18922 27082
rect 18922 27030 18932 27082
rect 18956 27030 18986 27082
rect 18986 27030 18998 27082
rect 18998 27030 19012 27082
rect 19036 27030 19050 27082
rect 19050 27030 19062 27082
rect 19062 27030 19092 27082
rect 19116 27030 19126 27082
rect 19126 27030 19172 27082
rect 18876 27028 18932 27030
rect 18956 27028 19012 27030
rect 19036 27028 19092 27030
rect 19116 27028 19172 27030
rect 18876 25994 18932 25996
rect 18956 25994 19012 25996
rect 19036 25994 19092 25996
rect 19116 25994 19172 25996
rect 18876 25942 18922 25994
rect 18922 25942 18932 25994
rect 18956 25942 18986 25994
rect 18986 25942 18998 25994
rect 18998 25942 19012 25994
rect 19036 25942 19050 25994
rect 19050 25942 19062 25994
rect 19062 25942 19092 25994
rect 19116 25942 19126 25994
rect 19126 25942 19172 25994
rect 18876 25940 18932 25942
rect 18956 25940 19012 25942
rect 19036 25940 19092 25942
rect 19116 25940 19172 25942
rect 18876 24906 18932 24908
rect 18956 24906 19012 24908
rect 19036 24906 19092 24908
rect 19116 24906 19172 24908
rect 18876 24854 18922 24906
rect 18922 24854 18932 24906
rect 18956 24854 18986 24906
rect 18986 24854 18998 24906
rect 18998 24854 19012 24906
rect 19036 24854 19050 24906
rect 19050 24854 19062 24906
rect 19062 24854 19092 24906
rect 19116 24854 19126 24906
rect 19126 24854 19172 24906
rect 18876 24852 18932 24854
rect 18956 24852 19012 24854
rect 19036 24852 19092 24854
rect 19116 24852 19172 24854
rect 18876 23818 18932 23820
rect 18956 23818 19012 23820
rect 19036 23818 19092 23820
rect 19116 23818 19172 23820
rect 18876 23766 18922 23818
rect 18922 23766 18932 23818
rect 18956 23766 18986 23818
rect 18986 23766 18998 23818
rect 18998 23766 19012 23818
rect 19036 23766 19050 23818
rect 19050 23766 19062 23818
rect 19062 23766 19092 23818
rect 19116 23766 19126 23818
rect 19126 23766 19172 23818
rect 18876 23764 18932 23766
rect 18956 23764 19012 23766
rect 19036 23764 19092 23766
rect 19116 23764 19172 23766
rect 18876 22730 18932 22732
rect 18956 22730 19012 22732
rect 19036 22730 19092 22732
rect 19116 22730 19172 22732
rect 18876 22678 18922 22730
rect 18922 22678 18932 22730
rect 18956 22678 18986 22730
rect 18986 22678 18998 22730
rect 18998 22678 19012 22730
rect 19036 22678 19050 22730
rect 19050 22678 19062 22730
rect 19062 22678 19092 22730
rect 19116 22678 19126 22730
rect 19126 22678 19172 22730
rect 18876 22676 18932 22678
rect 18956 22676 19012 22678
rect 19036 22676 19092 22678
rect 19116 22676 19172 22678
rect 18876 21642 18932 21644
rect 18956 21642 19012 21644
rect 19036 21642 19092 21644
rect 19116 21642 19172 21644
rect 18876 21590 18922 21642
rect 18922 21590 18932 21642
rect 18956 21590 18986 21642
rect 18986 21590 18998 21642
rect 18998 21590 19012 21642
rect 19036 21590 19050 21642
rect 19050 21590 19062 21642
rect 19062 21590 19092 21642
rect 19116 21590 19126 21642
rect 19126 21590 19172 21642
rect 18876 21588 18932 21590
rect 18956 21588 19012 21590
rect 19036 21588 19092 21590
rect 19116 21588 19172 21590
rect 18876 20554 18932 20556
rect 18956 20554 19012 20556
rect 19036 20554 19092 20556
rect 19116 20554 19172 20556
rect 18876 20502 18922 20554
rect 18922 20502 18932 20554
rect 18956 20502 18986 20554
rect 18986 20502 18998 20554
rect 18998 20502 19012 20554
rect 19036 20502 19050 20554
rect 19050 20502 19062 20554
rect 19062 20502 19092 20554
rect 19116 20502 19126 20554
rect 19126 20502 19172 20554
rect 18876 20500 18932 20502
rect 18956 20500 19012 20502
rect 19036 20500 19092 20502
rect 19116 20500 19172 20502
rect 18876 19466 18932 19468
rect 18956 19466 19012 19468
rect 19036 19466 19092 19468
rect 19116 19466 19172 19468
rect 18876 19414 18922 19466
rect 18922 19414 18932 19466
rect 18956 19414 18986 19466
rect 18986 19414 18998 19466
rect 18998 19414 19012 19466
rect 19036 19414 19050 19466
rect 19050 19414 19062 19466
rect 19062 19414 19092 19466
rect 19116 19414 19126 19466
rect 19126 19414 19172 19466
rect 18876 19412 18932 19414
rect 18956 19412 19012 19414
rect 19036 19412 19092 19414
rect 19116 19412 19172 19414
rect 18876 18378 18932 18380
rect 18956 18378 19012 18380
rect 19036 18378 19092 18380
rect 19116 18378 19172 18380
rect 18876 18326 18922 18378
rect 18922 18326 18932 18378
rect 18956 18326 18986 18378
rect 18986 18326 18998 18378
rect 18998 18326 19012 18378
rect 19036 18326 19050 18378
rect 19050 18326 19062 18378
rect 19062 18326 19092 18378
rect 19116 18326 19126 18378
rect 19126 18326 19172 18378
rect 18876 18324 18932 18326
rect 18956 18324 19012 18326
rect 19036 18324 19092 18326
rect 19116 18324 19172 18326
rect 18876 17290 18932 17292
rect 18956 17290 19012 17292
rect 19036 17290 19092 17292
rect 19116 17290 19172 17292
rect 18876 17238 18922 17290
rect 18922 17238 18932 17290
rect 18956 17238 18986 17290
rect 18986 17238 18998 17290
rect 18998 17238 19012 17290
rect 19036 17238 19050 17290
rect 19050 17238 19062 17290
rect 19062 17238 19092 17290
rect 19116 17238 19126 17290
rect 19126 17238 19172 17290
rect 18876 17236 18932 17238
rect 18956 17236 19012 17238
rect 19036 17236 19092 17238
rect 19116 17236 19172 17238
rect 18876 16202 18932 16204
rect 18956 16202 19012 16204
rect 19036 16202 19092 16204
rect 19116 16202 19172 16204
rect 18876 16150 18922 16202
rect 18922 16150 18932 16202
rect 18956 16150 18986 16202
rect 18986 16150 18998 16202
rect 18998 16150 19012 16202
rect 19036 16150 19050 16202
rect 19050 16150 19062 16202
rect 19062 16150 19092 16202
rect 19116 16150 19126 16202
rect 19126 16150 19172 16202
rect 18876 16148 18932 16150
rect 18956 16148 19012 16150
rect 19036 16148 19092 16150
rect 19116 16148 19172 16150
rect 18876 15114 18932 15116
rect 18956 15114 19012 15116
rect 19036 15114 19092 15116
rect 19116 15114 19172 15116
rect 18876 15062 18922 15114
rect 18922 15062 18932 15114
rect 18956 15062 18986 15114
rect 18986 15062 18998 15114
rect 18998 15062 19012 15114
rect 19036 15062 19050 15114
rect 19050 15062 19062 15114
rect 19062 15062 19092 15114
rect 19116 15062 19126 15114
rect 19126 15062 19172 15114
rect 18876 15060 18932 15062
rect 18956 15060 19012 15062
rect 19036 15060 19092 15062
rect 19116 15060 19172 15062
rect 18876 14026 18932 14028
rect 18956 14026 19012 14028
rect 19036 14026 19092 14028
rect 19116 14026 19172 14028
rect 18876 13974 18922 14026
rect 18922 13974 18932 14026
rect 18956 13974 18986 14026
rect 18986 13974 18998 14026
rect 18998 13974 19012 14026
rect 19036 13974 19050 14026
rect 19050 13974 19062 14026
rect 19062 13974 19092 14026
rect 19116 13974 19126 14026
rect 19126 13974 19172 14026
rect 18876 13972 18932 13974
rect 18956 13972 19012 13974
rect 19036 13972 19092 13974
rect 19116 13972 19172 13974
rect 21210 19616 21266 19672
rect 24338 24648 24394 24704
rect 25350 25056 25406 25112
rect 24430 22608 24486 22664
rect 23142 19616 23198 19672
rect 22314 17712 22370 17768
rect 21486 13632 21542 13688
rect 18876 12938 18932 12940
rect 18956 12938 19012 12940
rect 19036 12938 19092 12940
rect 19116 12938 19172 12940
rect 18876 12886 18922 12938
rect 18922 12886 18932 12938
rect 18956 12886 18986 12938
rect 18986 12886 18998 12938
rect 18998 12886 19012 12938
rect 19036 12886 19050 12938
rect 19050 12886 19062 12938
rect 19062 12886 19092 12938
rect 19116 12886 19126 12938
rect 19126 12886 19172 12938
rect 18876 12884 18932 12886
rect 18956 12884 19012 12886
rect 19036 12884 19092 12886
rect 19116 12884 19172 12886
rect 18876 11850 18932 11852
rect 18956 11850 19012 11852
rect 19036 11850 19092 11852
rect 19116 11850 19172 11852
rect 18876 11798 18922 11850
rect 18922 11798 18932 11850
rect 18956 11798 18986 11850
rect 18986 11798 18998 11850
rect 18998 11798 19012 11850
rect 19036 11798 19050 11850
rect 19050 11798 19062 11850
rect 19062 11798 19092 11850
rect 19116 11798 19126 11850
rect 19126 11798 19172 11850
rect 18876 11796 18932 11798
rect 18956 11796 19012 11798
rect 19036 11796 19092 11798
rect 19116 11796 19172 11798
rect 18876 10762 18932 10764
rect 18956 10762 19012 10764
rect 19036 10762 19092 10764
rect 19116 10762 19172 10764
rect 18876 10710 18922 10762
rect 18922 10710 18932 10762
rect 18956 10710 18986 10762
rect 18986 10710 18998 10762
rect 18998 10710 19012 10762
rect 19036 10710 19050 10762
rect 19050 10710 19062 10762
rect 19062 10710 19092 10762
rect 19116 10710 19126 10762
rect 19126 10710 19172 10762
rect 18876 10708 18932 10710
rect 18956 10708 19012 10710
rect 19036 10708 19092 10710
rect 19116 10708 19172 10710
rect 17622 7648 17678 7704
rect 18876 9674 18932 9676
rect 18956 9674 19012 9676
rect 19036 9674 19092 9676
rect 19116 9674 19172 9676
rect 18876 9622 18922 9674
rect 18922 9622 18932 9674
rect 18956 9622 18986 9674
rect 18986 9622 18998 9674
rect 18998 9622 19012 9674
rect 19036 9622 19050 9674
rect 19050 9622 19062 9674
rect 19062 9622 19092 9674
rect 19116 9622 19126 9674
rect 19126 9622 19172 9674
rect 18876 9620 18932 9622
rect 18956 9620 19012 9622
rect 19036 9620 19092 9622
rect 19116 9620 19172 9622
rect 18876 8586 18932 8588
rect 18956 8586 19012 8588
rect 19036 8586 19092 8588
rect 19116 8586 19172 8588
rect 18876 8534 18922 8586
rect 18922 8534 18932 8586
rect 18956 8534 18986 8586
rect 18986 8534 18998 8586
rect 18998 8534 19012 8586
rect 19036 8534 19050 8586
rect 19050 8534 19062 8586
rect 19062 8534 19092 8586
rect 19116 8534 19126 8586
rect 19126 8534 19172 8586
rect 18876 8532 18932 8534
rect 18956 8532 19012 8534
rect 19036 8532 19092 8534
rect 19116 8532 19172 8534
rect 18876 7498 18932 7500
rect 18956 7498 19012 7500
rect 19036 7498 19092 7500
rect 19116 7498 19172 7500
rect 18876 7446 18922 7498
rect 18922 7446 18932 7498
rect 18956 7446 18986 7498
rect 18986 7446 18998 7498
rect 18998 7446 19012 7498
rect 19036 7446 19050 7498
rect 19050 7446 19062 7498
rect 19062 7446 19092 7498
rect 19116 7446 19126 7498
rect 19126 7446 19172 7498
rect 18876 7444 18932 7446
rect 18956 7444 19012 7446
rect 19036 7444 19092 7446
rect 19116 7444 19172 7446
rect 18876 6410 18932 6412
rect 18956 6410 19012 6412
rect 19036 6410 19092 6412
rect 19116 6410 19172 6412
rect 18876 6358 18922 6410
rect 18922 6358 18932 6410
rect 18956 6358 18986 6410
rect 18986 6358 18998 6410
rect 18998 6358 19012 6410
rect 19036 6358 19050 6410
rect 19050 6358 19062 6410
rect 19062 6358 19092 6410
rect 19116 6358 19126 6410
rect 19126 6358 19172 6410
rect 18876 6356 18932 6358
rect 18956 6356 19012 6358
rect 19036 6356 19092 6358
rect 19116 6356 19172 6358
rect 18876 5322 18932 5324
rect 18956 5322 19012 5324
rect 19036 5322 19092 5324
rect 19116 5322 19172 5324
rect 18876 5270 18922 5322
rect 18922 5270 18932 5322
rect 18956 5270 18986 5322
rect 18986 5270 18998 5322
rect 18998 5270 19012 5322
rect 19036 5270 19050 5322
rect 19050 5270 19062 5322
rect 19062 5270 19092 5322
rect 19116 5270 19126 5322
rect 19126 5270 19172 5322
rect 18876 5268 18932 5270
rect 18956 5268 19012 5270
rect 19036 5268 19092 5270
rect 19116 5268 19172 5270
rect 25258 10096 25314 10152
rect 17254 4520 17310 4576
rect 17438 3704 17494 3760
rect 18876 4234 18932 4236
rect 18956 4234 19012 4236
rect 19036 4234 19092 4236
rect 19116 4234 19172 4236
rect 18876 4182 18922 4234
rect 18922 4182 18932 4234
rect 18956 4182 18986 4234
rect 18986 4182 18998 4234
rect 18998 4182 19012 4234
rect 19036 4182 19050 4234
rect 19050 4182 19062 4234
rect 19062 4182 19092 4234
rect 19116 4182 19126 4234
rect 19126 4182 19172 4234
rect 18876 4180 18932 4182
rect 18956 4180 19012 4182
rect 19036 4180 19092 4182
rect 19116 4180 19172 4182
rect 18082 3840 18138 3896
rect 18876 3146 18932 3148
rect 18956 3146 19012 3148
rect 19036 3146 19092 3148
rect 19116 3146 19172 3148
rect 18876 3094 18922 3146
rect 18922 3094 18932 3146
rect 18956 3094 18986 3146
rect 18986 3094 18998 3146
rect 18998 3094 19012 3146
rect 19036 3094 19050 3146
rect 19050 3094 19062 3146
rect 19062 3094 19092 3146
rect 19116 3094 19126 3146
rect 19126 3094 19172 3146
rect 18876 3092 18932 3094
rect 18956 3092 19012 3094
rect 19036 3092 19092 3094
rect 19116 3092 19172 3094
rect 17898 1800 17954 1856
rect 18082 1800 18138 1856
rect 18876 2058 18932 2060
rect 18956 2058 19012 2060
rect 19036 2058 19092 2060
rect 19116 2058 19172 2060
rect 18876 2006 18922 2058
rect 18922 2006 18932 2058
rect 18956 2006 18986 2058
rect 18986 2006 18998 2058
rect 18998 2006 19012 2058
rect 19036 2006 19050 2058
rect 19050 2006 19062 2058
rect 19062 2006 19092 2058
rect 19116 2006 19126 2058
rect 19126 2006 19172 2058
rect 18876 2004 18932 2006
rect 18956 2004 19012 2006
rect 19036 2004 19092 2006
rect 19116 2004 19172 2006
rect 18634 1120 18690 1176
rect 19278 1120 19334 1176
rect 18876 970 18932 972
rect 18956 970 19012 972
rect 19036 970 19092 972
rect 19116 970 19172 972
rect 18876 918 18922 970
rect 18922 918 18932 970
rect 18956 918 18986 970
rect 18986 918 18998 970
rect 18998 918 19012 970
rect 19036 918 19050 970
rect 19050 918 19062 970
rect 19062 918 19092 970
rect 19116 918 19126 970
rect 19126 918 19172 970
rect 18876 916 18932 918
rect 18956 916 19012 918
rect 19036 916 19092 918
rect 19116 916 19172 918
rect 23418 1936 23474 1992
rect 25442 19208 25498 19264
rect 26178 19344 26234 19400
rect 26178 18120 26234 18176
rect 26362 16624 26418 16680
rect 23510 1800 23566 1856
rect 24890 1140 24946 1176
rect 24890 1120 24892 1140
rect 24892 1120 24944 1140
rect 24944 1120 24946 1140
rect 3516 372 3572 374
rect 3596 372 3652 374
rect 3676 372 3732 374
rect 3756 372 3812 374
<< metal3 >>
rect 0 27018 432 27274
rect 18864 27088 19184 27104
rect 18864 27024 18872 27088
rect 18936 27024 18952 27088
rect 19016 27024 19032 27088
rect 19096 27024 19112 27088
rect 19176 27024 19184 27088
rect 873 27018 939 27021
rect 0 27016 939 27018
rect 0 26974 878 27016
rect 386 26960 878 26974
rect 934 26960 939 27016
rect 18864 27008 19184 27024
rect 386 26958 939 26960
rect 873 26955 939 26958
rect 3504 26544 3824 26560
rect 3504 26480 3512 26544
rect 3576 26480 3592 26544
rect 3656 26480 3672 26544
rect 3736 26480 3752 26544
rect 3816 26480 3824 26544
rect 3504 26464 3824 26480
rect 18864 26000 19184 26016
rect 18864 25936 18872 26000
rect 18936 25936 18952 26000
rect 19016 25936 19032 26000
rect 19096 25936 19112 26000
rect 19176 25936 19184 26000
rect 18864 25920 19184 25936
rect 27303 25658 27735 25914
rect 27289 25614 27735 25658
rect 3504 25456 3824 25472
rect 3504 25392 3512 25456
rect 3576 25392 3592 25456
rect 3656 25392 3672 25456
rect 3736 25392 3752 25456
rect 3816 25392 3824 25456
rect 3504 25376 3824 25392
rect 25345 25114 25411 25117
rect 27289 25114 27349 25614
rect 25345 25112 27349 25114
rect 25345 25056 25350 25112
rect 25406 25056 27349 25112
rect 25345 25054 27349 25056
rect 25345 25051 25411 25054
rect 18864 24912 19184 24928
rect 18864 24848 18872 24912
rect 18936 24848 18952 24912
rect 19016 24848 19032 24912
rect 19096 24848 19112 24912
rect 19176 24848 19184 24912
rect 18864 24832 19184 24848
rect 6485 24706 6551 24709
rect 24333 24706 24399 24709
rect 6485 24704 24399 24706
rect 6485 24648 6490 24704
rect 6546 24648 24338 24704
rect 24394 24648 24399 24704
rect 6485 24646 24399 24648
rect 6485 24643 6551 24646
rect 24333 24643 24399 24646
rect 3504 24368 3824 24384
rect 3504 24304 3512 24368
rect 3576 24304 3592 24368
rect 3656 24304 3672 24368
rect 3736 24304 3752 24368
rect 3816 24304 3824 24368
rect 3504 24288 3824 24304
rect 0 24026 432 24282
rect 1425 24026 1491 24029
rect 0 24024 1491 24026
rect 0 23982 1430 24024
rect 386 23968 1430 23982
rect 1486 23968 1491 24024
rect 386 23966 1491 23968
rect 1425 23963 1491 23966
rect 18864 23824 19184 23840
rect 18864 23760 18872 23824
rect 18936 23760 18952 23824
rect 19016 23760 19032 23824
rect 19096 23760 19112 23824
rect 19176 23760 19184 23824
rect 18864 23744 19184 23760
rect 3504 23280 3824 23296
rect 3504 23216 3512 23280
rect 3576 23216 3592 23280
rect 3656 23216 3672 23280
rect 3736 23216 3752 23280
rect 3816 23216 3824 23280
rect 3504 23200 3824 23216
rect 18864 22736 19184 22752
rect 18864 22672 18872 22736
rect 18936 22672 18952 22736
rect 19016 22672 19032 22736
rect 19096 22672 19112 22736
rect 19176 22672 19184 22736
rect 18864 22656 19184 22672
rect 24425 22666 24491 22669
rect 27303 22666 27735 22922
rect 24425 22664 27735 22666
rect 24425 22608 24430 22664
rect 24486 22622 27735 22664
rect 24486 22608 27349 22622
rect 24425 22606 27349 22608
rect 24425 22603 24491 22606
rect 3504 22192 3824 22208
rect 3504 22128 3512 22192
rect 3576 22128 3592 22192
rect 3656 22128 3672 22192
rect 3736 22128 3752 22192
rect 3816 22128 3824 22192
rect 3504 22112 3824 22128
rect 18864 21648 19184 21664
rect 18864 21584 18872 21648
rect 18936 21584 18952 21648
rect 19016 21584 19032 21648
rect 19096 21584 19112 21648
rect 19176 21584 19184 21648
rect 18864 21568 19184 21584
rect 0 21034 432 21290
rect 3504 21104 3824 21120
rect 3504 21040 3512 21104
rect 3576 21040 3592 21104
rect 3656 21040 3672 21104
rect 3736 21040 3752 21104
rect 3816 21040 3824 21104
rect 873 21034 939 21037
rect 0 21032 939 21034
rect 0 20990 878 21032
rect 386 20976 878 20990
rect 934 20976 939 21032
rect 3504 21024 3824 21040
rect 386 20974 939 20976
rect 873 20971 939 20974
rect 18864 20560 19184 20576
rect 18864 20496 18872 20560
rect 18936 20496 18952 20560
rect 19016 20496 19032 20560
rect 19096 20496 19112 20560
rect 19176 20496 19184 20560
rect 18864 20480 19184 20496
rect 3504 20016 3824 20032
rect 3504 19952 3512 20016
rect 3576 19952 3592 20016
rect 3656 19952 3672 20016
rect 3736 19952 3752 20016
rect 3816 19952 3824 20016
rect 3504 19936 3824 19952
rect 21205 19674 21271 19677
rect 23137 19674 23203 19677
rect 27303 19674 27735 19930
rect 21205 19672 23203 19674
rect 21205 19616 21210 19672
rect 21266 19616 23142 19672
rect 23198 19616 23203 19672
rect 21205 19614 23203 19616
rect 21205 19611 21271 19614
rect 23137 19611 23203 19614
rect 27289 19630 27735 19674
rect 18864 19472 19184 19488
rect 18864 19408 18872 19472
rect 18936 19408 18952 19472
rect 19016 19408 19032 19472
rect 19096 19408 19112 19472
rect 19176 19408 19184 19472
rect 18864 19392 19184 19408
rect 26173 19402 26239 19405
rect 27289 19402 27349 19630
rect 26173 19400 27349 19402
rect 26173 19344 26178 19400
rect 26234 19344 27349 19400
rect 26173 19342 27349 19344
rect 26173 19339 26239 19342
rect 13569 19266 13635 19269
rect 25437 19266 25503 19269
rect 13569 19264 25503 19266
rect 13569 19208 13574 19264
rect 13630 19208 25442 19264
rect 25498 19208 25503 19264
rect 13569 19206 25503 19208
rect 13569 19203 13635 19206
rect 25437 19203 25503 19206
rect 3504 18928 3824 18944
rect 3504 18864 3512 18928
rect 3576 18864 3592 18928
rect 3656 18864 3672 18928
rect 3736 18864 3752 18928
rect 3816 18864 3824 18928
rect 3504 18848 3824 18864
rect 18864 18384 19184 18400
rect 18864 18320 18872 18384
rect 18936 18320 18952 18384
rect 19016 18320 19032 18384
rect 19096 18320 19112 18384
rect 19176 18320 19184 18384
rect 18864 18304 19184 18320
rect 0 18042 432 18298
rect 9981 18178 10047 18181
rect 26173 18178 26239 18181
rect 9981 18176 26239 18178
rect 9981 18120 9986 18176
rect 10042 18120 26178 18176
rect 26234 18120 26239 18176
rect 9981 18118 26239 18120
rect 9981 18115 10047 18118
rect 26173 18115 26239 18118
rect 873 18042 939 18045
rect 0 18040 939 18042
rect 0 17998 878 18040
rect 386 17984 878 17998
rect 934 17984 939 18040
rect 386 17982 939 17984
rect 873 17979 939 17982
rect 3504 17840 3824 17856
rect 3504 17776 3512 17840
rect 3576 17776 3592 17840
rect 3656 17776 3672 17840
rect 3736 17776 3752 17840
rect 3816 17776 3824 17840
rect 3504 17760 3824 17776
rect 12373 17770 12439 17773
rect 22309 17770 22375 17773
rect 12373 17768 22375 17770
rect 12373 17712 12378 17768
rect 12434 17712 22314 17768
rect 22370 17712 22375 17768
rect 12373 17710 22375 17712
rect 12373 17707 12439 17710
rect 22309 17707 22375 17710
rect 2345 17634 2411 17637
rect 15133 17634 15199 17637
rect 2345 17632 15199 17634
rect 2345 17576 2350 17632
rect 2406 17576 15138 17632
rect 15194 17576 15199 17632
rect 2345 17574 15199 17576
rect 2345 17571 2411 17574
rect 15133 17571 15199 17574
rect 18864 17296 19184 17312
rect 18864 17232 18872 17296
rect 18936 17232 18952 17296
rect 19016 17232 19032 17296
rect 19096 17232 19112 17296
rect 19176 17232 19184 17296
rect 18864 17216 19184 17232
rect 3504 16752 3824 16768
rect 3504 16688 3512 16752
rect 3576 16688 3592 16752
rect 3656 16688 3672 16752
rect 3736 16688 3752 16752
rect 3816 16688 3824 16752
rect 3504 16672 3824 16688
rect 26357 16682 26423 16685
rect 27303 16682 27735 16938
rect 26357 16680 27735 16682
rect 26357 16624 26362 16680
rect 26418 16638 27735 16680
rect 26418 16624 27349 16638
rect 26357 16622 27349 16624
rect 26357 16619 26423 16622
rect 18864 16208 19184 16224
rect 18864 16144 18872 16208
rect 18936 16144 18952 16208
rect 19016 16144 19032 16208
rect 19096 16144 19112 16208
rect 19176 16144 19184 16208
rect 18864 16128 19184 16144
rect 3504 15664 3824 15680
rect 3504 15600 3512 15664
rect 3576 15600 3592 15664
rect 3656 15600 3672 15664
rect 3736 15600 3752 15664
rect 3816 15600 3824 15664
rect 3504 15584 3824 15600
rect 1977 15458 2043 15461
rect 2989 15458 3055 15461
rect 1977 15456 3055 15458
rect 1977 15400 1982 15456
rect 2038 15400 2994 15456
rect 3050 15400 3055 15456
rect 1977 15398 3055 15400
rect 1977 15395 2043 15398
rect 2989 15395 3055 15398
rect 0 15050 432 15306
rect 1701 15186 1767 15189
rect 7865 15186 7931 15189
rect 1701 15184 7931 15186
rect 1701 15128 1706 15184
rect 1762 15128 7870 15184
rect 7926 15128 7931 15184
rect 1701 15126 7931 15128
rect 1701 15123 1767 15126
rect 7865 15123 7931 15126
rect 18864 15120 19184 15136
rect 18864 15056 18872 15120
rect 18936 15056 18952 15120
rect 19016 15056 19032 15120
rect 19096 15056 19112 15120
rect 19176 15056 19184 15120
rect 873 15050 939 15053
rect 0 15048 939 15050
rect 0 15006 878 15048
rect 386 14992 878 15006
rect 934 14992 939 15048
rect 18864 15040 19184 15056
rect 386 14990 939 14992
rect 873 14987 939 14990
rect 4921 14642 4987 14645
rect 5197 14642 5263 14645
rect 4921 14640 5263 14642
rect 3504 14576 3824 14592
rect 4921 14584 4926 14640
rect 4982 14584 5202 14640
rect 5258 14584 5263 14640
rect 4921 14582 5263 14584
rect 4921 14579 4987 14582
rect 5197 14579 5263 14582
rect 3504 14512 3512 14576
rect 3576 14512 3592 14576
rect 3656 14512 3672 14576
rect 3736 14512 3752 14576
rect 3816 14512 3824 14576
rect 3504 14496 3824 14512
rect 3265 14234 3331 14237
rect 4277 14234 4343 14237
rect 3265 14232 4343 14234
rect 3265 14176 3270 14232
rect 3326 14176 4282 14232
rect 4338 14176 4343 14232
rect 3265 14174 4343 14176
rect 3265 14171 3331 14174
rect 4277 14171 4343 14174
rect 10625 14234 10691 14237
rect 12189 14234 12255 14237
rect 10625 14232 12255 14234
rect 10625 14176 10630 14232
rect 10686 14176 12194 14232
rect 12250 14176 12255 14232
rect 10625 14174 12255 14176
rect 10625 14171 10691 14174
rect 12189 14171 12255 14174
rect 6669 14098 6735 14101
rect 10165 14098 10231 14101
rect 10625 14098 10691 14101
rect 12833 14098 12899 14101
rect 6669 14096 10231 14098
rect 6669 14040 6674 14096
rect 6730 14040 10170 14096
rect 10226 14040 10231 14096
rect 6669 14038 10231 14040
rect 6669 14035 6735 14038
rect 10165 14035 10231 14038
rect 10398 14096 12899 14098
rect 10398 14040 10630 14096
rect 10686 14040 12838 14096
rect 12894 14040 12899 14096
rect 10398 14038 12899 14040
rect 9521 13962 9587 13965
rect 10398 13962 10458 14038
rect 10625 14035 10691 14038
rect 12833 14035 12899 14038
rect 9521 13960 10458 13962
rect 9521 13904 9526 13960
rect 9582 13904 10458 13960
rect 18864 14032 19184 14048
rect 18864 13968 18872 14032
rect 18936 13968 18952 14032
rect 19016 13968 19032 14032
rect 19096 13968 19112 14032
rect 19176 13968 19184 14032
rect 18864 13952 19184 13968
rect 9521 13902 10458 13904
rect 9521 13899 9587 13902
rect 21481 13690 21547 13693
rect 27303 13690 27735 13946
rect 21481 13688 27735 13690
rect 21481 13632 21486 13688
rect 21542 13646 27735 13688
rect 21542 13632 27349 13646
rect 21481 13630 27349 13632
rect 21481 13627 21547 13630
rect 3504 13488 3824 13504
rect 3504 13424 3512 13488
rect 3576 13424 3592 13488
rect 3656 13424 3672 13488
rect 3736 13424 3752 13488
rect 3816 13424 3824 13488
rect 3504 13408 3824 13424
rect 5657 13010 5723 13013
rect 6853 13010 6919 13013
rect 5657 13008 6919 13010
rect 5657 12952 5662 13008
rect 5718 12952 6858 13008
rect 6914 12952 6919 13008
rect 5657 12950 6919 12952
rect 5657 12947 5723 12950
rect 6853 12947 6919 12950
rect 18864 12944 19184 12960
rect 18864 12880 18872 12944
rect 18936 12880 18952 12944
rect 19016 12880 19032 12944
rect 19096 12880 19112 12944
rect 19176 12880 19184 12944
rect 18864 12864 19184 12880
rect 7129 12738 7195 12741
rect 8233 12738 8299 12741
rect 7129 12736 8299 12738
rect 7129 12680 7134 12736
rect 7190 12680 8238 12736
rect 8294 12680 8299 12736
rect 7129 12678 8299 12680
rect 7129 12675 7195 12678
rect 8233 12675 8299 12678
rect 3504 12400 3824 12416
rect 3504 12336 3512 12400
rect 3576 12336 3592 12400
rect 3656 12336 3672 12400
rect 3736 12336 3752 12400
rect 3816 12336 3824 12400
rect 3504 12320 3824 12336
rect 0 12058 432 12314
rect 689 12058 755 12061
rect 0 12056 755 12058
rect 0 12014 694 12056
rect 386 12000 694 12014
rect 750 12000 755 12056
rect 386 11998 755 12000
rect 689 11995 755 11998
rect 18864 11856 19184 11872
rect 18864 11792 18872 11856
rect 18936 11792 18952 11856
rect 19016 11792 19032 11856
rect 19096 11792 19112 11856
rect 19176 11792 19184 11856
rect 18864 11776 19184 11792
rect 3504 11312 3824 11328
rect 3504 11248 3512 11312
rect 3576 11248 3592 11312
rect 3656 11248 3672 11312
rect 3736 11248 3752 11312
rect 3816 11248 3824 11312
rect 3504 11232 3824 11248
rect 18864 10768 19184 10784
rect 18864 10704 18872 10768
rect 18936 10704 18952 10768
rect 19016 10704 19032 10768
rect 19096 10704 19112 10768
rect 19176 10704 19184 10768
rect 18864 10688 19184 10704
rect 27303 10698 27735 10954
rect 27289 10654 27735 10698
rect 3504 10224 3824 10240
rect 3504 10160 3512 10224
rect 3576 10160 3592 10224
rect 3656 10160 3672 10224
rect 3736 10160 3752 10224
rect 3816 10160 3824 10224
rect 3504 10144 3824 10160
rect 25253 10154 25319 10157
rect 27289 10154 27349 10654
rect 25253 10152 27349 10154
rect 25253 10096 25258 10152
rect 25314 10096 27349 10152
rect 25253 10094 27349 10096
rect 25253 10091 25319 10094
rect 18864 9680 19184 9696
rect 18864 9616 18872 9680
rect 18936 9616 18952 9680
rect 19016 9616 19032 9680
rect 19096 9616 19112 9680
rect 19176 9616 19184 9680
rect 18864 9600 19184 9616
rect 0 9066 432 9322
rect 3504 9136 3824 9152
rect 3504 9072 3512 9136
rect 3576 9072 3592 9136
rect 3656 9072 3672 9136
rect 3736 9072 3752 9136
rect 3816 9072 3824 9136
rect 689 9066 755 9069
rect 0 9064 755 9066
rect 0 9022 694 9064
rect 386 9008 694 9022
rect 750 9008 755 9064
rect 3504 9056 3824 9072
rect 386 9006 755 9008
rect 689 9003 755 9006
rect 18864 8592 19184 8608
rect 18864 8528 18872 8592
rect 18936 8528 18952 8592
rect 19016 8528 19032 8592
rect 19096 8528 19112 8592
rect 19176 8528 19184 8592
rect 18864 8512 19184 8528
rect 3504 8048 3824 8064
rect 3504 7984 3512 8048
rect 3576 7984 3592 8048
rect 3656 7984 3672 8048
rect 3736 7984 3752 8048
rect 3816 7984 3824 8048
rect 3504 7968 3824 7984
rect 17617 7706 17683 7709
rect 27303 7706 27735 7962
rect 17617 7704 27735 7706
rect 17617 7648 17622 7704
rect 17678 7662 27735 7704
rect 17678 7648 27349 7662
rect 17617 7646 27349 7648
rect 17617 7643 17683 7646
rect 18864 7504 19184 7520
rect 18864 7440 18872 7504
rect 18936 7440 18952 7504
rect 19016 7440 19032 7504
rect 19096 7440 19112 7504
rect 19176 7440 19184 7504
rect 18864 7424 19184 7440
rect 3504 6960 3824 6976
rect 3504 6896 3512 6960
rect 3576 6896 3592 6960
rect 3656 6896 3672 6960
rect 3736 6896 3752 6960
rect 3816 6896 3824 6960
rect 3504 6880 3824 6896
rect 18864 6416 19184 6432
rect 18864 6352 18872 6416
rect 18936 6352 18952 6416
rect 19016 6352 19032 6416
rect 19096 6352 19112 6416
rect 19176 6352 19184 6416
rect 18864 6336 19184 6352
rect 0 6074 432 6330
rect 873 6074 939 6077
rect 0 6072 939 6074
rect 0 6030 878 6072
rect 386 6016 878 6030
rect 934 6016 939 6072
rect 386 6014 939 6016
rect 873 6011 939 6014
rect 3504 5872 3824 5888
rect 3504 5808 3512 5872
rect 3576 5808 3592 5872
rect 3656 5808 3672 5872
rect 3736 5808 3752 5872
rect 3816 5808 3824 5872
rect 3504 5792 3824 5808
rect 18864 5328 19184 5344
rect 18864 5264 18872 5328
rect 18936 5264 18952 5328
rect 19016 5264 19032 5328
rect 19096 5264 19112 5328
rect 19176 5264 19184 5328
rect 18864 5248 19184 5264
rect 27303 4986 27735 5242
rect 27289 4942 27735 4986
rect 3504 4784 3824 4800
rect 3504 4720 3512 4784
rect 3576 4720 3592 4784
rect 3656 4720 3672 4784
rect 3736 4720 3752 4784
rect 3816 4720 3824 4784
rect 3504 4704 3824 4720
rect 17249 4578 17315 4581
rect 27289 4578 27349 4942
rect 17249 4576 27349 4578
rect 17249 4520 17254 4576
rect 17310 4520 27349 4576
rect 17249 4518 27349 4520
rect 17249 4515 17315 4518
rect 18864 4240 19184 4256
rect 18864 4176 18872 4240
rect 18936 4176 18952 4240
rect 19016 4176 19032 4240
rect 19096 4176 19112 4240
rect 19176 4176 19184 4240
rect 18864 4160 19184 4176
rect 1425 3898 1491 3901
rect 18077 3898 18143 3901
rect 1425 3896 18143 3898
rect 1425 3840 1430 3896
rect 1486 3840 18082 3896
rect 18138 3840 18143 3896
rect 1425 3838 18143 3840
rect 1425 3835 1491 3838
rect 18077 3835 18143 3838
rect 7037 3762 7103 3765
rect 17433 3762 17499 3765
rect 7037 3760 17499 3762
rect 3504 3696 3824 3712
rect 7037 3704 7042 3760
rect 7098 3704 17438 3760
rect 17494 3704 17499 3760
rect 7037 3702 17499 3704
rect 7037 3699 7103 3702
rect 17433 3699 17499 3702
rect 3504 3632 3512 3696
rect 3576 3632 3592 3696
rect 3656 3632 3672 3696
rect 3736 3632 3752 3696
rect 3816 3632 3824 3696
rect 3504 3616 3824 3632
rect 0 3085 432 3338
rect 18864 3152 19184 3168
rect 18864 3088 18872 3152
rect 18936 3088 18952 3152
rect 19016 3088 19032 3152
rect 19096 3088 19112 3152
rect 19176 3088 19184 3152
rect 0 3082 479 3085
rect 0 3080 576 3082
rect 0 3038 418 3080
rect 386 3024 418 3038
rect 474 3024 576 3080
rect 18864 3072 19184 3088
rect 386 3022 576 3024
rect 413 3019 479 3022
rect 3504 2608 3824 2624
rect 3504 2544 3512 2608
rect 3576 2544 3592 2608
rect 3656 2544 3672 2608
rect 3736 2544 3752 2608
rect 3816 2544 3824 2608
rect 3504 2528 3824 2544
rect 18864 2064 19184 2080
rect 18864 2000 18872 2064
rect 18936 2000 18952 2064
rect 19016 2000 19032 2064
rect 19096 2000 19112 2064
rect 19176 2000 19184 2064
rect 18864 1984 19184 2000
rect 23413 1994 23479 1997
rect 27303 1994 27735 2250
rect 23413 1992 27735 1994
rect 23413 1936 23418 1992
rect 23474 1950 27735 1992
rect 23474 1936 27349 1950
rect 23413 1934 27349 1936
rect 23413 1931 23479 1934
rect 413 1858 479 1861
rect 17893 1858 17959 1861
rect 18077 1858 18143 1861
rect 23505 1858 23571 1861
rect 413 1856 23571 1858
rect 413 1800 418 1856
rect 474 1800 17898 1856
rect 17954 1800 18082 1856
rect 18138 1800 23510 1856
rect 23566 1800 23571 1856
rect 413 1798 23571 1800
rect 413 1795 479 1798
rect 17893 1795 17959 1798
rect 18077 1795 18143 1798
rect 23505 1795 23571 1798
rect 3504 1520 3824 1536
rect 3504 1456 3512 1520
rect 3576 1456 3592 1520
rect 3656 1456 3672 1520
rect 3736 1456 3752 1520
rect 3816 1456 3824 1520
rect 3504 1440 3824 1456
rect 18629 1178 18695 1181
rect 19273 1178 19339 1181
rect 24885 1178 24951 1181
rect 18629 1176 24951 1178
rect 18629 1120 18634 1176
rect 18690 1120 19278 1176
rect 19334 1120 24890 1176
rect 24946 1120 24951 1176
rect 18629 1118 24951 1120
rect 18629 1115 18695 1118
rect 19273 1115 19339 1118
rect 24885 1115 24951 1118
rect 18864 976 19184 992
rect 18864 912 18872 976
rect 18936 912 18952 976
rect 19016 912 19032 976
rect 19096 912 19112 976
rect 19176 912 19184 976
rect 18864 896 19184 912
rect 3504 432 3824 448
rect 3504 368 3512 432
rect 3576 368 3592 432
rect 3656 368 3672 432
rect 3736 368 3752 432
rect 3816 368 3824 432
rect 3504 352 3824 368
<< via3 >>
rect 18872 27084 18936 27088
rect 18872 27028 18876 27084
rect 18876 27028 18932 27084
rect 18932 27028 18936 27084
rect 18872 27024 18936 27028
rect 18952 27084 19016 27088
rect 18952 27028 18956 27084
rect 18956 27028 19012 27084
rect 19012 27028 19016 27084
rect 18952 27024 19016 27028
rect 19032 27084 19096 27088
rect 19032 27028 19036 27084
rect 19036 27028 19092 27084
rect 19092 27028 19096 27084
rect 19032 27024 19096 27028
rect 19112 27084 19176 27088
rect 19112 27028 19116 27084
rect 19116 27028 19172 27084
rect 19172 27028 19176 27084
rect 19112 27024 19176 27028
rect 3512 26540 3576 26544
rect 3512 26484 3516 26540
rect 3516 26484 3572 26540
rect 3572 26484 3576 26540
rect 3512 26480 3576 26484
rect 3592 26540 3656 26544
rect 3592 26484 3596 26540
rect 3596 26484 3652 26540
rect 3652 26484 3656 26540
rect 3592 26480 3656 26484
rect 3672 26540 3736 26544
rect 3672 26484 3676 26540
rect 3676 26484 3732 26540
rect 3732 26484 3736 26540
rect 3672 26480 3736 26484
rect 3752 26540 3816 26544
rect 3752 26484 3756 26540
rect 3756 26484 3812 26540
rect 3812 26484 3816 26540
rect 3752 26480 3816 26484
rect 18872 25996 18936 26000
rect 18872 25940 18876 25996
rect 18876 25940 18932 25996
rect 18932 25940 18936 25996
rect 18872 25936 18936 25940
rect 18952 25996 19016 26000
rect 18952 25940 18956 25996
rect 18956 25940 19012 25996
rect 19012 25940 19016 25996
rect 18952 25936 19016 25940
rect 19032 25996 19096 26000
rect 19032 25940 19036 25996
rect 19036 25940 19092 25996
rect 19092 25940 19096 25996
rect 19032 25936 19096 25940
rect 19112 25996 19176 26000
rect 19112 25940 19116 25996
rect 19116 25940 19172 25996
rect 19172 25940 19176 25996
rect 19112 25936 19176 25940
rect 3512 25452 3576 25456
rect 3512 25396 3516 25452
rect 3516 25396 3572 25452
rect 3572 25396 3576 25452
rect 3512 25392 3576 25396
rect 3592 25452 3656 25456
rect 3592 25396 3596 25452
rect 3596 25396 3652 25452
rect 3652 25396 3656 25452
rect 3592 25392 3656 25396
rect 3672 25452 3736 25456
rect 3672 25396 3676 25452
rect 3676 25396 3732 25452
rect 3732 25396 3736 25452
rect 3672 25392 3736 25396
rect 3752 25452 3816 25456
rect 3752 25396 3756 25452
rect 3756 25396 3812 25452
rect 3812 25396 3816 25452
rect 3752 25392 3816 25396
rect 18872 24908 18936 24912
rect 18872 24852 18876 24908
rect 18876 24852 18932 24908
rect 18932 24852 18936 24908
rect 18872 24848 18936 24852
rect 18952 24908 19016 24912
rect 18952 24852 18956 24908
rect 18956 24852 19012 24908
rect 19012 24852 19016 24908
rect 18952 24848 19016 24852
rect 19032 24908 19096 24912
rect 19032 24852 19036 24908
rect 19036 24852 19092 24908
rect 19092 24852 19096 24908
rect 19032 24848 19096 24852
rect 19112 24908 19176 24912
rect 19112 24852 19116 24908
rect 19116 24852 19172 24908
rect 19172 24852 19176 24908
rect 19112 24848 19176 24852
rect 3512 24364 3576 24368
rect 3512 24308 3516 24364
rect 3516 24308 3572 24364
rect 3572 24308 3576 24364
rect 3512 24304 3576 24308
rect 3592 24364 3656 24368
rect 3592 24308 3596 24364
rect 3596 24308 3652 24364
rect 3652 24308 3656 24364
rect 3592 24304 3656 24308
rect 3672 24364 3736 24368
rect 3672 24308 3676 24364
rect 3676 24308 3732 24364
rect 3732 24308 3736 24364
rect 3672 24304 3736 24308
rect 3752 24364 3816 24368
rect 3752 24308 3756 24364
rect 3756 24308 3812 24364
rect 3812 24308 3816 24364
rect 3752 24304 3816 24308
rect 18872 23820 18936 23824
rect 18872 23764 18876 23820
rect 18876 23764 18932 23820
rect 18932 23764 18936 23820
rect 18872 23760 18936 23764
rect 18952 23820 19016 23824
rect 18952 23764 18956 23820
rect 18956 23764 19012 23820
rect 19012 23764 19016 23820
rect 18952 23760 19016 23764
rect 19032 23820 19096 23824
rect 19032 23764 19036 23820
rect 19036 23764 19092 23820
rect 19092 23764 19096 23820
rect 19032 23760 19096 23764
rect 19112 23820 19176 23824
rect 19112 23764 19116 23820
rect 19116 23764 19172 23820
rect 19172 23764 19176 23820
rect 19112 23760 19176 23764
rect 3512 23276 3576 23280
rect 3512 23220 3516 23276
rect 3516 23220 3572 23276
rect 3572 23220 3576 23276
rect 3512 23216 3576 23220
rect 3592 23276 3656 23280
rect 3592 23220 3596 23276
rect 3596 23220 3652 23276
rect 3652 23220 3656 23276
rect 3592 23216 3656 23220
rect 3672 23276 3736 23280
rect 3672 23220 3676 23276
rect 3676 23220 3732 23276
rect 3732 23220 3736 23276
rect 3672 23216 3736 23220
rect 3752 23276 3816 23280
rect 3752 23220 3756 23276
rect 3756 23220 3812 23276
rect 3812 23220 3816 23276
rect 3752 23216 3816 23220
rect 18872 22732 18936 22736
rect 18872 22676 18876 22732
rect 18876 22676 18932 22732
rect 18932 22676 18936 22732
rect 18872 22672 18936 22676
rect 18952 22732 19016 22736
rect 18952 22676 18956 22732
rect 18956 22676 19012 22732
rect 19012 22676 19016 22732
rect 18952 22672 19016 22676
rect 19032 22732 19096 22736
rect 19032 22676 19036 22732
rect 19036 22676 19092 22732
rect 19092 22676 19096 22732
rect 19032 22672 19096 22676
rect 19112 22732 19176 22736
rect 19112 22676 19116 22732
rect 19116 22676 19172 22732
rect 19172 22676 19176 22732
rect 19112 22672 19176 22676
rect 3512 22188 3576 22192
rect 3512 22132 3516 22188
rect 3516 22132 3572 22188
rect 3572 22132 3576 22188
rect 3512 22128 3576 22132
rect 3592 22188 3656 22192
rect 3592 22132 3596 22188
rect 3596 22132 3652 22188
rect 3652 22132 3656 22188
rect 3592 22128 3656 22132
rect 3672 22188 3736 22192
rect 3672 22132 3676 22188
rect 3676 22132 3732 22188
rect 3732 22132 3736 22188
rect 3672 22128 3736 22132
rect 3752 22188 3816 22192
rect 3752 22132 3756 22188
rect 3756 22132 3812 22188
rect 3812 22132 3816 22188
rect 3752 22128 3816 22132
rect 18872 21644 18936 21648
rect 18872 21588 18876 21644
rect 18876 21588 18932 21644
rect 18932 21588 18936 21644
rect 18872 21584 18936 21588
rect 18952 21644 19016 21648
rect 18952 21588 18956 21644
rect 18956 21588 19012 21644
rect 19012 21588 19016 21644
rect 18952 21584 19016 21588
rect 19032 21644 19096 21648
rect 19032 21588 19036 21644
rect 19036 21588 19092 21644
rect 19092 21588 19096 21644
rect 19032 21584 19096 21588
rect 19112 21644 19176 21648
rect 19112 21588 19116 21644
rect 19116 21588 19172 21644
rect 19172 21588 19176 21644
rect 19112 21584 19176 21588
rect 3512 21100 3576 21104
rect 3512 21044 3516 21100
rect 3516 21044 3572 21100
rect 3572 21044 3576 21100
rect 3512 21040 3576 21044
rect 3592 21100 3656 21104
rect 3592 21044 3596 21100
rect 3596 21044 3652 21100
rect 3652 21044 3656 21100
rect 3592 21040 3656 21044
rect 3672 21100 3736 21104
rect 3672 21044 3676 21100
rect 3676 21044 3732 21100
rect 3732 21044 3736 21100
rect 3672 21040 3736 21044
rect 3752 21100 3816 21104
rect 3752 21044 3756 21100
rect 3756 21044 3812 21100
rect 3812 21044 3816 21100
rect 3752 21040 3816 21044
rect 18872 20556 18936 20560
rect 18872 20500 18876 20556
rect 18876 20500 18932 20556
rect 18932 20500 18936 20556
rect 18872 20496 18936 20500
rect 18952 20556 19016 20560
rect 18952 20500 18956 20556
rect 18956 20500 19012 20556
rect 19012 20500 19016 20556
rect 18952 20496 19016 20500
rect 19032 20556 19096 20560
rect 19032 20500 19036 20556
rect 19036 20500 19092 20556
rect 19092 20500 19096 20556
rect 19032 20496 19096 20500
rect 19112 20556 19176 20560
rect 19112 20500 19116 20556
rect 19116 20500 19172 20556
rect 19172 20500 19176 20556
rect 19112 20496 19176 20500
rect 3512 20012 3576 20016
rect 3512 19956 3516 20012
rect 3516 19956 3572 20012
rect 3572 19956 3576 20012
rect 3512 19952 3576 19956
rect 3592 20012 3656 20016
rect 3592 19956 3596 20012
rect 3596 19956 3652 20012
rect 3652 19956 3656 20012
rect 3592 19952 3656 19956
rect 3672 20012 3736 20016
rect 3672 19956 3676 20012
rect 3676 19956 3732 20012
rect 3732 19956 3736 20012
rect 3672 19952 3736 19956
rect 3752 20012 3816 20016
rect 3752 19956 3756 20012
rect 3756 19956 3812 20012
rect 3812 19956 3816 20012
rect 3752 19952 3816 19956
rect 18872 19468 18936 19472
rect 18872 19412 18876 19468
rect 18876 19412 18932 19468
rect 18932 19412 18936 19468
rect 18872 19408 18936 19412
rect 18952 19468 19016 19472
rect 18952 19412 18956 19468
rect 18956 19412 19012 19468
rect 19012 19412 19016 19468
rect 18952 19408 19016 19412
rect 19032 19468 19096 19472
rect 19032 19412 19036 19468
rect 19036 19412 19092 19468
rect 19092 19412 19096 19468
rect 19032 19408 19096 19412
rect 19112 19468 19176 19472
rect 19112 19412 19116 19468
rect 19116 19412 19172 19468
rect 19172 19412 19176 19468
rect 19112 19408 19176 19412
rect 3512 18924 3576 18928
rect 3512 18868 3516 18924
rect 3516 18868 3572 18924
rect 3572 18868 3576 18924
rect 3512 18864 3576 18868
rect 3592 18924 3656 18928
rect 3592 18868 3596 18924
rect 3596 18868 3652 18924
rect 3652 18868 3656 18924
rect 3592 18864 3656 18868
rect 3672 18924 3736 18928
rect 3672 18868 3676 18924
rect 3676 18868 3732 18924
rect 3732 18868 3736 18924
rect 3672 18864 3736 18868
rect 3752 18924 3816 18928
rect 3752 18868 3756 18924
rect 3756 18868 3812 18924
rect 3812 18868 3816 18924
rect 3752 18864 3816 18868
rect 18872 18380 18936 18384
rect 18872 18324 18876 18380
rect 18876 18324 18932 18380
rect 18932 18324 18936 18380
rect 18872 18320 18936 18324
rect 18952 18380 19016 18384
rect 18952 18324 18956 18380
rect 18956 18324 19012 18380
rect 19012 18324 19016 18380
rect 18952 18320 19016 18324
rect 19032 18380 19096 18384
rect 19032 18324 19036 18380
rect 19036 18324 19092 18380
rect 19092 18324 19096 18380
rect 19032 18320 19096 18324
rect 19112 18380 19176 18384
rect 19112 18324 19116 18380
rect 19116 18324 19172 18380
rect 19172 18324 19176 18380
rect 19112 18320 19176 18324
rect 3512 17836 3576 17840
rect 3512 17780 3516 17836
rect 3516 17780 3572 17836
rect 3572 17780 3576 17836
rect 3512 17776 3576 17780
rect 3592 17836 3656 17840
rect 3592 17780 3596 17836
rect 3596 17780 3652 17836
rect 3652 17780 3656 17836
rect 3592 17776 3656 17780
rect 3672 17836 3736 17840
rect 3672 17780 3676 17836
rect 3676 17780 3732 17836
rect 3732 17780 3736 17836
rect 3672 17776 3736 17780
rect 3752 17836 3816 17840
rect 3752 17780 3756 17836
rect 3756 17780 3812 17836
rect 3812 17780 3816 17836
rect 3752 17776 3816 17780
rect 18872 17292 18936 17296
rect 18872 17236 18876 17292
rect 18876 17236 18932 17292
rect 18932 17236 18936 17292
rect 18872 17232 18936 17236
rect 18952 17292 19016 17296
rect 18952 17236 18956 17292
rect 18956 17236 19012 17292
rect 19012 17236 19016 17292
rect 18952 17232 19016 17236
rect 19032 17292 19096 17296
rect 19032 17236 19036 17292
rect 19036 17236 19092 17292
rect 19092 17236 19096 17292
rect 19032 17232 19096 17236
rect 19112 17292 19176 17296
rect 19112 17236 19116 17292
rect 19116 17236 19172 17292
rect 19172 17236 19176 17292
rect 19112 17232 19176 17236
rect 3512 16748 3576 16752
rect 3512 16692 3516 16748
rect 3516 16692 3572 16748
rect 3572 16692 3576 16748
rect 3512 16688 3576 16692
rect 3592 16748 3656 16752
rect 3592 16692 3596 16748
rect 3596 16692 3652 16748
rect 3652 16692 3656 16748
rect 3592 16688 3656 16692
rect 3672 16748 3736 16752
rect 3672 16692 3676 16748
rect 3676 16692 3732 16748
rect 3732 16692 3736 16748
rect 3672 16688 3736 16692
rect 3752 16748 3816 16752
rect 3752 16692 3756 16748
rect 3756 16692 3812 16748
rect 3812 16692 3816 16748
rect 3752 16688 3816 16692
rect 18872 16204 18936 16208
rect 18872 16148 18876 16204
rect 18876 16148 18932 16204
rect 18932 16148 18936 16204
rect 18872 16144 18936 16148
rect 18952 16204 19016 16208
rect 18952 16148 18956 16204
rect 18956 16148 19012 16204
rect 19012 16148 19016 16204
rect 18952 16144 19016 16148
rect 19032 16204 19096 16208
rect 19032 16148 19036 16204
rect 19036 16148 19092 16204
rect 19092 16148 19096 16204
rect 19032 16144 19096 16148
rect 19112 16204 19176 16208
rect 19112 16148 19116 16204
rect 19116 16148 19172 16204
rect 19172 16148 19176 16204
rect 19112 16144 19176 16148
rect 3512 15660 3576 15664
rect 3512 15604 3516 15660
rect 3516 15604 3572 15660
rect 3572 15604 3576 15660
rect 3512 15600 3576 15604
rect 3592 15660 3656 15664
rect 3592 15604 3596 15660
rect 3596 15604 3652 15660
rect 3652 15604 3656 15660
rect 3592 15600 3656 15604
rect 3672 15660 3736 15664
rect 3672 15604 3676 15660
rect 3676 15604 3732 15660
rect 3732 15604 3736 15660
rect 3672 15600 3736 15604
rect 3752 15660 3816 15664
rect 3752 15604 3756 15660
rect 3756 15604 3812 15660
rect 3812 15604 3816 15660
rect 3752 15600 3816 15604
rect 18872 15116 18936 15120
rect 18872 15060 18876 15116
rect 18876 15060 18932 15116
rect 18932 15060 18936 15116
rect 18872 15056 18936 15060
rect 18952 15116 19016 15120
rect 18952 15060 18956 15116
rect 18956 15060 19012 15116
rect 19012 15060 19016 15116
rect 18952 15056 19016 15060
rect 19032 15116 19096 15120
rect 19032 15060 19036 15116
rect 19036 15060 19092 15116
rect 19092 15060 19096 15116
rect 19032 15056 19096 15060
rect 19112 15116 19176 15120
rect 19112 15060 19116 15116
rect 19116 15060 19172 15116
rect 19172 15060 19176 15116
rect 19112 15056 19176 15060
rect 3512 14572 3576 14576
rect 3512 14516 3516 14572
rect 3516 14516 3572 14572
rect 3572 14516 3576 14572
rect 3512 14512 3576 14516
rect 3592 14572 3656 14576
rect 3592 14516 3596 14572
rect 3596 14516 3652 14572
rect 3652 14516 3656 14572
rect 3592 14512 3656 14516
rect 3672 14572 3736 14576
rect 3672 14516 3676 14572
rect 3676 14516 3732 14572
rect 3732 14516 3736 14572
rect 3672 14512 3736 14516
rect 3752 14572 3816 14576
rect 3752 14516 3756 14572
rect 3756 14516 3812 14572
rect 3812 14516 3816 14572
rect 3752 14512 3816 14516
rect 18872 14028 18936 14032
rect 18872 13972 18876 14028
rect 18876 13972 18932 14028
rect 18932 13972 18936 14028
rect 18872 13968 18936 13972
rect 18952 14028 19016 14032
rect 18952 13972 18956 14028
rect 18956 13972 19012 14028
rect 19012 13972 19016 14028
rect 18952 13968 19016 13972
rect 19032 14028 19096 14032
rect 19032 13972 19036 14028
rect 19036 13972 19092 14028
rect 19092 13972 19096 14028
rect 19032 13968 19096 13972
rect 19112 14028 19176 14032
rect 19112 13972 19116 14028
rect 19116 13972 19172 14028
rect 19172 13972 19176 14028
rect 19112 13968 19176 13972
rect 3512 13484 3576 13488
rect 3512 13428 3516 13484
rect 3516 13428 3572 13484
rect 3572 13428 3576 13484
rect 3512 13424 3576 13428
rect 3592 13484 3656 13488
rect 3592 13428 3596 13484
rect 3596 13428 3652 13484
rect 3652 13428 3656 13484
rect 3592 13424 3656 13428
rect 3672 13484 3736 13488
rect 3672 13428 3676 13484
rect 3676 13428 3732 13484
rect 3732 13428 3736 13484
rect 3672 13424 3736 13428
rect 3752 13484 3816 13488
rect 3752 13428 3756 13484
rect 3756 13428 3812 13484
rect 3812 13428 3816 13484
rect 3752 13424 3816 13428
rect 18872 12940 18936 12944
rect 18872 12884 18876 12940
rect 18876 12884 18932 12940
rect 18932 12884 18936 12940
rect 18872 12880 18936 12884
rect 18952 12940 19016 12944
rect 18952 12884 18956 12940
rect 18956 12884 19012 12940
rect 19012 12884 19016 12940
rect 18952 12880 19016 12884
rect 19032 12940 19096 12944
rect 19032 12884 19036 12940
rect 19036 12884 19092 12940
rect 19092 12884 19096 12940
rect 19032 12880 19096 12884
rect 19112 12940 19176 12944
rect 19112 12884 19116 12940
rect 19116 12884 19172 12940
rect 19172 12884 19176 12940
rect 19112 12880 19176 12884
rect 3512 12396 3576 12400
rect 3512 12340 3516 12396
rect 3516 12340 3572 12396
rect 3572 12340 3576 12396
rect 3512 12336 3576 12340
rect 3592 12396 3656 12400
rect 3592 12340 3596 12396
rect 3596 12340 3652 12396
rect 3652 12340 3656 12396
rect 3592 12336 3656 12340
rect 3672 12396 3736 12400
rect 3672 12340 3676 12396
rect 3676 12340 3732 12396
rect 3732 12340 3736 12396
rect 3672 12336 3736 12340
rect 3752 12396 3816 12400
rect 3752 12340 3756 12396
rect 3756 12340 3812 12396
rect 3812 12340 3816 12396
rect 3752 12336 3816 12340
rect 18872 11852 18936 11856
rect 18872 11796 18876 11852
rect 18876 11796 18932 11852
rect 18932 11796 18936 11852
rect 18872 11792 18936 11796
rect 18952 11852 19016 11856
rect 18952 11796 18956 11852
rect 18956 11796 19012 11852
rect 19012 11796 19016 11852
rect 18952 11792 19016 11796
rect 19032 11852 19096 11856
rect 19032 11796 19036 11852
rect 19036 11796 19092 11852
rect 19092 11796 19096 11852
rect 19032 11792 19096 11796
rect 19112 11852 19176 11856
rect 19112 11796 19116 11852
rect 19116 11796 19172 11852
rect 19172 11796 19176 11852
rect 19112 11792 19176 11796
rect 3512 11308 3576 11312
rect 3512 11252 3516 11308
rect 3516 11252 3572 11308
rect 3572 11252 3576 11308
rect 3512 11248 3576 11252
rect 3592 11308 3656 11312
rect 3592 11252 3596 11308
rect 3596 11252 3652 11308
rect 3652 11252 3656 11308
rect 3592 11248 3656 11252
rect 3672 11308 3736 11312
rect 3672 11252 3676 11308
rect 3676 11252 3732 11308
rect 3732 11252 3736 11308
rect 3672 11248 3736 11252
rect 3752 11308 3816 11312
rect 3752 11252 3756 11308
rect 3756 11252 3812 11308
rect 3812 11252 3816 11308
rect 3752 11248 3816 11252
rect 18872 10764 18936 10768
rect 18872 10708 18876 10764
rect 18876 10708 18932 10764
rect 18932 10708 18936 10764
rect 18872 10704 18936 10708
rect 18952 10764 19016 10768
rect 18952 10708 18956 10764
rect 18956 10708 19012 10764
rect 19012 10708 19016 10764
rect 18952 10704 19016 10708
rect 19032 10764 19096 10768
rect 19032 10708 19036 10764
rect 19036 10708 19092 10764
rect 19092 10708 19096 10764
rect 19032 10704 19096 10708
rect 19112 10764 19176 10768
rect 19112 10708 19116 10764
rect 19116 10708 19172 10764
rect 19172 10708 19176 10764
rect 19112 10704 19176 10708
rect 3512 10220 3576 10224
rect 3512 10164 3516 10220
rect 3516 10164 3572 10220
rect 3572 10164 3576 10220
rect 3512 10160 3576 10164
rect 3592 10220 3656 10224
rect 3592 10164 3596 10220
rect 3596 10164 3652 10220
rect 3652 10164 3656 10220
rect 3592 10160 3656 10164
rect 3672 10220 3736 10224
rect 3672 10164 3676 10220
rect 3676 10164 3732 10220
rect 3732 10164 3736 10220
rect 3672 10160 3736 10164
rect 3752 10220 3816 10224
rect 3752 10164 3756 10220
rect 3756 10164 3812 10220
rect 3812 10164 3816 10220
rect 3752 10160 3816 10164
rect 18872 9676 18936 9680
rect 18872 9620 18876 9676
rect 18876 9620 18932 9676
rect 18932 9620 18936 9676
rect 18872 9616 18936 9620
rect 18952 9676 19016 9680
rect 18952 9620 18956 9676
rect 18956 9620 19012 9676
rect 19012 9620 19016 9676
rect 18952 9616 19016 9620
rect 19032 9676 19096 9680
rect 19032 9620 19036 9676
rect 19036 9620 19092 9676
rect 19092 9620 19096 9676
rect 19032 9616 19096 9620
rect 19112 9676 19176 9680
rect 19112 9620 19116 9676
rect 19116 9620 19172 9676
rect 19172 9620 19176 9676
rect 19112 9616 19176 9620
rect 3512 9132 3576 9136
rect 3512 9076 3516 9132
rect 3516 9076 3572 9132
rect 3572 9076 3576 9132
rect 3512 9072 3576 9076
rect 3592 9132 3656 9136
rect 3592 9076 3596 9132
rect 3596 9076 3652 9132
rect 3652 9076 3656 9132
rect 3592 9072 3656 9076
rect 3672 9132 3736 9136
rect 3672 9076 3676 9132
rect 3676 9076 3732 9132
rect 3732 9076 3736 9132
rect 3672 9072 3736 9076
rect 3752 9132 3816 9136
rect 3752 9076 3756 9132
rect 3756 9076 3812 9132
rect 3812 9076 3816 9132
rect 3752 9072 3816 9076
rect 18872 8588 18936 8592
rect 18872 8532 18876 8588
rect 18876 8532 18932 8588
rect 18932 8532 18936 8588
rect 18872 8528 18936 8532
rect 18952 8588 19016 8592
rect 18952 8532 18956 8588
rect 18956 8532 19012 8588
rect 19012 8532 19016 8588
rect 18952 8528 19016 8532
rect 19032 8588 19096 8592
rect 19032 8532 19036 8588
rect 19036 8532 19092 8588
rect 19092 8532 19096 8588
rect 19032 8528 19096 8532
rect 19112 8588 19176 8592
rect 19112 8532 19116 8588
rect 19116 8532 19172 8588
rect 19172 8532 19176 8588
rect 19112 8528 19176 8532
rect 3512 8044 3576 8048
rect 3512 7988 3516 8044
rect 3516 7988 3572 8044
rect 3572 7988 3576 8044
rect 3512 7984 3576 7988
rect 3592 8044 3656 8048
rect 3592 7988 3596 8044
rect 3596 7988 3652 8044
rect 3652 7988 3656 8044
rect 3592 7984 3656 7988
rect 3672 8044 3736 8048
rect 3672 7988 3676 8044
rect 3676 7988 3732 8044
rect 3732 7988 3736 8044
rect 3672 7984 3736 7988
rect 3752 8044 3816 8048
rect 3752 7988 3756 8044
rect 3756 7988 3812 8044
rect 3812 7988 3816 8044
rect 3752 7984 3816 7988
rect 18872 7500 18936 7504
rect 18872 7444 18876 7500
rect 18876 7444 18932 7500
rect 18932 7444 18936 7500
rect 18872 7440 18936 7444
rect 18952 7500 19016 7504
rect 18952 7444 18956 7500
rect 18956 7444 19012 7500
rect 19012 7444 19016 7500
rect 18952 7440 19016 7444
rect 19032 7500 19096 7504
rect 19032 7444 19036 7500
rect 19036 7444 19092 7500
rect 19092 7444 19096 7500
rect 19032 7440 19096 7444
rect 19112 7500 19176 7504
rect 19112 7444 19116 7500
rect 19116 7444 19172 7500
rect 19172 7444 19176 7500
rect 19112 7440 19176 7444
rect 3512 6956 3576 6960
rect 3512 6900 3516 6956
rect 3516 6900 3572 6956
rect 3572 6900 3576 6956
rect 3512 6896 3576 6900
rect 3592 6956 3656 6960
rect 3592 6900 3596 6956
rect 3596 6900 3652 6956
rect 3652 6900 3656 6956
rect 3592 6896 3656 6900
rect 3672 6956 3736 6960
rect 3672 6900 3676 6956
rect 3676 6900 3732 6956
rect 3732 6900 3736 6956
rect 3672 6896 3736 6900
rect 3752 6956 3816 6960
rect 3752 6900 3756 6956
rect 3756 6900 3812 6956
rect 3812 6900 3816 6956
rect 3752 6896 3816 6900
rect 18872 6412 18936 6416
rect 18872 6356 18876 6412
rect 18876 6356 18932 6412
rect 18932 6356 18936 6412
rect 18872 6352 18936 6356
rect 18952 6412 19016 6416
rect 18952 6356 18956 6412
rect 18956 6356 19012 6412
rect 19012 6356 19016 6412
rect 18952 6352 19016 6356
rect 19032 6412 19096 6416
rect 19032 6356 19036 6412
rect 19036 6356 19092 6412
rect 19092 6356 19096 6412
rect 19032 6352 19096 6356
rect 19112 6412 19176 6416
rect 19112 6356 19116 6412
rect 19116 6356 19172 6412
rect 19172 6356 19176 6412
rect 19112 6352 19176 6356
rect 3512 5868 3576 5872
rect 3512 5812 3516 5868
rect 3516 5812 3572 5868
rect 3572 5812 3576 5868
rect 3512 5808 3576 5812
rect 3592 5868 3656 5872
rect 3592 5812 3596 5868
rect 3596 5812 3652 5868
rect 3652 5812 3656 5868
rect 3592 5808 3656 5812
rect 3672 5868 3736 5872
rect 3672 5812 3676 5868
rect 3676 5812 3732 5868
rect 3732 5812 3736 5868
rect 3672 5808 3736 5812
rect 3752 5868 3816 5872
rect 3752 5812 3756 5868
rect 3756 5812 3812 5868
rect 3812 5812 3816 5868
rect 3752 5808 3816 5812
rect 18872 5324 18936 5328
rect 18872 5268 18876 5324
rect 18876 5268 18932 5324
rect 18932 5268 18936 5324
rect 18872 5264 18936 5268
rect 18952 5324 19016 5328
rect 18952 5268 18956 5324
rect 18956 5268 19012 5324
rect 19012 5268 19016 5324
rect 18952 5264 19016 5268
rect 19032 5324 19096 5328
rect 19032 5268 19036 5324
rect 19036 5268 19092 5324
rect 19092 5268 19096 5324
rect 19032 5264 19096 5268
rect 19112 5324 19176 5328
rect 19112 5268 19116 5324
rect 19116 5268 19172 5324
rect 19172 5268 19176 5324
rect 19112 5264 19176 5268
rect 3512 4780 3576 4784
rect 3512 4724 3516 4780
rect 3516 4724 3572 4780
rect 3572 4724 3576 4780
rect 3512 4720 3576 4724
rect 3592 4780 3656 4784
rect 3592 4724 3596 4780
rect 3596 4724 3652 4780
rect 3652 4724 3656 4780
rect 3592 4720 3656 4724
rect 3672 4780 3736 4784
rect 3672 4724 3676 4780
rect 3676 4724 3732 4780
rect 3732 4724 3736 4780
rect 3672 4720 3736 4724
rect 3752 4780 3816 4784
rect 3752 4724 3756 4780
rect 3756 4724 3812 4780
rect 3812 4724 3816 4780
rect 3752 4720 3816 4724
rect 18872 4236 18936 4240
rect 18872 4180 18876 4236
rect 18876 4180 18932 4236
rect 18932 4180 18936 4236
rect 18872 4176 18936 4180
rect 18952 4236 19016 4240
rect 18952 4180 18956 4236
rect 18956 4180 19012 4236
rect 19012 4180 19016 4236
rect 18952 4176 19016 4180
rect 19032 4236 19096 4240
rect 19032 4180 19036 4236
rect 19036 4180 19092 4236
rect 19092 4180 19096 4236
rect 19032 4176 19096 4180
rect 19112 4236 19176 4240
rect 19112 4180 19116 4236
rect 19116 4180 19172 4236
rect 19172 4180 19176 4236
rect 19112 4176 19176 4180
rect 3512 3692 3576 3696
rect 3512 3636 3516 3692
rect 3516 3636 3572 3692
rect 3572 3636 3576 3692
rect 3512 3632 3576 3636
rect 3592 3692 3656 3696
rect 3592 3636 3596 3692
rect 3596 3636 3652 3692
rect 3652 3636 3656 3692
rect 3592 3632 3656 3636
rect 3672 3692 3736 3696
rect 3672 3636 3676 3692
rect 3676 3636 3732 3692
rect 3732 3636 3736 3692
rect 3672 3632 3736 3636
rect 3752 3692 3816 3696
rect 3752 3636 3756 3692
rect 3756 3636 3812 3692
rect 3812 3636 3816 3692
rect 3752 3632 3816 3636
rect 18872 3148 18936 3152
rect 18872 3092 18876 3148
rect 18876 3092 18932 3148
rect 18932 3092 18936 3148
rect 18872 3088 18936 3092
rect 18952 3148 19016 3152
rect 18952 3092 18956 3148
rect 18956 3092 19012 3148
rect 19012 3092 19016 3148
rect 18952 3088 19016 3092
rect 19032 3148 19096 3152
rect 19032 3092 19036 3148
rect 19036 3092 19092 3148
rect 19092 3092 19096 3148
rect 19032 3088 19096 3092
rect 19112 3148 19176 3152
rect 19112 3092 19116 3148
rect 19116 3092 19172 3148
rect 19172 3092 19176 3148
rect 19112 3088 19176 3092
rect 3512 2604 3576 2608
rect 3512 2548 3516 2604
rect 3516 2548 3572 2604
rect 3572 2548 3576 2604
rect 3512 2544 3576 2548
rect 3592 2604 3656 2608
rect 3592 2548 3596 2604
rect 3596 2548 3652 2604
rect 3652 2548 3656 2604
rect 3592 2544 3656 2548
rect 3672 2604 3736 2608
rect 3672 2548 3676 2604
rect 3676 2548 3732 2604
rect 3732 2548 3736 2604
rect 3672 2544 3736 2548
rect 3752 2604 3816 2608
rect 3752 2548 3756 2604
rect 3756 2548 3812 2604
rect 3812 2548 3816 2604
rect 3752 2544 3816 2548
rect 18872 2060 18936 2064
rect 18872 2004 18876 2060
rect 18876 2004 18932 2060
rect 18932 2004 18936 2060
rect 18872 2000 18936 2004
rect 18952 2060 19016 2064
rect 18952 2004 18956 2060
rect 18956 2004 19012 2060
rect 19012 2004 19016 2060
rect 18952 2000 19016 2004
rect 19032 2060 19096 2064
rect 19032 2004 19036 2060
rect 19036 2004 19092 2060
rect 19092 2004 19096 2060
rect 19032 2000 19096 2004
rect 19112 2060 19176 2064
rect 19112 2004 19116 2060
rect 19116 2004 19172 2060
rect 19172 2004 19176 2060
rect 19112 2000 19176 2004
rect 3512 1516 3576 1520
rect 3512 1460 3516 1516
rect 3516 1460 3572 1516
rect 3572 1460 3576 1516
rect 3512 1456 3576 1460
rect 3592 1516 3656 1520
rect 3592 1460 3596 1516
rect 3596 1460 3652 1516
rect 3652 1460 3656 1516
rect 3592 1456 3656 1460
rect 3672 1516 3736 1520
rect 3672 1460 3676 1516
rect 3676 1460 3732 1516
rect 3732 1460 3736 1516
rect 3672 1456 3736 1460
rect 3752 1516 3816 1520
rect 3752 1460 3756 1516
rect 3756 1460 3812 1516
rect 3812 1460 3816 1516
rect 3752 1456 3816 1460
rect 18872 972 18936 976
rect 18872 916 18876 972
rect 18876 916 18932 972
rect 18932 916 18936 972
rect 18872 912 18936 916
rect 18952 972 19016 976
rect 18952 916 18956 972
rect 18956 916 19012 972
rect 19012 916 19016 972
rect 18952 912 19016 916
rect 19032 972 19096 976
rect 19032 916 19036 972
rect 19036 916 19092 972
rect 19092 916 19096 972
rect 19032 912 19096 916
rect 19112 972 19176 976
rect 19112 916 19116 972
rect 19116 916 19172 972
rect 19172 916 19176 972
rect 19112 912 19176 916
rect 3512 428 3576 432
rect 3512 372 3516 428
rect 3516 372 3572 428
rect 3572 372 3576 428
rect 3512 368 3576 372
rect 3592 428 3656 432
rect 3592 372 3596 428
rect 3596 372 3652 428
rect 3652 372 3656 428
rect 3592 368 3656 372
rect 3672 428 3736 432
rect 3672 372 3676 428
rect 3676 372 3732 428
rect 3732 372 3736 428
rect 3672 368 3736 372
rect 3752 428 3816 432
rect 3752 372 3756 428
rect 3756 372 3812 428
rect 3812 372 3816 428
rect 3752 368 3816 372
<< metal4 >>
rect 18864 27088 19184 27104
rect 3504 26544 3824 27056
rect 3504 26480 3512 26544
rect 3576 26480 3592 26544
rect 3656 26480 3672 26544
rect 3736 26480 3752 26544
rect 3816 26480 3824 26544
rect 3504 25456 3824 26480
rect 3504 25392 3512 25456
rect 3576 25392 3592 25456
rect 3656 25392 3672 25456
rect 3736 25392 3752 25456
rect 3816 25392 3824 25456
rect 3504 24368 3824 25392
rect 3504 24304 3512 24368
rect 3576 24304 3592 24368
rect 3656 24304 3672 24368
rect 3736 24304 3752 24368
rect 3816 24304 3824 24368
rect 3504 23280 3824 24304
rect 3504 23216 3512 23280
rect 3576 23216 3592 23280
rect 3656 23216 3672 23280
rect 3736 23216 3752 23280
rect 3816 23216 3824 23280
rect 3504 22192 3824 23216
rect 3504 22128 3512 22192
rect 3576 22128 3592 22192
rect 3656 22128 3672 22192
rect 3736 22128 3752 22192
rect 3816 22128 3824 22192
rect 3504 21104 3824 22128
rect 3504 21040 3512 21104
rect 3576 21040 3592 21104
rect 3656 21040 3672 21104
rect 3736 21040 3752 21104
rect 3816 21040 3824 21104
rect 3504 20016 3824 21040
rect 3504 19952 3512 20016
rect 3576 19952 3592 20016
rect 3656 19952 3672 20016
rect 3736 19952 3752 20016
rect 3816 19952 3824 20016
rect 3504 18928 3824 19952
rect 3504 18864 3512 18928
rect 3576 18864 3592 18928
rect 3656 18864 3672 18928
rect 3736 18864 3752 18928
rect 3816 18864 3824 18928
rect 3504 17840 3824 18864
rect 3504 17776 3512 17840
rect 3576 17776 3592 17840
rect 3656 17776 3672 17840
rect 3736 17776 3752 17840
rect 3816 17776 3824 17840
rect 3504 16752 3824 17776
rect 3504 16688 3512 16752
rect 3576 16688 3592 16752
rect 3656 16688 3672 16752
rect 3736 16688 3752 16752
rect 3816 16688 3824 16752
rect 3504 15664 3824 16688
rect 3504 15600 3512 15664
rect 3576 15600 3592 15664
rect 3656 15600 3672 15664
rect 3736 15600 3752 15664
rect 3816 15600 3824 15664
rect 3504 14576 3824 15600
rect 3504 14512 3512 14576
rect 3576 14512 3592 14576
rect 3656 14512 3672 14576
rect 3736 14512 3752 14576
rect 3816 14512 3824 14576
rect 3504 13488 3824 14512
rect 3504 13424 3512 13488
rect 3576 13424 3592 13488
rect 3656 13424 3672 13488
rect 3736 13424 3752 13488
rect 3816 13424 3824 13488
rect 3504 12400 3824 13424
rect 3504 12336 3512 12400
rect 3576 12336 3592 12400
rect 3656 12336 3672 12400
rect 3736 12336 3752 12400
rect 3816 12336 3824 12400
rect 3504 11312 3824 12336
rect 3504 11248 3512 11312
rect 3576 11248 3592 11312
rect 3656 11248 3672 11312
rect 3736 11248 3752 11312
rect 3816 11248 3824 11312
rect 3504 10224 3824 11248
rect 3504 10160 3512 10224
rect 3576 10160 3592 10224
rect 3656 10160 3672 10224
rect 3736 10160 3752 10224
rect 3816 10160 3824 10224
rect 3504 9136 3824 10160
rect 3504 9072 3512 9136
rect 3576 9072 3592 9136
rect 3656 9072 3672 9136
rect 3736 9072 3752 9136
rect 3816 9072 3824 9136
rect 3504 8048 3824 9072
rect 3504 7984 3512 8048
rect 3576 7984 3592 8048
rect 3656 7984 3672 8048
rect 3736 7984 3752 8048
rect 3816 7984 3824 8048
rect 3504 6960 3824 7984
rect 3504 6896 3512 6960
rect 3576 6896 3592 6960
rect 3656 6896 3672 6960
rect 3736 6896 3752 6960
rect 3816 6896 3824 6960
rect 3504 5872 3824 6896
rect 3504 5808 3512 5872
rect 3576 5808 3592 5872
rect 3656 5808 3672 5872
rect 3736 5808 3752 5872
rect 3816 5808 3824 5872
rect 3504 4784 3824 5808
rect 3504 4720 3512 4784
rect 3576 4720 3592 4784
rect 3656 4720 3672 4784
rect 3736 4720 3752 4784
rect 3816 4720 3824 4784
rect 3504 3848 3824 4720
rect 3504 3696 3546 3848
rect 3782 3696 3824 3848
rect 3504 3632 3512 3696
rect 3816 3632 3824 3696
rect 3504 3612 3546 3632
rect 3782 3612 3824 3632
rect 3504 2608 3824 3612
rect 3504 2544 3512 2608
rect 3576 2544 3592 2608
rect 3656 2544 3672 2608
rect 3736 2544 3752 2608
rect 3816 2544 3824 2608
rect 3504 1520 3824 2544
rect 3504 1456 3512 1520
rect 3576 1456 3592 1520
rect 3656 1456 3672 1520
rect 3736 1456 3752 1520
rect 3816 1456 3824 1520
rect 3504 432 3824 1456
rect 3504 368 3512 432
rect 3576 368 3592 432
rect 3656 368 3672 432
rect 3736 368 3752 432
rect 3816 368 3824 432
rect 18864 27024 18872 27088
rect 18936 27024 18952 27088
rect 19016 27024 19032 27088
rect 19096 27024 19112 27088
rect 19176 27024 19184 27088
rect 18864 26000 19184 27024
rect 18864 25936 18872 26000
rect 18936 25936 18952 26000
rect 19016 25936 19032 26000
rect 19096 25936 19112 26000
rect 19176 25936 19184 26000
rect 18864 24912 19184 25936
rect 18864 24848 18872 24912
rect 18936 24848 18952 24912
rect 19016 24848 19032 24912
rect 19096 24848 19112 24912
rect 19176 24848 19184 24912
rect 18864 23824 19184 24848
rect 18864 23760 18872 23824
rect 18936 23760 18952 23824
rect 19016 23760 19032 23824
rect 19096 23760 19112 23824
rect 19176 23760 19184 23824
rect 18864 22736 19184 23760
rect 18864 22672 18872 22736
rect 18936 22672 18952 22736
rect 19016 22672 19032 22736
rect 19096 22672 19112 22736
rect 19176 22672 19184 22736
rect 18864 21648 19184 22672
rect 18864 21584 18872 21648
rect 18936 21584 18952 21648
rect 19016 21584 19032 21648
rect 19096 21584 19112 21648
rect 19176 21584 19184 21648
rect 18864 20560 19184 21584
rect 18864 20496 18872 20560
rect 18936 20496 18952 20560
rect 19016 20496 19032 20560
rect 19096 20496 19112 20560
rect 19176 20496 19184 20560
rect 18864 19472 19184 20496
rect 18864 19408 18872 19472
rect 18936 19408 18952 19472
rect 19016 19408 19032 19472
rect 19096 19408 19112 19472
rect 19176 19408 19184 19472
rect 18864 19166 19184 19408
rect 18864 18930 18906 19166
rect 19142 18930 19184 19166
rect 18864 18384 19184 18930
rect 18864 18320 18872 18384
rect 18936 18320 18952 18384
rect 19016 18320 19032 18384
rect 19096 18320 19112 18384
rect 19176 18320 19184 18384
rect 18864 17296 19184 18320
rect 18864 17232 18872 17296
rect 18936 17232 18952 17296
rect 19016 17232 19032 17296
rect 19096 17232 19112 17296
rect 19176 17232 19184 17296
rect 18864 16208 19184 17232
rect 18864 16144 18872 16208
rect 18936 16144 18952 16208
rect 19016 16144 19032 16208
rect 19096 16144 19112 16208
rect 19176 16144 19184 16208
rect 18864 15120 19184 16144
rect 18864 15056 18872 15120
rect 18936 15056 18952 15120
rect 19016 15056 19032 15120
rect 19096 15056 19112 15120
rect 19176 15056 19184 15120
rect 18864 14032 19184 15056
rect 18864 13968 18872 14032
rect 18936 13968 18952 14032
rect 19016 13968 19032 14032
rect 19096 13968 19112 14032
rect 19176 13968 19184 14032
rect 18864 12944 19184 13968
rect 18864 12880 18872 12944
rect 18936 12880 18952 12944
rect 19016 12880 19032 12944
rect 19096 12880 19112 12944
rect 19176 12880 19184 12944
rect 18864 11856 19184 12880
rect 18864 11792 18872 11856
rect 18936 11792 18952 11856
rect 19016 11792 19032 11856
rect 19096 11792 19112 11856
rect 19176 11792 19184 11856
rect 18864 10768 19184 11792
rect 18864 10704 18872 10768
rect 18936 10704 18952 10768
rect 19016 10704 19032 10768
rect 19096 10704 19112 10768
rect 19176 10704 19184 10768
rect 18864 9680 19184 10704
rect 18864 9616 18872 9680
rect 18936 9616 18952 9680
rect 19016 9616 19032 9680
rect 19096 9616 19112 9680
rect 19176 9616 19184 9680
rect 18864 8592 19184 9616
rect 18864 8528 18872 8592
rect 18936 8528 18952 8592
rect 19016 8528 19032 8592
rect 19096 8528 19112 8592
rect 19176 8528 19184 8592
rect 18864 7504 19184 8528
rect 18864 7440 18872 7504
rect 18936 7440 18952 7504
rect 19016 7440 19032 7504
rect 19096 7440 19112 7504
rect 19176 7440 19184 7504
rect 18864 6416 19184 7440
rect 18864 6352 18872 6416
rect 18936 6352 18952 6416
rect 19016 6352 19032 6416
rect 19096 6352 19112 6416
rect 19176 6352 19184 6416
rect 18864 5328 19184 6352
rect 18864 5264 18872 5328
rect 18936 5264 18952 5328
rect 19016 5264 19032 5328
rect 19096 5264 19112 5328
rect 19176 5264 19184 5328
rect 18864 4240 19184 5264
rect 18864 4176 18872 4240
rect 18936 4176 18952 4240
rect 19016 4176 19032 4240
rect 19096 4176 19112 4240
rect 19176 4176 19184 4240
rect 18864 3152 19184 4176
rect 18864 3088 18872 3152
rect 18936 3088 18952 3152
rect 19016 3088 19032 3152
rect 19096 3088 19112 3152
rect 19176 3088 19184 3152
rect 18864 2064 19184 3088
rect 18864 2000 18872 2064
rect 18936 2000 18952 2064
rect 19016 2000 19032 2064
rect 19096 2000 19112 2064
rect 19176 2000 19184 2064
rect 18864 976 19184 2000
rect 18864 912 18872 976
rect 18936 912 18952 976
rect 19016 912 19032 976
rect 19096 912 19112 976
rect 19176 912 19184 976
rect 18864 400 19184 912
rect 3504 352 3824 368
<< via4 >>
rect 3546 3696 3782 3848
rect 3546 3632 3576 3696
rect 3576 3632 3592 3696
rect 3592 3632 3656 3696
rect 3656 3632 3672 3696
rect 3672 3632 3736 3696
rect 3736 3632 3752 3696
rect 3752 3632 3782 3696
rect 3546 3612 3782 3632
rect 18906 18930 19142 19166
<< metal5 >>
rect 400 19166 27264 19208
rect 400 18930 18906 19166
rect 19142 18930 27264 19166
rect 400 18888 27264 18930
rect 400 3848 27264 3890
rect 400 3612 3546 3848
rect 3782 3612 27264 3848
rect 400 3570 27264 3612
use sky130_fd_sc_hd__decap_3  PHY_2 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 400 0 1 944
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1586547711
transform 1 0 400 0 -1 944
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL1380x2720 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 676 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1313 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 768 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL4140x0
timestamp 1586547711
transform 1 0 1228 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_976
timestamp 1586547711
transform 1 0 952 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_611
timestamp 1586547711
transform 1 0 1136 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_977
timestamp 1586547711
transform 1 0 1320 0 -1 944
box 0 -48 184 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen1 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 1320 0 1 944
box 0 -48 644 592
use sky130_fd_sc_hd__decap_6  FILL1380x0 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 676 0 -1 944
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_62
timestamp 1586547711
transform 1 0 1964 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_73
timestamp 1586547711
transform 1 0 2148 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1314
timestamp 1586547711
transform 1 0 1504 0 -1 944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL9660x2720
timestamp 1586547711
transform 1 0 2332 0 1 944
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL6440x0 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 1688 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL14720x0
timestamp 1586547711
transform 1 0 3344 0 -1 944
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL12420x2720
timestamp 1586547711
transform 1 0 2884 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL13800x0
timestamp 1586547711
transform 1 0 3160 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_936
timestamp 1586547711
transform 1 0 2976 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 3252 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL11960x0 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 2792 0 -1 944
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _287_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 3160 0 1 944
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1586547711
transform 1 0 3804 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1586547711
transform 1 0 3988 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_61
timestamp 1586547711
transform 1 0 4172 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_74
timestamp 1586547711
transform 1 0 4356 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_600
timestamp 1586547711
transform 1 0 3620 0 -1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_970
timestamp 1586547711
transform 1 0 3804 0 -1 944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL20700x2720 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 4540 0 1 944
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILL17940x0
timestamp 1586547711
transform 1 0 3988 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1301
timestamp 1586547711
transform 1 0 5460 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1300
timestamp 1586547711
transform 1 0 5644 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL24380x2720 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 5276 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL23460x0
timestamp 1586547711
transform 1 0 5092 0 -1 944
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL28060x0
timestamp 1586547711
transform 1 0 6012 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_972
timestamp 1586547711
transform 1 0 5828 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_971
timestamp 1586547711
transform 1 0 6748 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1311
timestamp 1586547711
transform 1 0 5828 0 -1 944
box 0 -48 184 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen1
timestamp 1586547711
transform 1 0 6104 0 1 944
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1586547711
transform 1 0 6012 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1586547711
transform 1 0 6104 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL28980x0
timestamp 1586547711
transform 1 0 6196 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1299
timestamp 1586547711
transform 1 0 6932 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1298
timestamp 1586547711
transform 1 0 7760 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL33580x2720
timestamp 1586547711
transform 1 0 7116 0 1 944
box 0 -48 368 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[6\].id.delayint0 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 7484 0 1 944
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL40480x2720
timestamp 1586547711
transform 1 0 8496 0 1 944
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1302
timestamp 1586547711
transform 1 0 7944 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1304
timestamp 1586547711
transform 1 0 8128 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1309
timestamp 1586547711
transform 1 0 8312 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_964
timestamp 1586547711
transform 1 0 8772 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL40020x0
timestamp 1586547711
transform 1 0 8404 0 -1 944
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL34500x0
timestamp 1586547711
transform 1 0 7300 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_59
timestamp 1586547711
transform 1 0 8956 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_76
timestamp 1586547711
transform 1 0 9140 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_581
timestamp 1586547711
transform 1 0 9692 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1292
timestamp 1586547711
transform 1 0 9876 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1586547711
transform 1 0 8956 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[6\].id.delaybuf0 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 9324 0 1 944
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILL51980x2720
timestamp 1586547711
transform 1 0 10796 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1308
timestamp 1586547711
transform 1 0 10060 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_965
timestamp 1586547711
transform 1 0 10888 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL49220x2720
timestamp 1586547711
transform 1 0 10244 0 1 944
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL43240x0
timestamp 1586547711
transform 1 0 9048 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL48760x0
timestamp 1586547711
transform 1 0 10152 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1270
timestamp 1586547711
transform 1 0 11072 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1271
timestamp 1586547711
transform 1 0 11256 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1269
timestamp 1586547711
transform 1 0 11992 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL54280x0
timestamp 1586547711
transform 1 0 11256 0 -1 944
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1586547711
transform 1 0 11624 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1586547711
transform 1 0 11808 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL55200x2720
timestamp 1586547711
transform 1 0 11440 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 11716 0 1 944
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL59800x2720
timestamp 1586547711
transform 1 0 12360 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1280
timestamp 1586547711
transform 1 0 12176 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_60
timestamp 1586547711
transform 1 0 12452 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_75
timestamp 1586547711
transform 1 0 12636 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_592
timestamp 1586547711
transform 1 0 12820 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_967
timestamp 1586547711
transform 1 0 13004 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL57500x0
timestamp 1586547711
transform 1 0 11900 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL63020x0
timestamp 1586547711
transform 1 0 13004 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1286
timestamp 1586547711
transform 1 0 13924 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1285
timestamp 1586547711
transform 1 0 14108 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL68540x0
timestamp 1586547711
transform 1 0 14108 0 -1 944
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL63940x2720
timestamp 1586547711
transform 1 0 13188 0 1 944
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1284
timestamp 1586547711
transform 1 0 14292 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_968
timestamp 1586547711
transform 1 0 15120 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1297
timestamp 1586547711
transform 1 0 14752 0 -1 944
box 0 -48 184 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen1
timestamp 1586547711
transform 1 0 14476 0 1 944
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1586547711
transform 1 0 14660 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL72680x0
timestamp 1586547711
transform 1 0 14936 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_969
timestamp 1586547711
transform 1 0 15304 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1287
timestamp 1586547711
transform 1 0 16132 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL75440x2720
timestamp 1586547711
transform 1 0 15488 0 1 944
box 0 -48 368 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[5\].id.delayint0
timestamp 1586547711
transform 1 0 15856 0 1 944
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1283
timestamp 1586547711
transform 1 0 16316 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1289
timestamp 1586547711
transform 1 0 16500 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1295
timestamp 1586547711
transform 1 0 16684 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL84640x2720
timestamp 1586547711
transform 1 0 17328 0 1 944
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1586547711
transform 1 0 17236 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL82340x2720
timestamp 1586547711
transform 1 0 16868 0 1 944
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILL83720x0
timestamp 1586547711
transform 1 0 17144 0 -1 944
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL78200x0
timestamp 1586547711
transform 1 0 16040 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1586547711
transform 1 0 18340 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1586547711
transform 1 0 17512 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  irb /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 17880 0 1 944
box 0 -48 460 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1170
timestamp 1586547711
transform 1 0 18524 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1586547711
transform 1 0 18708 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_627
timestamp 1586547711
transform 1 0 18892 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_628
timestamp 1586547711
transform 1 0 19444 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp10 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 19076 0 1 944
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL86020x0
timestamp 1586547711
transform 1 0 17604 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL91540x0
timestamp 1586547711
transform 1 0 18708 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL99820x2720
timestamp 1586547711
transform 1 0 20364 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1173
timestamp 1586547711
transform 1 0 19628 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1293
timestamp 1586547711
transform 1 0 19812 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1174
timestamp 1586547711
transform 1 0 20456 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL97060x0
timestamp 1586547711
transform 1 0 19812 0 -1 944
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1586547711
transform 1 0 20364 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL97980x2720
timestamp 1586547711
transform 1 0 19996 0 1 944
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1586547711
transform 1 0 21100 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1586547711
transform 1 0 21284 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_227
timestamp 1586547711
transform 1 0 21468 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _267_
timestamp 1586547711
transform 1 0 20640 0 1 944
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL100280x0
timestamp 1586547711
transform 1 0 20456 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL105800x0
timestamp 1586547711
transform 1 0 21560 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL111780x2720
timestamp 1586547711
transform 1 0 22756 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL112700x2720
timestamp 1586547711
transform 1 0 22940 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_620
timestamp 1586547711
transform 1 0 23032 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1586547711
transform 1 0 22848 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL115920x2720
timestamp 1586547711
transform 1 0 23584 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1586547711
transform 1 0 23216 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1586547711
transform 1 0 23400 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1586547711
transform 1 0 23676 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1586547711
transform 1 0 23216 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL111320x0
timestamp 1586547711
transform 1 0 22664 0 -1 944
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL114540x0
timestamp 1586547711
transform 1 0 23308 0 -1 944
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILL106260x2720
timestamp 1586547711
transform 1 0 21652 0 1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1586547711
transform 1 0 23860 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1018
timestamp 1586547711
transform 1 0 24044 0 -1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1167
timestamp 1586547711
transform 1 0 24228 0 -1 944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL125580x0
timestamp 1586547711
transform 1 0 25516 0 -1 944
box 0 -48 552 592
use sky130_fd_sc_hd__dfrbp_1  idiv2 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 24044 0 1 944
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_12  FILL120060x0
timestamp 1586547711
transform 1 0 24412 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1586547711
transform 1 0 26988 0 1 944
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1586547711
transform 1 0 26988 0 -1 944
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL132480x2720
timestamp 1586547711
transform 1 0 26896 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL132480x0
timestamp 1586547711
transform 1 0 26896 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1586547711
transform 1 0 26160 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_291
timestamp 1586547711
transform 1 0 26344 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1586547711
transform 1 0 26068 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL130640x2720
timestamp 1586547711
transform 1 0 26528 0 1 944
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILL128800x0
timestamp 1586547711
transform 1 0 26160 0 -1 944
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1586547711
transform 1 0 400 0 -1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL4140x5440
timestamp 1586547711
transform 1 0 1228 0 -1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL1380x5440
timestamp 1586547711
transform 1 0 676 0 -1 2032
box 0 -48 552 592
use sky130_fd_sc_hd__a21bo_4  _403_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 1320 0 -1 2032
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_8  FILL10580x5440
timestamp 1586547711
transform 1 0 2516 0 -1 2032
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL14720x5440
timestamp 1586547711
transform 1 0 3344 0 -1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1586547711
transform 1 0 3252 0 -1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__a21bo_4  _397_
timestamp 1586547711
transform 1 0 3620 0 -1 2032
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_3  FILL25760x5440
timestamp 1586547711
transform 1 0 5552 0 -1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[6\].id.delayenb1 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 5828 0 -1 2032
box 0 -48 1012 592
use sky130_fd_sc_hd__decap_8  FILL22080x5440
timestamp 1586547711
transform 1 0 4816 0 -1 2032
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL34500x5440
timestamp 1586547711
transform 1 0 7300 0 -1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL40940x5440
timestamp 1586547711
transform 1 0 8588 0 -1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL32200x5440
timestamp 1586547711
transform 1 0 6840 0 -1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1303
timestamp 1586547711
transform 1 0 6932 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1305
timestamp 1586547711
transform 1 0 7116 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1586547711
transform 1 0 8864 0 -1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp 1586547711
transform 1 0 7576 0 -1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL37260x5440
timestamp 1586547711
transform 1 0 7852 0 -1 2032
box 0 -48 736 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen1
timestamp 1586547711
transform 1 0 10888 0 -1 2032
box 0 -48 644 592
use sky130_fd_sc_hd__a21bo_4  _388_
timestamp 1586547711
transform 1 0 8956 0 -1 2032
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_8  FILL48760x5440
timestamp 1586547711
transform 1 0 10152 0 -1 2032
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1281
timestamp 1586547711
transform 1 0 11716 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL57500x5440
timestamp 1586547711
transform 1 0 11900 0 -1 2032
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILL55660x5440
timestamp 1586547711
transform 1 0 11532 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _393_
timestamp 1586547711
transform 1 0 12452 0 -1 2032
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_1  FILL69920x5440
timestamp 1586547711
transform 1 0 14384 0 -1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1586547711
transform 1 0 14476 0 -1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[5\].id.delayenb1
timestamp 1586547711
transform 1 0 14568 0 -1 2032
box 0 -48 1012 592
use sky130_fd_sc_hd__decap_8  FILL66240x5440
timestamp 1586547711
transform 1 0 13648 0 -1 2032
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1291
timestamp 1586547711
transform 1 0 15580 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL76820x5440
timestamp 1586547711
transform 1 0 15764 0 -1 2032
box 0 -48 552 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp 1586547711
transform 1 0 16316 0 -1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL80960x5440
timestamp 1586547711
transform 1 0 16592 0 -1 2032
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL86480x5440
timestamp 1586547711
transform 1 0 17696 0 -1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1166
timestamp 1586547711
transform 1 0 17788 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1586547711
transform 1 0 17972 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1586547711
transform 1 0 18156 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_629
timestamp 1586547711
transform 1 0 18340 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1021
timestamp 1586547711
transform 1 0 18524 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _417_
timestamp 1586547711
transform 1 0 18708 0 -1 2032
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL94760x5440
timestamp 1586547711
transform 1 0 19352 0 -1 2032
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_625
timestamp 1586547711
transform 1 0 20548 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1586547711
transform 1 0 20088 0 -1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL98900x5440
timestamp 1586547711
transform 1 0 20180 0 -1 2032
box 0 -48 368 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp11 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 20732 0 -1 2032
box 0 -48 1196 592
use sky130_fd_sc_hd__or2_4  _413_
timestamp 1586547711
transform 1 0 23216 0 -1 2032
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILL113160x5440
timestamp 1586547711
transform 1 0 23032 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL107640x5440
timestamp 1586547711
transform 1 0 21928 0 -1 2032
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_225
timestamp 1586547711
transform 1 0 23860 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1586547711
transform 1 0 24044 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_618
timestamp 1586547711
transform 1 0 24228 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1168
timestamp 1586547711
transform 1 0 24412 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1586547711
transform 1 0 25700 0 -1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _284_
timestamp 1586547711
transform 1 0 25792 0 -1 2032
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL120980x5440
timestamp 1586547711
transform 1 0 24596 0 -1 2032
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1586547711
transform 1 0 26988 0 -1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL129260x5440
timestamp 1586547711
transform 1 0 26252 0 -1 2032
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1586547711
transform 1 0 400 0 1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL1380x8160
timestamp 1586547711
transform 1 0 676 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1316
timestamp 1586547711
transform 1 0 768 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1315
timestamp 1586547711
transform 1 0 952 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_978
timestamp 1586547711
transform 1 0 1136 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1325
timestamp 1586547711
transform 1 0 2332 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL10580x8160
timestamp 1586547711
transform 1 0 2516 0 1 2032
box 0 -48 552 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[7\].id.delayenb1
timestamp 1586547711
transform 1 0 1320 0 1 2032
box 0 -48 1012 592
use sky130_fd_sc_hd__fill_1  FILL19320x8160
timestamp 1586547711
transform 1 0 4264 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1312
timestamp 1586547711
transform 1 0 3344 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1323
timestamp 1586547711
transform 1 0 3528 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL16560x8160
timestamp 1586547711
transform 1 0 3712 0 1 2032
box 0 -48 552 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[7\].id.delaybuf0
timestamp 1586547711
transform 1 0 4356 0 1 2032
box 0 -48 368 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp 1586547711
transform 1 0 3068 0 1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1307
timestamp 1586547711
transform 1 0 4724 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1322
timestamp 1586547711
transform 1 0 4908 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1360
timestamp 1586547711
transform 1 0 5092 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL24380x8160
timestamp 1586547711
transform 1 0 5276 0 1 2032
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL28520x8160
timestamp 1586547711
transform 1 0 6104 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1310
timestamp 1586547711
transform 1 0 6196 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1008
timestamp 1586547711
transform 1 0 6380 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1007
timestamp 1586547711
transform 1 0 6564 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1586547711
transform 1 0 6012 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[6\].id.delayenb0 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 6748 0 1 2032
box 0 -48 1656 592
use sky130_fd_sc_hd__decap_12  FILL40020x8160
timestamp 1586547711
transform 1 0 8404 0 1 2032
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1272
timestamp 1586547711
transform 1 0 9508 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_966
timestamp 1586547711
transform 1 0 9692 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL52440x8160
timestamp 1586547711
transform 1 0 10888 0 1 2032
box 0 -48 368 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[4\].id.delayenb1
timestamp 1586547711
transform 1 0 9876 0 1 2032
box 0 -48 1012 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1277
timestamp 1586547711
transform 1 0 11256 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1276
timestamp 1586547711
transform 1 0 11440 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1002
timestamp 1586547711
transform 1 0 11716 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1001
timestamp 1586547711
transform 1 0 12544 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1274
timestamp 1586547711
transform 1 0 12728 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen0
timestamp 1586547711
transform 1 0 11900 0 1 2032
box 0 -48 644 592
use sky130_fd_sc_hd__decap_6  FILL62560x8160
timestamp 1586547711
transform 1 0 12912 0 1 2032
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1586547711
transform 1 0 11624 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL65320x8160
timestamp 1586547711
transform 1 0 13464 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1294
timestamp 1586547711
transform 1 0 13556 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1278
timestamp 1586547711
transform 1 0 14108 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1288
timestamp 1586547711
transform 1 0 14292 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1005
timestamp 1586547711
transform 1 0 14476 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1004
timestamp 1586547711
transform 1 0 14660 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[5\].id.delaybuf0
timestamp 1586547711
transform 1 0 13740 0 1 2032
box 0 -48 368 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[5\].id.delayenb0
timestamp 1586547711
transform 1 0 14844 0 1 2032
box 0 -48 1656 592
use sky130_fd_sc_hd__fill_1  FILL84640x8160
timestamp 1586547711
transform 1 0 17328 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1296
timestamp 1586547711
transform 1 0 16500 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1586547711
transform 1 0 17052 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1586547711
transform 1 0 17236 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL81420x8160
timestamp 1586547711
transform 1 0 16684 0 1 2032
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1586547711
transform 1 0 17420 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1586547711
transform 1 0 17604 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1586547711
transform 1 0 17788 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__dfrbp_1  idiv16
timestamp 1586547711
transform 1 0 17972 0 1 2032
box 0 -48 2116 592
use sky130_fd_sc_hd__fill_1  FILL98440x8160
timestamp 1586547711
transform 1 0 20088 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_619
timestamp 1586547711
transform 1 0 20180 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_228
timestamp 1586547711
transform 1 0 20364 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp 1586547711
transform 1 0 20548 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1586547711
transform 1 0 20732 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _415_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 20916 0 1 2032
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_621
timestamp 1586547711
transform 1 0 22020 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL109940x8160
timestamp 1586547711
transform 1 0 22388 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_623
timestamp 1586547711
transform 1 0 22204 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_224
timestamp 1586547711
transform 1 0 22480 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1586547711
transform 1 0 22664 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1586547711
transform 1 0 22848 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _266_
timestamp 1586547711
transform 1 0 22940 0 1 2032
box 0 -48 460 592
use sky130_fd_sc_hd__fill_1  FILL115000x8160
timestamp 1586547711
transform 1 0 23400 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL116380x8160
timestamp 1586547711
transform 1 0 23676 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1586547711
transform 1 0 23492 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1586547711
transform 1 0 23768 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1586547711
transform 1 0 23952 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__dfrbp_1  idiv4
timestamp 1586547711
transform 1 0 24136 0 1 2032
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1586547711
transform 1 0 26988 0 1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL129260x8160
timestamp 1586547711
transform 1 0 26252 0 1 2032
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1586547711
transform 1 0 400 0 -1 3120
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1320
timestamp 1586547711
transform 1 0 676 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1319
timestamp 1586547711
transform 1 0 860 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1324
timestamp 1586547711
transform 1 0 1044 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1318
timestamp 1586547711
transform 1 0 1688 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL4140x10880
timestamp 1586547711
transform 1 0 1228 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[7\].id.delayint0
timestamp 1586547711
transform 1 0 1412 0 -1 3120
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL7360x10880
timestamp 1586547711
transform 1 0 1872 0 -1 3120
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL12880x10880
timestamp 1586547711
transform 1 0 2976 0 -1 3120
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1586547711
transform 1 0 3252 0 -1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__conb_1  ringosc.iss.const1 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 4448 0 -1 3120
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL14720x10880
timestamp 1586547711
transform 1 0 3344 0 -1 3120
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1306
timestamp 1586547711
transform 1 0 6748 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL30820x10880
timestamp 1586547711
transform 1 0 6564 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL21620x10880
timestamp 1586547711
transform 1 0 4724 0 -1 3120
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL27140x10880
timestamp 1586547711
transform 1 0 5828 0 -1 3120
box 0 -48 736 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen0
timestamp 1586547711
transform 1 0 6932 0 -1 3120
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1586547711
transform 1 0 8864 0 -1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL41400x10880
timestamp 1586547711
transform 1 0 8680 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL35880x10880
timestamp 1586547711
transform 1 0 7576 0 -1 3120
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1183
timestamp 1586547711
transform 1 0 8956 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1282
timestamp 1586547711
transform 1 0 9876 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL48300x10880
timestamp 1586547711
transform 1 0 10060 0 -1 3120
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL43700x10880
timestamp 1586547711
transform 1 0 9140 0 -1 3120
box 0 -48 736 592
use sky130_fd_sc_hd__decap_6  FILL53820x10880
timestamp 1586547711
transform 1 0 11164 0 -1 3120
box 0 -48 552 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[4\].id.delayenb0
timestamp 1586547711
transform 1 0 11716 0 -1 3120
box 0 -48 1656 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen0
timestamp 1586547711
transform 1 0 14936 0 -1 3120
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1586547711
transform 1 0 14476 0 -1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL70840x10880
timestamp 1586547711
transform 1 0 14568 0 -1 3120
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL64860x10880
timestamp 1586547711
transform 1 0 13372 0 -1 3120
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1290
timestamp 1586547711
transform 1 0 15580 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL76820x10880
timestamp 1586547711
transform 1 0 15764 0 -1 3120
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL82340x10880
timestamp 1586547711
transform 1 0 16868 0 -1 3120
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL86020x10880
timestamp 1586547711
transform 1 0 17604 0 -1 3120
box 0 -48 276 592
use sky130_fd_sc_hd__a21bo_4  _418_
timestamp 1586547711
transform 1 0 17880 0 -1 3120
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_8  FILL93380x10880
timestamp 1586547711
transform 1 0 19076 0 -1 3120
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL97060x10880
timestamp 1586547711
transform 1 0 19812 0 -1 3120
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_626
timestamp 1586547711
transform 1 0 20364 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_624
timestamp 1586547711
transform 1 0 20548 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1586547711
transform 1 0 20088 0 -1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL98900x10880
timestamp 1586547711
transform 1 0 20180 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__a32oi_4  _416_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 20732 0 -1 3120
box 0 -48 2024 592
use sky130_fd_sc_hd__or2_4  _412_
timestamp 1586547711
transform 1 0 23492 0 -1 3120
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL111780x10880
timestamp 1586547711
transform 1 0 22756 0 -1 3120
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL126040x10880
timestamp 1586547711
transform 1 0 25608 0 -1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1586547711
transform 1 0 24136 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1019
timestamp 1586547711
transform 1 0 24320 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1586547711
transform 1 0 25700 0 -1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL120520x10880
timestamp 1586547711
transform 1 0 24504 0 -1 3120
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL126960x10880
timestamp 1586547711
transform 1 0 25792 0 -1 3120
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1586547711
transform 1 0 26988 0 -1 3120
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL132480x10880
timestamp 1586547711
transform 1 0 26896 0 -1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1586547711
transform 1 0 400 0 1 3120
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1011
timestamp 1586547711
transform 1 0 676 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1010
timestamp 1586547711
transform 1 0 1504 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1317
timestamp 1586547711
transform 1 0 1688 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen0
timestamp 1586547711
transform 1 0 860 0 1 3120
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL7360x13600
timestamp 1586547711
transform 1 0 1872 0 1 3120
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL17480x13600
timestamp 1586547711
transform 1 0 3896 0 1 3120
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_938
timestamp 1586547711
transform 1 0 3344 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_950
timestamp 1586547711
transform 1 0 3528 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1351
timestamp 1586547711
transform 1 0 3712 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_939
timestamp 1586547711
transform 1 0 4632 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL12880x13600
timestamp 1586547711
transform 1 0 2976 0 1 3120
box 0 -48 368 592
use sky130_fd_sc_hd__einvp_1  ringosc.iss.reseten0 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 4172 0 1 3120
box 0 -48 460 592
use sky130_fd_sc_hd__fill_1  FILL25760x13600
timestamp 1586547711
transform 1 0 5552 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1186
timestamp 1586547711
transform 1 0 4816 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1361
timestamp 1586547711
transform 1 0 5000 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_937
timestamp 1586547711
transform 1 0 5644 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_134
timestamp 1586547711
transform 1 0 5828 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1586547711
transform 1 0 6012 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL23920x13600
timestamp 1586547711
transform 1 0 5184 0 1 3120
box 0 -48 368 592
use sky130_fd_sc_hd__nor2_4  _288_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 6104 0 1 3120
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  FILL37260x13600
timestamp 1586547711
transform 1 0 7852 0 1 3120
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp 1586547711
transform 1 0 6932 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1172
timestamp 1586547711
transform 1 0 8128 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1047
timestamp 1586547711
transform 1 0 8312 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp01
timestamp 1586547711
transform 1 0 8496 0 1 3120
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_8  FILL33580x13600
timestamp 1586547711
transform 1 0 7116 0 1 3120
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1171
timestamp 1586547711
transform 1 0 9692 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL52900x13600
timestamp 1586547711
transform 1 0 10980 0 1 3120
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL47380x13600
timestamp 1586547711
transform 1 0 9876 0 1 3120
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL55660x13600
timestamp 1586547711
transform 1 0 11532 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1273
timestamp 1586547711
transform 1 0 11992 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1275
timestamp 1586547711
transform 1 0 12176 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1586547711
transform 1 0 11624 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[4\].id.delayint0
timestamp 1586547711
transform 1 0 11716 0 1 3120
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL59800x13600
timestamp 1586547711
transform 1 0 12360 0 1 3120
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL73600x13600
timestamp 1586547711
transform 1 0 15120 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_127
timestamp 1586547711
transform 1 0 15212 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL70840x13600
timestamp 1586547711
transform 1 0 14568 0 1 3120
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL65320x13600
timestamp 1586547711
transform 1 0 13464 0 1 3120
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_909
timestamp 1586547711
transform 1 0 15396 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1032
timestamp 1586547711
transform 1 0 15580 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1129
timestamp 1586547711
transform 1 0 15764 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1586547711
transform 1 0 17236 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL83260x13600
timestamp 1586547711
transform 1 0 17052 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _532_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 17328 0 1 3120
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL77740x13600
timestamp 1586547711
transform 1 0 15948 0 1 3120
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_143
timestamp 1586547711
transform 1 0 17880 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_908
timestamp 1586547711
transform 1 0 18064 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL89240x13600
timestamp 1586547711
transform 1 0 18248 0 1 3120
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL94760x13600
timestamp 1586547711
transform 1 0 19352 0 1 3120
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL102120x13600
timestamp 1586547711
transform 1 0 20824 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1022
timestamp 1586547711
transform 1 0 20916 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL100280x13600
timestamp 1586547711
transform 1 0 20456 0 1 3120
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL103500x13600
timestamp 1586547711
transform 1 0 21100 0 1 3120
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_622
timestamp 1586547711
transform 1 0 22388 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1586547711
transform 1 0 22572 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL109020x13600
timestamp 1586547711
transform 1 0 22204 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL111780x13600
timestamp 1586547711
transform 1 0 22756 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL113620x13600
timestamp 1586547711
transform 1 0 23124 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_226
timestamp 1586547711
transform 1 0 22940 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1586547711
transform 1 0 23216 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1586547711
transform 1 0 23400 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1586547711
transform 1 0 22848 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__dfrbp_1  idiv8
timestamp 1586547711
transform 1 0 23584 0 1 3120
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_12  FILL126500x13600
timestamp 1586547711
transform 1 0 25700 0 1 3120
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1586547711
transform 1 0 26988 0 1 3120
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILL132020x13600
timestamp 1586547711
transform 1 0 26804 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1586547711
transform 1 0 400 0 1 4208
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL6900x19040
timestamp 1586547711
transform 1 0 1780 0 1 4208
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1586547711
transform 1 0 400 0 -1 4208
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1221
timestamp 1586547711
transform 1 0 2056 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1185
timestamp 1586547711
transform 1 0 2240 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__einvn_8  ringosc.iss.delayenb0
timestamp 1586547711
transform 1 0 2424 0 1 4208
box 0 -48 1656 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[7\].id.delayenb0
timestamp 1586547711
transform 1 0 676 0 -1 4208
box 0 -48 1656 592
use sky130_fd_sc_hd__decap_12  FILL1380x19040
timestamp 1586547711
transform 1 0 676 0 1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL9660x16320
timestamp 1586547711
transform 1 0 2332 0 -1 4208
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL18400x19040
timestamp 1586547711
transform 1 0 4080 0 1 4208
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_948
timestamp 1586547711
transform 1 0 4356 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1219
timestamp 1586547711
transform 1 0 4540 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1586547711
transform 1 0 3252 0 -1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL13340x16320
timestamp 1586547711
transform 1 0 3068 0 -1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__or2_2  ringosc.iss.ctrlen0 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 3344 0 -1 4208
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL17020x16320
timestamp 1586547711
transform 1 0 3804 0 -1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL31280x19040
timestamp 1586547711
transform 1 0 6656 0 1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1225
timestamp 1586547711
transform 1 0 4724 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1215
timestamp 1586547711
transform 1 0 6748 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL28520x19040
timestamp 1586547711
transform 1 0 6104 0 1 4208
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1586547711
transform 1 0 6012 0 1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL22540x19040
timestamp 1586547711
transform 1 0 4908 0 1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL22540x16320
timestamp 1586547711
transform 1 0 4908 0 -1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL28060x16320
timestamp 1586547711
transform 1 0 6012 0 -1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL41860x16320
timestamp 1586547711
transform 1 0 8772 0 -1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1217
timestamp 1586547711
transform 1 0 6932 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL39100x16320
timestamp 1586547711
transform 1 0 8220 0 -1 4208
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1586547711
transform 1 0 8864 0 -1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL33580x19040
timestamp 1586547711
transform 1 0 7116 0 1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL33580x16320
timestamp 1586547711
transform 1 0 7116 0 -1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL39100x19040
timestamp 1586547711
transform 1 0 8220 0 1 4208
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL42780x19040
timestamp 1586547711
transform 1 0 8956 0 1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_146
timestamp 1586547711
transform 1 0 9048 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_914
timestamp 1586547711
transform 1 0 9232 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_129
timestamp 1586547711
transform 1 0 10888 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL50600x19040
timestamp 1586547711
transform 1 0 10520 0 1 4208
box 0 -48 368 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp00
timestamp 1586547711
transform 1 0 8956 0 -1 4208
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL45080x19040
timestamp 1586547711
transform 1 0 9416 0 1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL44620x16320
timestamp 1586547711
transform 1 0 9324 0 -1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL50140x16320
timestamp 1586547711
transform 1 0 10428 0 -1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL56580x19040
timestamp 1586547711
transform 1 0 11716 0 1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_911
timestamp 1586547711
transform 1 0 11072 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1033
timestamp 1586547711
transform 1 0 11256 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1135
timestamp 1586547711
transform 1 0 11440 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1586547711
transform 1 0 11624 0 1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _533_
timestamp 1586547711
transform 1 0 11808 0 1 4208
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_144
timestamp 1586547711
transform 1 0 12360 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_910
timestamp 1586547711
transform 1 0 12544 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL61640x19040
timestamp 1586547711
transform 1 0 12728 0 1 4208
box 0 -48 368 592
use sky130_fd_sc_hd__inv_4  _512_
timestamp 1586547711
transform 1 0 13096 0 1 4208
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL55660x16320
timestamp 1586547711
transform 1 0 11532 0 -1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL61180x16320
timestamp 1586547711
transform 1 0 12636 0 -1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_870
timestamp 1586547711
transform 1 0 13556 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_872
timestamp 1586547711
transform 1 0 13740 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL67620x19040
timestamp 1586547711
transform 1 0 13924 0 1 4208
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL66700x16320
timestamp 1586547711
transform 1 0 13740 0 -1 4208
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL70380x19040
timestamp 1586547711
transform 1 0 14476 0 1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL73600x16320
timestamp 1586547711
transform 1 0 15120 0 -1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_866
timestamp 1586547711
transform 1 0 14568 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_867
timestamp 1586547711
transform 1 0 14752 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL70840x16320
timestamp 1586547711
transform 1 0 14568 0 -1 4208
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1586547711
transform 1 0 14476 0 -1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL72680x19040
timestamp 1586547711
transform 1 0 14936 0 1 4208
box 0 -48 736 592
use sky130_fd_sc_hd__dfrtp_4  _555_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 15212 0 -1 4208
box 0 -48 2116 592
use sky130_fd_sc_hd__fill_1  FILL76360x19040
timestamp 1586547711
transform 1 0 15672 0 1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_825
timestamp 1586547711
transform 1 0 15764 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_854
timestamp 1586547711
transform 1 0 15948 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_862
timestamp 1586547711
transform 1 0 16132 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1586547711
transform 1 0 17236 0 1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL83260x19040
timestamp 1586547711
transform 1 0 17052 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL84640x19040
timestamp 1586547711
transform 1 0 17328 0 1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL84640x16320
timestamp 1586547711
transform 1 0 17328 0 -1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL79580x19040
timestamp 1586547711
transform 1 0 16316 0 1 4208
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL90160x19040
timestamp 1586547711
transform 1 0 18432 0 1 4208
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL93380x19040
timestamp 1586547711
transform 1 0 19076 0 1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_297
timestamp 1586547711
transform 1 0 18708 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1161
timestamp 1586547711
transform 1 0 18892 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _530_
timestamp 1586547711
transform 1 0 19168 0 1 4208
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL90160x16320
timestamp 1586547711
transform 1 0 18432 0 -1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_141
timestamp 1586547711
transform 1 0 19720 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_904
timestamp 1586547711
transform 1 0 19904 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL95680x16320
timestamp 1586547711
transform 1 0 19536 0 -1 4208
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1586547711
transform 1 0 20088 0 -1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL98440x19040
timestamp 1586547711
transform 1 0 20088 0 1 4208
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_121
timestamp 1586547711
transform 1 0 21008 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_903
timestamp 1586547711
transform 1 0 21192 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1029
timestamp 1586547711
transform 1 0 21376 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1160
timestamp 1586547711
transform 1 0 21560 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL102120x19040
timestamp 1586547711
transform 1 0 20824 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL98900x16320
timestamp 1586547711
transform 1 0 20180 0 -1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL104420x16320
timestamp 1586547711
transform 1 0 21284 0 -1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1586547711
transform 1 0 23584 0 -1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1586547711
transform 1 0 22848 0 1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL114080x16320
timestamp 1586547711
transform 1 0 23216 0 -1 4208
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _414_
timestamp 1586547711
transform 1 0 22572 0 -1 4208
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILL109940x16320
timestamp 1586547711
transform 1 0 22388 0 -1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL106720x19040
timestamp 1586547711
transform 1 0 21744 0 1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL112700x19040
timestamp 1586547711
transform 1 0 22940 0 1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_152
timestamp 1586547711
transform 1 0 24412 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_926
timestamp 1586547711
transform 1 0 24596 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1020
timestamp 1586547711
transform 1 0 23768 0 -1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1169
timestamp 1586547711
transform 1 0 23952 0 -1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL118220x19040
timestamp 1586547711
transform 1 0 24044 0 1 4208
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILL126040x16320
timestamp 1586547711
transform 1 0 25608 0 -1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1586547711
transform 1 0 25700 0 -1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL124200x16320
timestamp 1586547711
transform 1 0 25240 0 -1 4208
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL121900x19040
timestamp 1586547711
transform 1 0 24780 0 1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL118680x16320
timestamp 1586547711
transform 1 0 24136 0 -1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL126960x16320
timestamp 1586547711
transform 1 0 25792 0 -1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1586547711
transform 1 0 26988 0 1 4208
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1586547711
transform 1 0 26988 0 -1 4208
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL132480x16320
timestamp 1586547711
transform 1 0 26896 0 -1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL127420x19040
timestamp 1586547711
transform 1 0 25884 0 1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1586547711
transform 1 0 400 0 -1 5296
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL9660x21760
timestamp 1586547711
transform 1 0 2332 0 -1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1352
timestamp 1586547711
transform 1 0 2424 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL6900x21760
timestamp 1586547711
transform 1 0 1780 0 -1 5296
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL1380x21760
timestamp 1586547711
transform 1 0 676 0 -1 5296
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL13800x21760
timestamp 1586547711
transform 1 0 3160 0 -1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL19320x21760
timestamp 1586547711
transform 1 0 4264 0 -1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1353
timestamp 1586547711
transform 1 0 3344 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_946
timestamp 1586547711
transform 1 0 4080 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL11040x21760
timestamp 1586547711
transform 1 0 2608 0 -1 5296
box 0 -48 552 592
use sky130_fd_sc_hd__decap_6  FILL15640x21760
timestamp 1586547711
transform 1 0 3528 0 -1 5296
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1586547711
transform 1 0 3252 0 -1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[11\].id.delayenb0
timestamp 1586547711
transform 1 0 4356 0 -1 5296
box 0 -48 1656 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1214
timestamp 1586547711
transform 1 0 6380 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL28060x21760
timestamp 1586547711
transform 1 0 6012 0 -1 5296
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL30820x21760
timestamp 1586547711
transform 1 0 6564 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[11\].id.delayint0
timestamp 1586547711
transform 1 0 6748 0 -1 5296
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1158
timestamp 1586547711
transform 1 0 8680 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL38640x21760
timestamp 1586547711
transform 1 0 8128 0 -1 5296
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1586547711
transform 1 0 8864 0 -1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL33120x21760
timestamp 1586547711
transform 1 0 7024 0 -1 5296
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL42780x21760
timestamp 1586547711
transform 1 0 8956 0 -1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_132
timestamp 1586547711
transform 1 0 9600 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_889
timestamp 1586547711
transform 1 0 9784 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_891
timestamp 1586547711
transform 1 0 9968 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1157
timestamp 1586547711
transform 1 0 10152 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL49680x21760
timestamp 1586547711
transform 1 0 10336 0 -1 5296
box 0 -48 552 592
use sky130_fd_sc_hd__buf_4  _535_
timestamp 1586547711
transform 1 0 9048 0 -1 5296
box 0 -48 552 592
use sky130_fd_sc_hd__dfrtp_4  _556_
timestamp 1586547711
transform 1 0 10888 0 -1 5296
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_12  FILL63020x21760
timestamp 1586547711
transform 1 0 13004 0 -1 5296
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_864
timestamp 1586547711
transform 1 0 15028 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_869
timestamp 1586547711
transform 1 0 15212 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1586547711
transform 1 0 14476 0 -1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL68540x21760
timestamp 1586547711
transform 1 0 14108 0 -1 5296
box 0 -48 368 592
use sky130_fd_sc_hd__inv_4  _509_
timestamp 1586547711
transform 1 0 14568 0 -1 5296
box 0 -48 460 592
use sky130_fd_sc_hd__decap_4  FILL74980x21760
timestamp 1586547711
transform 1 0 15396 0 -1 5296
box 0 -48 368 592
use sky130_fd_sc_hd__and2_4  _507_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 15764 0 -1 5296
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL80040x21760
timestamp 1586547711
transform 1 0 16408 0 -1 5296
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL85560x21760
timestamp 1586547711
transform 1 0 17512 0 -1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1112
timestamp 1586547711
transform 1 0 17604 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1164
timestamp 1586547711
transform 1 0 17788 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_905
timestamp 1586547711
transform 1 0 17972 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1030
timestamp 1586547711
transform 1 0 18156 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1165
timestamp 1586547711
transform 1 0 18340 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL90620x21760
timestamp 1586547711
transform 1 0 18524 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _286_
timestamp 1586547711
transform 1 0 18708 0 -1 5296
box 0 -48 460 592
use sky130_fd_sc_hd__decap_8  FILL93840x21760
timestamp 1586547711
transform 1 0 19168 0 -1 5296
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL102580x21760
timestamp 1586547711
transform 1 0 20916 0 -1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1586547711
transform 1 0 20088 0 -1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL97520x21760
timestamp 1586547711
transform 1 0 19904 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _552_
timestamp 1586547711
transform 1 0 21008 0 -1 5296
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_8  FILL98900x21760
timestamp 1586547711
transform 1 0 20180 0 -1 5296
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL113620x21760
timestamp 1586547711
transform 1 0 23124 0 -1 5296
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1041
timestamp 1586547711
transform 1 0 23860 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_94
timestamp 1586547711
transform 1 0 24228 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1586547711
transform 1 0 25700 0 -1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL118220x21760
timestamp 1586547711
transform 1 0 24044 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _541_
timestamp 1586547711
transform 1 0 24412 0 -1 5296
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL126960x21760
timestamp 1586547711
transform 1 0 25792 0 -1 5296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL122820x21760
timestamp 1586547711
transform 1 0 24964 0 -1 5296
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1586547711
transform 1 0 26988 0 -1 5296
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL132480x21760
timestamp 1586547711
transform 1 0 26896 0 -1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1586547711
transform 1 0 400 0 1 5296
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL8740x24480
timestamp 1586547711
transform 1 0 2148 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_49
timestamp 1586547711
transform 1 0 676 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_86
timestamp 1586547711
transform 1 0 860 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_478
timestamp 1586547711
transform 1 0 1044 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1009
timestamp 1586547711
transform 1 0 1228 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1358
timestamp 1586547711
transform 1 0 2240 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen0
timestamp 1586547711
transform 1 0 2424 0 1 5296
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL5060x24480
timestamp 1586547711
transform 1 0 1412 0 1 5296
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL16100x24480
timestamp 1586547711
transform 1 0 3620 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_951
timestamp 1586547711
transform 1 0 3068 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1184
timestamp 1586547711
transform 1 0 3252 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1220
timestamp 1586547711
transform 1 0 3436 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_82
timestamp 1586547711
transform 1 0 3712 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_53
timestamp 1586547711
transform 1 0 3896 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _349_
timestamp 1586547711
transform 1 0 4080 0 1 5296
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA_947
timestamp 1586547711
transform 1 0 5276 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1216
timestamp 1586547711
transform 1 0 5460 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1218
timestamp 1586547711
transform 1 0 5644 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1226
timestamp 1586547711
transform 1 0 5828 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL28520x24480
timestamp 1586547711
transform 1 0 6104 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL30820x24480
timestamp 1586547711
transform 1 0 6564 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1213
timestamp 1586547711
transform 1 0 6196 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_990
timestamp 1586547711
transform 1 0 6380 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1586547711
transform 1 0 6012 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen1
timestamp 1586547711
transform 1 0 6656 0 1 5296
box 0 -48 644 592
use sky130_fd_sc_hd__fill_1  FILL39100x24480
timestamp 1586547711
transform 1 0 8220 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_989
timestamp 1586547711
transform 1 0 7300 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1212
timestamp 1586547711
transform 1 0 7484 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_915
timestamp 1586547711
transform 1 0 8312 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_133
timestamp 1586547711
transform 1 0 8496 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL36340x24480
timestamp 1586547711
transform 1 0 7668 0 1 5296
box 0 -48 552 592
use sky130_fd_sc_hd__dfrtp_4  _558_
timestamp 1586547711
transform 1 0 8680 0 1 5296
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_3  FILL51980x24480
timestamp 1586547711
transform 1 0 10796 0 1 5296
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_873
timestamp 1586547711
transform 1 0 11072 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_168
timestamp 1586547711
transform 1 0 11256 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_128
timestamp 1586547711
transform 1 0 11440 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL63020x24480
timestamp 1586547711
transform 1 0 13004 0 1 5296
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1586547711
transform 1 0 11624 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _513_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 11716 0 1 5296
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA_868
timestamp 1586547711
transform 1 0 13556 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_861
timestamp 1586547711
transform 1 0 13740 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_850
timestamp 1586547711
transform 1 0 13924 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_849
timestamp 1586547711
transform 1 0 14108 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_126
timestamp 1586547711
transform 1 0 14292 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _510_
timestamp 1586547711
transform 1 0 14476 0 1 5296
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_1  FILL84640x24480
timestamp 1586547711
transform 1 0 17328 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1127
timestamp 1586547711
transform 1 0 15764 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_824
timestamp 1586547711
transform 1 0 15948 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_859
timestamp 1586547711
transform 1 0 16132 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_860
timestamp 1586547711
transform 1 0 16316 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1126
timestamp 1586547711
transform 1 0 17052 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL80500x24480
timestamp 1586547711
transform 1 0 16500 0 1 5296
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1586547711
transform 1 0 17236 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_852
timestamp 1586547711
transform 1 0 17420 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_796
timestamp 1586547711
transform 1 0 17604 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_123
timestamp 1586547711
transform 1 0 17788 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _553_
timestamp 1586547711
transform 1 0 17972 0 1 5296
box 0 -48 2116 592
use sky130_fd_sc_hd__fill_1  FILL98440x24480
timestamp 1586547711
transform 1 0 20088 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL104420x24480
timestamp 1586547711
transform 1 0 21284 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_795
timestamp 1586547711
transform 1 0 20180 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_797
timestamp 1586547711
transform 1 0 20364 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1162
timestamp 1586547711
transform 1 0 20548 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_902
timestamp 1586547711
transform 1 0 21376 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL101660x24480
timestamp 1586547711
transform 1 0 20732 0 1 5296
box 0 -48 552 592
use sky130_fd_sc_hd__buf_4  _529_
timestamp 1586547711
transform 1 0 21560 0 1 5296
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_140
timestamp 1586547711
transform 1 0 22112 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_282
timestamp 1586547711
transform 1 0 22296 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1159
timestamp 1586547711
transform 1 0 22480 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1096
timestamp 1586547711
transform 1 0 23308 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_632
timestamp 1586547711
transform 1 0 23492 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_95
timestamp 1586547711
transform 1 0 23676 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1586547711
transform 1 0 22848 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL112700x24480
timestamp 1586547711
transform 1 0 22940 0 1 5296
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL111320x24480
timestamp 1586547711
transform 1 0 22664 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _564_
timestamp 1586547711
transform 1 0 23860 0 1 5296
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_3  FILL131560x24480
timestamp 1586547711
transform 1 0 26712 0 1 5296
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1586547711
transform 1 0 26988 0 1 5296
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL127880x24480
timestamp 1586547711
transform 1 0 25976 0 1 5296
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1586547711
transform 1 0 400 0 -1 6384
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1355
timestamp 1586547711
transform 1 0 1872 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _344_
timestamp 1586547711
transform 1 0 676 0 -1 6384
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_12  FILL8280x27200
timestamp 1586547711
transform 1 0 2056 0 -1 6384
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL13800x27200
timestamp 1586547711
transform 1 0 3160 0 -1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL17940x27200
timestamp 1586547711
transform 1 0 3988 0 -1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_461
timestamp 1586547711
transform 1 0 4080 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL19320x27200
timestamp 1586547711
transform 1 0 4264 0 -1 6384
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1586547711
transform 1 0 3252 0 -1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL16100x27200
timestamp 1586547711
transform 1 0 3620 0 -1 6384
box 0 -48 368 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.iss.delaybuf0
timestamp 1586547711
transform 1 0 3344 0 -1 6384
box 0 -48 276 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen0
timestamp 1586547711
transform 1 0 4816 0 -1 6384
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILL28980x27200
timestamp 1586547711
transform 1 0 6196 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[11\].id.delayenb1
timestamp 1586547711
transform 1 0 6380 0 -1 6384
box 0 -48 1012 592
use sky130_fd_sc_hd__decap_8  FILL25300x27200
timestamp 1586547711
transform 1 0 5460 0 -1 6384
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1035
timestamp 1586547711
transform 1 0 8680 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1586547711
transform 1 0 8864 0 -1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL40480x27200
timestamp 1586547711
transform 1 0 8496 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL34960x27200
timestamp 1586547711
transform 1 0 7392 0 -1 6384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILL42780x27200
timestamp 1586547711
transform 1 0 8956 0 -1 6384
box 0 -48 368 592
use sky130_fd_sc_hd__a21bo_4  _523_
timestamp 1586547711
transform 1 0 9324 0 -1 6384
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_12  FILL50600x27200
timestamp 1586547711
transform 1 0 10520 0 -1 6384
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL56120x27200
timestamp 1586547711
transform 1 0 11624 0 -1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_871
timestamp 1586547711
transform 1 0 11716 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1134
timestamp 1586547711
transform 1 0 11900 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL58420x27200
timestamp 1586547711
transform 1 0 12084 0 -1 6384
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_856
timestamp 1586547711
transform 1 0 15212 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1586547711
transform 1 0 14476 0 -1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _511_
timestamp 1586547711
transform 1 0 14568 0 -1 6384
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILL69460x27200
timestamp 1586547711
transform 1 0 14292 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL63940x27200
timestamp 1586547711
transform 1 0 13188 0 -1 6384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL84640x27200
timestamp 1586547711
transform 1 0 17328 0 -1 6384
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_865
timestamp 1586547711
transform 1 0 15396 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL75900x27200
timestamp 1586547711
transform 1 0 15580 0 -1 6384
box 0 -48 368 592
use sky130_fd_sc_hd__and2_4  _506_
timestamp 1586547711
transform 1 0 15948 0 -1 6384
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL80960x27200
timestamp 1586547711
transform 1 0 16592 0 -1 6384
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_792
timestamp 1586547711
transform 1 0 18432 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_805
timestamp 1586547711
transform 1 0 18616 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _503_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 17604 0 -1 6384
box 0 -48 828 592
use sky130_fd_sc_hd__decap_12  FILL92000x27200
timestamp 1586547711
transform 1 0 18800 0 -1 6384
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_789
timestamp 1586547711
transform 1 0 20824 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1586547711
transform 1 0 20088 0 -1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _484_
timestamp 1586547711
transform 1 0 20180 0 -1 6384
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILL97520x27200
timestamp 1586547711
transform 1 0 19904 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL103040x27200
timestamp 1586547711
transform 1 0 21008 0 -1 6384
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL106720x27200
timestamp 1586547711
transform 1 0 21744 0 -1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL115000x27200
timestamp 1586547711
transform 1 0 23400 0 -1 6384
box 0 -48 368 592
use sky130_fd_sc_hd__inv_4  _281_
timestamp 1586547711
transform 1 0 21836 0 -1 6384
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL109480x27200
timestamp 1586547711
transform 1 0 22296 0 -1 6384
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL116840x27200
timestamp 1586547711
transform 1 0 23768 0 -1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL126040x27200
timestamp 1586547711
transform 1 0 25608 0 -1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_927
timestamp 1586547711
transform 1 0 23860 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1097
timestamp 1586547711
transform 1 0 24044 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1586547711
transform 1 0 25700 0 -1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _421_
timestamp 1586547711
transform 1 0 24228 0 -1 6384
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL126960x27200
timestamp 1586547711
transform 1 0 25792 0 -1 6384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL122360x27200
timestamp 1586547711
transform 1 0 24872 0 -1 6384
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1586547711
transform 1 0 26988 0 -1 6384
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL132480x27200
timestamp 1586547711
transform 1 0 26896 0 -1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1586547711
transform 1 0 400 0 1 6384
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1354
timestamp 1586547711
transform 1 0 860 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1222
timestamp 1586547711
transform 1 0 1044 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_993
timestamp 1586547711
transform 1 0 1228 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_992
timestamp 1586547711
transform 1 0 2424 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL1380x29920
timestamp 1586547711
transform 1 0 676 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__einvn_4  ringosc.iss.delayenb1
timestamp 1586547711
transform 1 0 1412 0 1 6384
box 0 -48 1012 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1357
timestamp 1586547711
transform 1 0 3436 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1359
timestamp 1586547711
transform 1 0 3620 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL11040x29920
timestamp 1586547711
transform 1 0 2608 0 1 6384
box 0 -48 552 592
use sky130_fd_sc_hd__clkinv_1  ringosc.iss.delayint0
timestamp 1586547711
transform 1 0 3160 0 1 6384
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL17020x29920
timestamp 1586547711
transform 1 0 3804 0 1 6384
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_512
timestamp 1586547711
transform 1 0 5828 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_589
timestamp 1586547711
transform 1 0 6104 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_591
timestamp 1586547711
transform 1 0 6288 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1124
timestamp 1586547711
transform 1 0 6472 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1586547711
transform 1 0 6012 0 1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL26220x29920
timestamp 1586547711
transform 1 0 5644 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL31280x29920
timestamp 1586547711
transform 1 0 6656 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL22540x29920
timestamp 1586547711
transform 1 0 4908 0 1 6384
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1211
timestamp 1586547711
transform 1 0 7116 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1224
timestamp 1586547711
transform 1 0 7300 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1155
timestamp 1586547711
transform 1 0 8588 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1140
timestamp 1586547711
transform 1 0 8772 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp 1586547711
transform 1 0 6840 0 1 6384
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL35420x29920
timestamp 1586547711
transform 1 0 7484 0 1 6384
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_66
timestamp 1586547711
transform 1 0 8956 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_69
timestamp 1586547711
transform 1 0 9140 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_189
timestamp 1586547711
transform 1 0 9324 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_988
timestamp 1586547711
transform 1 0 9508 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_888
timestamp 1586547711
transform 1 0 10336 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_890
timestamp 1586547711
transform 1 0 10520 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1156
timestamp 1586547711
transform 1 0 10704 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL52440x29920
timestamp 1586547711
transform 1 0 10888 0 1 6384
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _522_
timestamp 1586547711
transform 1 0 9692 0 1 6384
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  FILL60260x29920
timestamp 1586547711
transform 1 0 12452 0 1 6384
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_163
timestamp 1586547711
transform 1 0 11256 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1130
timestamp 1586547711
transform 1 0 11440 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_169
timestamp 1586547711
transform 1 0 12728 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_857
timestamp 1586547711
transform 1 0 12912 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_874
timestamp 1586547711
transform 1 0 13096 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1586547711
transform 1 0 11624 0 1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL56580x29920
timestamp 1586547711
transform 1 0 11716 0 1 6384
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL68080x29920
timestamp 1586547711
transform 1 0 14016 0 1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_863
timestamp 1586547711
transform 1 0 14108 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_858
timestamp 1586547711
transform 1 0 14292 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_843
timestamp 1586547711
transform 1 0 14476 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_819
timestamp 1586547711
transform 1 0 14660 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_781
timestamp 1586547711
transform 1 0 14844 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__or3_4  _505_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 15028 0 1 6384
box 0 -48 828 592
use sky130_fd_sc_hd__decap_8  FILL64400x29920
timestamp 1586547711
transform 1 0 13280 0 1 6384
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL82800x29920
timestamp 1586547711
transform 1 0 16960 0 1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL84640x29920
timestamp 1586547711
transform 1 0 17328 0 1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_801
timestamp 1586547711
transform 1 0 15856 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1113
timestamp 1586547711
transform 1 0 16040 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_841
timestamp 1586547711
transform 1 0 17052 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1586547711
transform 1 0 17236 0 1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL79120x29920
timestamp 1586547711
transform 1 0 16224 0 1 6384
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_799
timestamp 1586547711
transform 1 0 17420 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_299
timestamp 1586547711
transform 1 0 17604 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_285
timestamp 1586547711
transform 1 0 17788 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_221
timestamp 1586547711
transform 1 0 18800 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_298
timestamp 1586547711
transform 1 0 18984 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL93840x29920
timestamp 1586547711
transform 1 0 19168 0 1 6384
box 0 -48 368 592
use sky130_fd_sc_hd__or3_4  _500_
timestamp 1586547711
transform 1 0 17972 0 1 6384
box 0 -48 828 592
use sky130_fd_sc_hd__fill_1  FILL95680x29920
timestamp 1586547711
transform 1 0 19536 0 1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_790
timestamp 1586547711
transform 1 0 19628 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_774
timestamp 1586547711
transform 1 0 19812 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_284
timestamp 1586547711
transform 1 0 19996 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_283
timestamp 1586547711
transform 1 0 20180 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_120
timestamp 1586547711
transform 1 0 20364 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__o22ai_4  _483_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 20548 0 1 6384
box 0 -48 1472 592
use sky130_fd_sc_hd__decap_3  FILL116380x29920
timestamp 1586547711
transform 1 0 23676 0 1 6384
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL111780x29920
timestamp 1586547711
transform 1 0 22756 0 1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_791
timestamp 1586547711
transform 1 0 22020 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_793
timestamp 1586547711
transform 1 0 22204 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1586547711
transform 1 0 22848 0 1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL109940x29920
timestamp 1586547711
transform 1 0 22388 0 1 6384
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILL112700x29920
timestamp 1586547711
transform 1 0 22940 0 1 6384
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_229
timestamp 1586547711
transform 1 0 24412 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1095
timestamp 1586547711
transform 1 0 24596 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_153
timestamp 1586547711
transform 1 0 25700 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL121900x29920
timestamp 1586547711
transform 1 0 24780 0 1 6384
box 0 -48 368 592
use sky130_fd_sc_hd__inv_4  _268_
timestamp 1586547711
transform 1 0 23952 0 1 6384
box 0 -48 460 592
use sky130_fd_sc_hd__buf_4  _542_
timestamp 1586547711
transform 1 0 25148 0 1 6384
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1586547711
transform 1 0 26988 0 1 6384
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_928
timestamp 1586547711
transform 1 0 25884 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL132020x29920
timestamp 1586547711
transform 1 0 26804 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL128340x29920
timestamp 1586547711
transform 1 0 26068 0 1 6384
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1586547711
transform 1 0 400 0 -1 7472
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1356
timestamp 1586547711
transform 1 0 1412 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen1
timestamp 1586547711
transform 1 0 1596 0 -1 7472
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL1380x32640
timestamp 1586547711
transform 1 0 676 0 -1 7472
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL9200x32640
timestamp 1586547711
transform 1 0 2240 0 -1 7472
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL12880x32640
timestamp 1586547711
transform 1 0 2976 0 -1 7472
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1586547711
transform 1 0 3252 0 -1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL14720x32640
timestamp 1586547711
transform 1 0 3344 0 -1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL20240x32640
timestamp 1586547711
transform 1 0 4448 0 -1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL25760x32640
timestamp 1586547711
transform 1 0 5552 0 -1 7472
box 0 -48 276 592
use sky130_fd_sc_hd__a21o_4  _392_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 5828 0 -1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL41860x32640
timestamp 1586547711
transform 1 0 8772 0 -1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1586547711
transform 1 0 8864 0 -1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL32660x32640
timestamp 1586547711
transform 1 0 6932 0 -1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL38180x32640
timestamp 1586547711
transform 1 0 8036 0 -1 7472
box 0 -48 736 592
use sky130_fd_sc_hd__a32o_4  _409_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 8956 0 -1 7472
box 0 -48 1564 592
use sky130_fd_sc_hd__decap_8  FILL50600x32640
timestamp 1586547711
transform 1 0 10520 0 -1 7472
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL59340x32640
timestamp 1586547711
transform 1 0 12268 0 -1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_880
timestamp 1586547711
transform 1 0 12360 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_887
timestamp 1586547711
transform 1 0 12544 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL56580x32640
timestamp 1586547711
transform 1 0 11716 0 -1 7472
box 0 -48 552 592
use sky130_fd_sc_hd__inv_4  _260_
timestamp 1586547711
transform 1 0 11256 0 -1 7472
box 0 -48 460 592
use sky130_fd_sc_hd__and2_4  _514_
timestamp 1586547711
transform 1 0 12728 0 -1 7472
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1586547711
transform 1 0 14476 0 -1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL70840x32640
timestamp 1586547711
transform 1 0 14568 0 -1 7472
box 0 -48 368 592
use sky130_fd_sc_hd__a211o_4  _508_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 14936 0 -1 7472
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL64860x32640
timestamp 1586547711
transform 1 0 13372 0 -1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILL84640x32640
timestamp 1586547711
transform 1 0 17328 0 -1 7472
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL79120x32640
timestamp 1586547711
transform 1 0 16224 0 -1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL87400x32640
timestamp 1586547711
transform 1 0 17880 0 -1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL88780x32640
timestamp 1586547711
transform 1 0 18156 0 -1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_823
timestamp 1586547711
transform 1 0 17696 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_785
timestamp 1586547711
transform 1 0 17972 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _486_
timestamp 1586547711
transform 1 0 18248 0 -1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL94760x32640
timestamp 1586547711
transform 1 0 19352 0 -1 7472
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_777
timestamp 1586547711
transform 1 0 20824 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_794
timestamp 1586547711
transform 1 0 21008 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1586547711
transform 1 0 20088 0 -1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL103960x32640
timestamp 1586547711
transform 1 0 21192 0 -1 7472
box 0 -48 368 592
use sky130_fd_sc_hd__inv_4  _482_
timestamp 1586547711
transform 1 0 21560 0 -1 7472
box 0 -48 460 592
use sky130_fd_sc_hd__and2_4  _481_
timestamp 1586547711
transform 1 0 20180 0 -1 7472
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL108100x32640
timestamp 1586547711
transform 1 0 22020 0 -1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL113620x32640
timestamp 1586547711
transform 1 0 23124 0 -1 7472
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL117300x32640
timestamp 1586547711
transform 1 0 23860 0 -1 7472
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL125120x32640
timestamp 1586547711
transform 1 0 25424 0 -1 7472
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_929
timestamp 1586547711
transform 1 0 24136 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1042
timestamp 1586547711
transform 1 0 24320 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1099
timestamp 1586547711
transform 1 0 24504 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1586547711
transform 1 0 25700 0 -1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL126960x32640
timestamp 1586547711
transform 1 0 25792 0 -1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL121440x32640
timestamp 1586547711
transform 1 0 24688 0 -1 7472
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1586547711
transform 1 0 26988 0 -1 7472
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL132480x32640
timestamp 1586547711
transform 1 0 26896 0 -1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1586547711
transform 1 0 400 0 -1 8560
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1586547711
transform 1 0 400 0 1 7472
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_68
timestamp 1586547711
transform 1 0 676 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_991
timestamp 1586547711
transform 1 0 860 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_460
timestamp 1586547711
transform 1 0 1412 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL3220x38080
timestamp 1586547711
transform 1 0 1044 0 -1 8560
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _343_
timestamp 1586547711
transform 1 0 1412 0 -1 8560
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL1380x35360
timestamp 1586547711
transform 1 0 676 0 1 7472
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_475
timestamp 1586547711
transform 1 0 1596 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_477
timestamp 1586547711
transform 1 0 1780 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL8280x38080
timestamp 1586547711
transform 1 0 2056 0 -1 8560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL7820x35360
timestamp 1586547711
transform 1 0 1964 0 1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL13800x38080
timestamp 1586547711
transform 1 0 3160 0 -1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1586547711
transform 1 0 3252 0 -1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL14720x38080
timestamp 1586547711
transform 1 0 3344 0 -1 8560
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILL13340x35360
timestamp 1586547711
transform 1 0 3068 0 1 7472
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL17020x35360
timestamp 1586547711
transform 1 0 3804 0 1 7472
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL16560x38080
timestamp 1586547711
transform 1 0 3712 0 -1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL17940x38080
timestamp 1586547711
transform 1 0 3988 0 -1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_601
timestamp 1586547711
transform 1 0 3804 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_192
timestamp 1586547711
transform 1 0 4080 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_209
timestamp 1586547711
transform 1 0 4264 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_317
timestamp 1586547711
transform 1 0 4448 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _294_
timestamp 1586547711
transform 1 0 4080 0 -1 8560
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL21160x35360
timestamp 1586547711
transform 1 0 4632 0 1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL25300x38080
timestamp 1586547711
transform 1 0 5460 0 -1 8560
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL21620x38080
timestamp 1586547711
transform 1 0 4724 0 -1 8560
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL27600x35360
timestamp 1586547711
transform 1 0 5920 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_517
timestamp 1586547711
transform 1 0 6196 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_606
timestamp 1586547711
transform 1 0 6380 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1149
timestamp 1586547711
transform 1 0 6564 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_318
timestamp 1586547711
transform 1 0 5736 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_320
timestamp 1586547711
transform 1 0 6104 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1586547711
transform 1 0 6012 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _295_
timestamp 1586547711
transform 1 0 5736 0 -1 8560
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL31740x38080
timestamp 1586547711
transform 1 0 6748 0 -1 8560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL29440x35360
timestamp 1586547711
transform 1 0 6288 0 1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL40940x38080
timestamp 1586547711
transform 1 0 8588 0 -1 8560
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL42320x35360
timestamp 1586547711
transform 1 0 8864 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1586547711
transform 1 0 8864 0 -1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL40480x35360
timestamp 1586547711
transform 1 0 8496 0 1 7472
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL34960x35360
timestamp 1586547711
transform 1 0 7392 0 1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL37260x38080
timestamp 1586547711
transform 1 0 7852 0 -1 8560
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_190
timestamp 1586547711
transform 1 0 8956 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1116
timestamp 1586547711
transform 1 0 9140 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _263_
timestamp 1586547711
transform 1 0 8956 0 -1 8560
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL45080x38080
timestamp 1586547711
transform 1 0 9416 0 -1 8560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL44620x35360
timestamp 1586547711
transform 1 0 9324 0 1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL50600x38080
timestamp 1586547711
transform 1 0 10520 0 -1 8560
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL50140x35360
timestamp 1586547711
transform 1 0 10428 0 1 7472
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL53820x35360
timestamp 1586547711
transform 1 0 11164 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL57500x35360
timestamp 1586547711
transform 1 0 11900 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_161
timestamp 1586547711
transform 1 0 11256 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_166
timestamp 1586547711
transform 1 0 11440 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_462
timestamp 1586547711
transform 1 0 11716 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_820
timestamp 1586547711
transform 1 0 11992 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1586547711
transform 1 0 11624 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL57500x38080
timestamp 1586547711
transform 1 0 11900 0 -1 8560
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _339_
timestamp 1586547711
transform 1 0 11256 0 -1 8560
box 0 -48 644 592
use sky130_fd_sc_hd__fill_1  FILL59340x38080
timestamp 1586547711
transform 1 0 12268 0 -1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_851
timestamp 1586547711
transform 1 0 12360 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_875
timestamp 1586547711
transform 1 0 12544 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_881
timestamp 1586547711
transform 1 0 12728 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_464
timestamp 1586547711
transform 1 0 12176 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__a211o_4  _521_
timestamp 1586547711
transform 1 0 12360 0 1 7472
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL62560x38080
timestamp 1586547711
transform 1 0 12912 0 -1 8560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILL68080x38080
timestamp 1586547711
transform 1 0 14016 0 -1 8560
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILL66240x35360
timestamp 1586547711
transform 1 0 13648 0 1 7472
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL69920x38080
timestamp 1586547711
transform 1 0 14384 0 -1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_877
timestamp 1586547711
transform 1 0 14568 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_848
timestamp 1586547711
transform 1 0 14568 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_780
timestamp 1586547711
transform 1 0 14752 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_818
timestamp 1586547711
transform 1 0 14936 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_845
timestamp 1586547711
transform 1 0 15120 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1586547711
transform 1 0 14476 0 -1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL69920x35360
timestamp 1586547711
transform 1 0 14384 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _502_
timestamp 1586547711
transform 1 0 14752 0 -1 8560
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL74520x35360
timestamp 1586547711
transform 1 0 15304 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_853
timestamp 1586547711
transform 1 0 15856 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_855
timestamp 1586547711
transform 1 0 16040 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL79120x35360
timestamp 1586547711
transform 1 0 16224 0 1 7472
box 0 -48 552 592
use sky130_fd_sc_hd__inv_4  _504_
timestamp 1586547711
transform 1 0 15396 0 1 7472
box 0 -48 460 592
use sky130_fd_sc_hd__fill_1  FILL81880x35360
timestamp 1586547711
transform 1 0 16776 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL84640x35360
timestamp 1586547711
transform 1 0 17328 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_832
timestamp 1586547711
transform 1 0 16868 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_829
timestamp 1586547711
transform 1 0 17052 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1586547711
transform 1 0 17236 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL82800x38080
timestamp 1586547711
transform 1 0 16960 0 -1 8560
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILL77280x38080
timestamp 1586547711
transform 1 0 15856 0 -1 8560
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_833
timestamp 1586547711
transform 1 0 18524 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1163
timestamp 1586547711
transform 1 0 18708 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_807
timestamp 1586547711
transform 1 0 17420 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_778
timestamp 1586547711
transform 1 0 17604 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_122
timestamp 1586547711
transform 1 0 17788 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__a32o_4  _495_
timestamp 1586547711
transform 1 0 17972 0 1 7472
box 0 -48 1564 592
use sky130_fd_sc_hd__nand2_4  _494_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 17696 0 -1 8560
box 0 -48 828 592
use sky130_fd_sc_hd__decap_12  FILL92460x38080
timestamp 1586547711
transform 1 0 18892 0 -1 8560
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL97980x38080
timestamp 1586547711
transform 1 0 19996 0 -1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_788
timestamp 1586547711
transform 1 0 20456 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1586547711
transform 1 0 20088 0 -1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL99360x35360
timestamp 1586547711
transform 1 0 20272 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL95680x35360
timestamp 1586547711
transform 1 0 19536 0 1 7472
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_773
timestamp 1586547711
transform 1 0 21284 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_784
timestamp 1586547711
transform 1 0 21468 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _480_
timestamp 1586547711
transform 1 0 20640 0 1 7472
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL98900x38080
timestamp 1586547711
transform 1 0 20180 0 -1 8560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL104420x38080
timestamp 1586547711
transform 1 0 21284 0 -1 8560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILL109940x38080
timestamp 1586547711
transform 1 0 22388 0 -1 8560
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILL112700x38080
timestamp 1586547711
transform 1 0 22940 0 -1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL111780x35360
timestamp 1586547711
transform 1 0 22756 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL112700x35360
timestamp 1586547711
transform 1 0 22940 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_237
timestamp 1586547711
transform 1 0 23032 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_645
timestamp 1586547711
transform 1 0 23032 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_96
timestamp 1586547711
transform 1 0 23216 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_230
timestamp 1586547711
transform 1 0 23400 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_233
timestamp 1586547711
transform 1 0 23584 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1586547711
transform 1 0 22848 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__o22ai_4  _422_
timestamp 1586547711
transform 1 0 23216 0 -1 8560
box 0 -48 1472 592
use sky130_fd_sc_hd__decap_12  FILL106260x35360
timestamp 1586547711
transform 1 0 21652 0 1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL125120x38080
timestamp 1586547711
transform 1 0 25424 0 -1 8560
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_633
timestamp 1586547711
transform 1 0 23768 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_97
timestamp 1586547711
transform 1 0 23952 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1586547711
transform 1 0 25700 0 -1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _269_
timestamp 1586547711
transform 1 0 25792 0 -1 8560
box 0 -48 460 592
use sky130_fd_sc_hd__dfrtp_4  _565_
timestamp 1586547711
transform 1 0 24136 0 1 7472
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_8  FILL121440x38080
timestamp 1586547711
transform 1 0 24688 0 -1 8560
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1586547711
transform 1 0 26988 0 -1 8560
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1586547711
transform 1 0 26988 0 1 7472
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_232
timestamp 1586547711
transform 1 0 26252 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1098
timestamp 1586547711
transform 1 0 26436 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL131100x35360
timestamp 1586547711
transform 1 0 26620 0 1 7472
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILL129260x38080
timestamp 1586547711
transform 1 0 26252 0 -1 8560
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1586547711
transform 1 0 400 0 1 8560
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_560
timestamp 1586547711
transform 1 0 1872 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_597
timestamp 1586547711
transform 1 0 2056 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_599
timestamp 1586547711
transform 1 0 2240 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL10120x40800
timestamp 1586547711
transform 1 0 2424 0 1 8560
box 0 -48 368 592
use sky130_fd_sc_hd__a21bo_4  _411_
timestamp 1586547711
transform 1 0 676 0 1 8560
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_1  FILL11960x40800
timestamp 1586547711
transform 1 0 2792 0 1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1153
timestamp 1586547711
transform 1 0 2884 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1125
timestamp 1586547711
transform 1 0 3068 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_519
timestamp 1586547711
transform 1 0 3252 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_513
timestamp 1586547711
transform 1 0 3436 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_336
timestamp 1586547711
transform 1 0 3620 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_204
timestamp 1586547711
transform 1 0 3804 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_319
timestamp 1586547711
transform 1 0 4632 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _362_
timestamp 1586547711
transform 1 0 3988 0 1 8560
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  FILL23000x40800
timestamp 1586547711
transform 1 0 5000 0 1 8560
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_509
timestamp 1586547711
transform 1 0 4816 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1108
timestamp 1586547711
transform 1 0 5276 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_605
timestamp 1586547711
transform 1 0 5460 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_400
timestamp 1586547711
transform 1 0 5644 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_334
timestamp 1586547711
transform 1 0 5828 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1586547711
transform 1 0 6012 0 1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _361_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 6104 0 1 8560
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  FILL34500x40800
timestamp 1586547711
transform 1 0 7300 0 1 8560
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_201
timestamp 1586547711
transform 1 0 6932 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1154
timestamp 1586547711
transform 1 0 7116 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_604
timestamp 1586547711
transform 1 0 7576 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_167
timestamp 1586547711
transform 1 0 8404 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_205
timestamp 1586547711
transform 1 0 8588 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL41860x40800
timestamp 1586547711
transform 1 0 8772 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _399_
timestamp 1586547711
transform 1 0 7760 0 1 8560
box 0 -48 644 592
use sky130_fd_sc_hd__fill_1  FILL52900x40800
timestamp 1586547711
transform 1 0 10980 0 1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_308
timestamp 1586547711
transform 1 0 8956 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_507
timestamp 1586547711
transform 1 0 9140 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1148
timestamp 1586547711
transform 1 0 9324 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL51060x40800
timestamp 1586547711
transform 1 0 10612 0 1 8560
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL45540x40800
timestamp 1586547711
transform 1 0 9508 0 1 8560
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL56580x40800
timestamp 1586547711
transform 1 0 11716 0 1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_159
timestamp 1586547711
transform 1 0 11072 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_327
timestamp 1586547711
transform 1 0 11256 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1132
timestamp 1586547711
transform 1 0 11440 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1136
timestamp 1586547711
transform 1 0 11808 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_879
timestamp 1586547711
transform 1 0 11992 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1586547711
transform 1 0 11624 0 1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_162
timestamp 1586547711
transform 1 0 12176 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_158
timestamp 1586547711
transform 1 0 12360 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _517_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 12544 0 1 8560
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA_878
timestamp 1586547711
transform 1 0 13924 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_844
timestamp 1586547711
transform 1 0 14108 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_842
timestamp 1586547711
transform 1 0 14292 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_206
timestamp 1586547711
transform 1 0 15120 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _501_
timestamp 1586547711
transform 1 0 14476 0 1 8560
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILL66700x40800
timestamp 1586547711
transform 1 0 13740 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL79120x40800
timestamp 1586547711
transform 1 0 16224 0 1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_826
timestamp 1586547711
transform 1 0 15304 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_817
timestamp 1586547711
transform 1 0 16316 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_821
timestamp 1586547711
transform 1 0 16500 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL81420x40800
timestamp 1586547711
transform 1 0 16684 0 1 8560
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1586547711
transform 1 0 17236 0 1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL84640x40800
timestamp 1586547711
transform 1 0 17328 0 1 8560
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILL75440x40800
timestamp 1586547711
transform 1 0 15488 0 1 8560
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_828
timestamp 1586547711
transform 1 0 17696 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_806
timestamp 1586547711
transform 1 0 18524 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_822
timestamp 1586547711
transform 1 0 18708 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_831
timestamp 1586547711
transform 1 0 18892 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_836
timestamp 1586547711
transform 1 0 19076 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_839
timestamp 1586547711
transform 1 0 19260 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _493_
timestamp 1586547711
transform 1 0 17880 0 1 8560
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL95220x40800
timestamp 1586547711
transform 1 0 19444 0 1 8560
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL102580x40800
timestamp 1586547711
transform 1 0 20916 0 1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_776
timestamp 1586547711
transform 1 0 21468 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL100740x40800
timestamp 1586547711
transform 1 0 20548 0 1 8560
box 0 -48 368 592
use sky130_fd_sc_hd__inv_4  _479_
timestamp 1586547711
transform 1 0 21008 0 1 8560
box 0 -48 460 592
use sky130_fd_sc_hd__decap_3  FILL107180x40800
timestamp 1586547711
transform 1 0 21836 0 1 8560
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_783
timestamp 1586547711
transform 1 0 21652 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_634
timestamp 1586547711
transform 1 0 22112 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_238
timestamp 1586547711
transform 1 0 22296 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_235
timestamp 1586547711
transform 1 0 22480 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_234
timestamp 1586547711
transform 1 0 22664 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_98
timestamp 1586547711
transform 1 0 22940 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1586547711
transform 1 0 22848 0 1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__or4_4  _478_
timestamp 1586547711
transform 1 0 23124 0 1 8560
box 0 -48 828 592
use sky130_fd_sc_hd__fill_1  FILL121440x40800
timestamp 1586547711
transform 1 0 24688 0 1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_231
timestamp 1586547711
transform 1 0 23952 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_646
timestamp 1586547711
transform 1 0 24136 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_653
timestamp 1586547711
transform 1 0 24320 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_775
timestamp 1586547711
transform 1 0 24504 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_236
timestamp 1586547711
transform 1 0 25240 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1100
timestamp 1586547711
transform 1 0 25424 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _270_
timestamp 1586547711
transform 1 0 24780 0 1 8560
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL126040x40800
timestamp 1586547711
transform 1 0 25608 0 1 8560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL131560x40800
timestamp 1586547711
transform 1 0 26712 0 1 8560
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1586547711
transform 1 0 26988 0 1 8560
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1586547711
transform 1 0 400 0 -1 9648
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL5980x43520
timestamp 1586547711
transform 1 0 1596 0 -1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_67
timestamp 1586547711
transform 1 0 676 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_617
timestamp 1586547711
transform 1 0 860 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_616
timestamp 1586547711
transform 1 0 1688 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL3220x43520
timestamp 1586547711
transform 1 0 1044 0 -1 9648
box 0 -48 552 592
use sky130_fd_sc_hd__or2_4  _396_
timestamp 1586547711
transform 1 0 1872 0 -1 9648
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL10580x43520
timestamp 1586547711
transform 1 0 2516 0 -1 9648
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL16560x43520
timestamp 1586547711
transform 1 0 3712 0 -1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1586547711
transform 1 0 3252 0 -1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL14720x43520
timestamp 1586547711
transform 1 0 3344 0 -1 9648
box 0 -48 368 592
use sky130_fd_sc_hd__a32o_4  _398_
timestamp 1586547711
transform 1 0 3804 0 -1 9648
box 0 -48 1564 592
use sky130_fd_sc_hd__o21a_4  _400_
timestamp 1586547711
transform 1 0 6104 0 -1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL24840x43520
timestamp 1586547711
transform 1 0 5368 0 -1 9648
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL39560x43520
timestamp 1586547711
transform 1 0 8312 0 -1 9648
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL41860x43520
timestamp 1586547711
transform 1 0 8772 0 -1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_415
timestamp 1586547711
transform 1 0 8588 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1586547711
transform 1 0 8864 0 -1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL34040x43520
timestamp 1586547711
transform 1 0 7208 0 -1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILL51520x43520
timestamp 1586547711
transform 1 0 10704 0 -1 9648
box 0 -48 368 592
use sky130_fd_sc_hd__and2_4  _359_
timestamp 1586547711
transform 1 0 8956 0 -1 9648
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL46000x43520
timestamp 1586547711
transform 1 0 9600 0 -1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__inv_4  _259_
timestamp 1586547711
transform 1 0 12452 0 -1 9648
box 0 -48 460 592
use sky130_fd_sc_hd__and2_4  _297_
timestamp 1586547711
transform 1 0 11072 0 -1 9648
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL62560x43520
timestamp 1586547711
transform 1 0 12912 0 -1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL56580x43520
timestamp 1586547711
transform 1 0 11716 0 -1 9648
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL68080x43520
timestamp 1586547711
transform 1 0 14016 0 -1 9648
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1142
timestamp 1586547711
transform 1 0 14292 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_847
timestamp 1586547711
transform 1 0 15212 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1586547711
transform 1 0 14476 0 -1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _516_
timestamp 1586547711
transform 1 0 14568 0 -1 9648
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_884
timestamp 1586547711
transform 1 0 15396 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1110
timestamp 1586547711
transform 1 0 17328 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL81880x43520
timestamp 1586547711
transform 1 0 16776 0 -1 9648
box 0 -48 552 592
use sky130_fd_sc_hd__inv_4  _492_
timestamp 1586547711
transform 1 0 16316 0 -1 9648
box 0 -48 460 592
use sky130_fd_sc_hd__decap_8  FILL75900x43520
timestamp 1586547711
transform 1 0 15580 0 -1 9648
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL91080x43520
timestamp 1586547711
transform 1 0 18616 0 -1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_840
timestamp 1586547711
transform 1 0 19352 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _498_
timestamp 1586547711
transform 1 0 18708 0 -1 9648
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL85560x43520
timestamp 1586547711
transform 1 0 17512 0 -1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1115
timestamp 1586547711
transform 1 0 20180 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL95680x43520
timestamp 1586547711
transform 1 0 19536 0 -1 9648
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1586547711
transform 1 0 20088 0 -1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL99820x43520
timestamp 1586547711
transform 1 0 20364 0 -1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL105340x43520
timestamp 1586547711
transform 1 0 21468 0 -1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL112700x43520
timestamp 1586547711
transform 1 0 22940 0 -1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL110860x43520
timestamp 1586547711
transform 1 0 22572 0 -1 9648
box 0 -48 368 592
use sky130_fd_sc_hd__o22ai_4  _423_
timestamp 1586547711
transform 1 0 23032 0 -1 9648
box 0 -48 1472 592
use sky130_fd_sc_hd__fill_1  FILL126040x43520
timestamp 1586547711
transform 1 0 25608 0 -1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_154
timestamp 1586547711
transform 1 0 24504 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_930
timestamp 1586547711
transform 1 0 24688 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1586547711
transform 1 0 25700 0 -1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL126960x43520
timestamp 1586547711
transform 1 0 25792 0 -1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL122360x43520
timestamp 1586547711
transform 1 0 24872 0 -1 9648
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1586547711
transform 1 0 26988 0 -1 9648
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL132480x43520
timestamp 1586547711
transform 1 0 26896 0 -1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1586547711
transform 1 0 400 0 1 9648
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL4140x46240
timestamp 1586547711
transform 1 0 1228 0 1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_584
timestamp 1586547711
transform 1 0 1320 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_521
timestamp 1586547711
transform 1 0 1504 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_458
timestamp 1586547711
transform 1 0 2516 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL1380x46240
timestamp 1586547711
transform 1 0 676 0 1 9648
box 0 -48 552 592
use sky130_fd_sc_hd__or4_4  _410_
timestamp 1586547711
transform 1 0 1688 0 1 9648
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA_554
timestamp 1586547711
transform 1 0 2884 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_532
timestamp 1586547711
transform 1 0 3068 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_459
timestamp 1586547711
transform 1 0 3252 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_435
timestamp 1586547711
transform 1 0 4080 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_454
timestamp 1586547711
transform 1 0 4264 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_494
timestamp 1586547711
transform 1 0 4448 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL21160x46240
timestamp 1586547711
transform 1 0 4632 0 1 9648
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _338_
timestamp 1586547711
transform 1 0 3436 0 1 9648
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILL11500x46240
timestamp 1586547711
transform 1 0 2700 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL23000x46240
timestamp 1586547711
transform 1 0 5000 0 1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL31280x46240
timestamp 1586547711
transform 1 0 6656 0 1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_518
timestamp 1586547711
transform 1 0 5092 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_520
timestamp 1586547711
transform 1 0 5276 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_522
timestamp 1586547711
transform 1 0 5460 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_397
timestamp 1586547711
transform 1 0 6748 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL28520x46240
timestamp 1586547711
transform 1 0 6104 0 1 9648
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1586547711
transform 1 0 6012 0 1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL26220x46240
timestamp 1586547711
transform 1 0 5644 0 1 9648
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILL37720x46240
timestamp 1586547711
transform 1 0 7944 0 1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_322
timestamp 1586547711
transform 1 0 7576 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_331
timestamp 1586547711
transform 1 0 7760 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_380
timestamp 1586547711
transform 1 0 8036 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_197
timestamp 1586547711
transform 1 0 8220 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_165
timestamp 1586547711
transform 1 0 8404 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _313_
timestamp 1586547711
transform 1 0 6932 0 1 9648
box 0 -48 644 592
use sky130_fd_sc_hd__and4_4  _318_
timestamp 1586547711
transform 1 0 8588 0 1 9648
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA_164
timestamp 1586547711
transform 1 0 9416 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_177
timestamp 1586547711
transform 1 0 9600 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_321
timestamp 1586547711
transform 1 0 9784 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1138
timestamp 1586547711
transform 1 0 9968 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1139
timestamp 1586547711
transform 1 0 10152 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL49680x46240
timestamp 1586547711
transform 1 0 10336 0 1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL58880x46240
timestamp 1586547711
transform 1 0 12176 0 1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_465
timestamp 1586547711
transform 1 0 11440 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_310
timestamp 1586547711
transform 1 0 12268 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_463
timestamp 1586547711
transform 1 0 12452 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_470
timestamp 1586547711
transform 1 0 12636 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_846
timestamp 1586547711
transform 1 0 12820 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_883
timestamp 1586547711
transform 1 0 13004 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1586547711
transform 1 0 11624 0 1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _340_
timestamp 1586547711
transform 1 0 11716 0 1 9648
box 0 -48 460 592
use sky130_fd_sc_hd__diode_2  ANTENNA_882
timestamp 1586547711
transform 1 0 13556 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_827
timestamp 1586547711
transform 1 0 13740 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_787
timestamp 1586547711
transform 1 0 13924 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_782
timestamp 1586547711
transform 1 0 14108 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_130
timestamp 1586547711
transform 1 0 14292 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL63940x46240
timestamp 1586547711
transform 1 0 13188 0 1 9648
box 0 -48 368 592
use sky130_fd_sc_hd__a32o_4  _520_
timestamp 1586547711
transform 1 0 14476 0 1 9648
box 0 -48 1564 592
use sky130_fd_sc_hd__fill_1  FILL81880x46240
timestamp 1586547711
transform 1 0 16776 0 1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_885
timestamp 1586547711
transform 1 0 16040 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_886
timestamp 1586547711
transform 1 0 16224 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_834
timestamp 1586547711
transform 1 0 16868 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_804
timestamp 1586547711
transform 1 0 17052 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_220
timestamp 1586547711
transform 1 0 17328 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1586547711
transform 1 0 17236 0 1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL80040x46240
timestamp 1586547711
transform 1 0 16408 0 1 9648
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILL86480x46240
timestamp 1586547711
transform 1 0 17696 0 1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL91080x46240
timestamp 1586547711
transform 1 0 18616 0 1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_800
timestamp 1586547711
transform 1 0 17512 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_798
timestamp 1586547711
transform 1 0 18248 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_803
timestamp 1586547711
transform 1 0 18432 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_779
timestamp 1586547711
transform 1 0 18708 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_124
timestamp 1586547711
transform 1 0 18892 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _485_
timestamp 1586547711
transform 1 0 17788 0 1 9648
box 0 -48 460 592
use sky130_fd_sc_hd__a32o_4  _499_
timestamp 1586547711
transform 1 0 19076 0 1 9648
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA_125
timestamp 1586547711
transform 1 0 20640 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_907
timestamp 1586547711
transform 1 0 20824 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1031
timestamp 1586547711
transform 1 0 21008 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL103960x46240
timestamp 1586547711
transform 1 0 21192 0 1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL112700x46240
timestamp 1586547711
transform 1 0 22940 0 1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_631
timestamp 1586547711
transform 1 0 23032 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_644
timestamp 1586547711
transform 1 0 23216 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_931
timestamp 1586547711
transform 1 0 23400 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_99
timestamp 1586547711
transform 1 0 23584 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL109480x46240
timestamp 1586547711
transform 1 0 22296 0 1 9648
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1586547711
transform 1 0 22848 0 1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _566_
timestamp 1586547711
transform 1 0 23768 0 1 9648
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1586547711
transform 1 0 26988 0 1 9648
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL127420x46240
timestamp 1586547711
transform 1 0 25884 0 1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1586547711
transform 1 0 400 0 -1 10736
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL5060x48960
timestamp 1586547711
transform 1 0 1412 0 -1 10736
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_598
timestamp 1586547711
transform 1 0 1688 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_558
timestamp 1586547711
transform 1 0 2056 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL7360x48960
timestamp 1586547711
transform 1 0 1872 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL1380x48960
timestamp 1586547711
transform 1 0 676 0 -1 10736
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL9200x48960
timestamp 1586547711
transform 1 0 2240 0 -1 10736
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL12880x48960
timestamp 1586547711
transform 1 0 2976 0 -1 10736
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_530
timestamp 1586547711
transform 1 0 4356 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_608
timestamp 1586547711
transform 1 0 4540 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1586547711
transform 1 0 3252 0 -1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL14720x48960
timestamp 1586547711
transform 1 0 3344 0 -1 10736
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _374_
timestamp 1586547711
transform 1 0 3712 0 -1 10736
box 0 -48 644 592
use sky130_fd_sc_hd__decap_4  FILL21620x48960
timestamp 1586547711
transform 1 0 4724 0 -1 10736
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _363_
timestamp 1586547711
transform 1 0 5092 0 -1 10736
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL26680x48960
timestamp 1586547711
transform 1 0 5736 0 -1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL34040x48960
timestamp 1586547711
transform 1 0 7208 0 -1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL41860x48960
timestamp 1586547711
transform 1 0 8772 0 -1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_514
timestamp 1586547711
transform 1 0 7300 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_214
timestamp 1586547711
transform 1 0 8588 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1586547711
transform 1 0 8864 0 -1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL32200x48960
timestamp 1586547711
transform 1 0 6840 0 -1 10736
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL35420x48960
timestamp 1586547711
transform 1 0 7484 0 -1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__and4_4  _308_
timestamp 1586547711
transform 1 0 8956 0 -1 10736
box 0 -48 828 592
use sky130_fd_sc_hd__decap_12  FILL46920x48960
timestamp 1586547711
transform 1 0 9784 0 -1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL52440x48960
timestamp 1586547711
transform 1 0 10888 0 -1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL57960x48960
timestamp 1586547711
transform 1 0 11992 0 -1 10736
box 0 -48 276 592
use sky130_fd_sc_hd__nor3_4  _518_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 12268 0 -1 10736
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_1  FILL69000x48960
timestamp 1586547711
transform 1 0 14200 0 -1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1141
timestamp 1586547711
transform 1 0 14292 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1586547711
transform 1 0 14476 0 -1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__a211o_4  _519_
timestamp 1586547711
transform 1 0 14568 0 -1 10736
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_8  FILL65320x48960
timestamp 1586547711
transform 1 0 13464 0 -1 10736
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILL82800x48960
timestamp 1586547711
transform 1 0 16960 0 -1 10736
box 0 -48 368 592
use sky130_fd_sc_hd__o22a_4  _496_
timestamp 1586547711
transform 1 0 17328 0 -1 10736
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL77280x48960
timestamp 1586547711
transform 1 0 15856 0 -1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL92920x48960
timestamp 1586547711
transform 1 0 18984 0 -1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_786
timestamp 1586547711
transform 1 0 19076 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_838
timestamp 1586547711
transform 1 0 19260 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1111
timestamp 1586547711
transform 1 0 19444 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL91080x48960
timestamp 1586547711
transform 1 0 18616 0 -1 10736
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILL97980x48960
timestamp 1586547711
transform 1 0 19996 0 -1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1586547711
transform 1 0 20088 0 -1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL96140x48960
timestamp 1586547711
transform 1 0 19628 0 -1 10736
box 0 -48 368 592
use sky130_fd_sc_hd__dfrtp_4  _554_
timestamp 1586547711
transform 1 0 20180 0 -1 10736
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_3  FILL115460x48960
timestamp 1586547711
transform 1 0 23492 0 -1 10736
box 0 -48 276 592
use sky130_fd_sc_hd__inv_4  _420_
timestamp 1586547711
transform 1 0 23032 0 -1 10736
box 0 -48 460 592
use sky130_fd_sc_hd__decap_8  FILL109480x48960
timestamp 1586547711
transform 1 0 22296 0 -1 10736
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL118680x48960
timestamp 1586547711
transform 1 0 24136 0 -1 10736
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1043
timestamp 1586547711
transform 1 0 23768 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1101
timestamp 1586547711
transform 1 0 23952 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1586547711
transform 1 0 25700 0 -1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _543_
timestamp 1586547711
transform 1 0 24412 0 -1 10736
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL126960x48960
timestamp 1586547711
transform 1 0 25792 0 -1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL122820x48960
timestamp 1586547711
transform 1 0 24964 0 -1 10736
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1586547711
transform 1 0 26988 0 -1 10736
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL132480x48960
timestamp 1586547711
transform 1 0 26896 0 -1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1586547711
transform 1 0 400 0 -1 11824
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1586547711
transform 1 0 400 0 1 10736
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL1380x54400
timestamp 1586547711
transform 1 0 676 0 -1 11824
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL1380x51680
timestamp 1586547711
transform 1 0 676 0 1 10736
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL5060x54400
timestamp 1586547711
transform 1 0 1412 0 -1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL5060x51680
timestamp 1586547711
transform 1 0 1412 0 1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_382
timestamp 1586547711
transform 1 0 1504 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_472
timestamp 1586547711
transform 1 0 1688 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_474
timestamp 1586547711
transform 1 0 1872 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _342_
timestamp 1586547711
transform 1 0 1504 0 -1 11824
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_545
timestamp 1586547711
transform 1 0 2148 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_610
timestamp 1586547711
transform 1 0 2332 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _375_
timestamp 1586547711
transform 1 0 2056 0 1 10736
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL10580x54400
timestamp 1586547711
transform 1 0 2516 0 -1 11824
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL14720x54400
timestamp 1586547711
transform 1 0 3344 0 -1 11824
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL13340x51680
timestamp 1586547711
transform 1 0 3068 0 1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_455
timestamp 1586547711
transform 1 0 2700 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_555
timestamp 1586547711
transform 1 0 2884 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_607
timestamp 1586547711
transform 1 0 3160 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_602
timestamp 1586547711
transform 1 0 3344 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1586547711
transform 1 0 3252 0 -1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL17020x54400
timestamp 1586547711
transform 1 0 3804 0 -1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL18400x54400
timestamp 1586547711
transform 1 0 4080 0 -1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_471
timestamp 1586547711
transform 1 0 3620 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_549
timestamp 1586547711
transform 1 0 3896 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_529
timestamp 1586547711
transform 1 0 3528 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_469
timestamp 1586547711
transform 1 0 3712 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _401_
timestamp 1586547711
transform 1 0 3896 0 1 10736
box 0 -48 828 592
use sky130_fd_sc_hd__and4_4  _365_
timestamp 1586547711
transform 1 0 4172 0 -1 11824
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA_185
timestamp 1586547711
transform 1 0 4724 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_217
timestamp 1586547711
transform 1 0 4908 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1122
timestamp 1586547711
transform 1 0 5092 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL23000x54400
timestamp 1586547711
transform 1 0 5000 0 -1 11824
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL24380x51680
timestamp 1586547711
transform 1 0 5276 0 1 10736
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_399
timestamp 1586547711
transform 1 0 6104 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_417
timestamp 1586547711
transform 1 0 6288 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_537
timestamp 1586547711
transform 1 0 6472 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1150
timestamp 1586547711
transform 1 0 6656 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1586547711
transform 1 0 6012 0 1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL26680x54400
timestamp 1586547711
transform 1 0 5736 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _367_
timestamp 1586547711
transform 1 0 5920 0 -1 11824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL33120x54400
timestamp 1586547711
transform 1 0 7024 0 -1 11824
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL32200x51680
timestamp 1586547711
transform 1 0 6840 0 1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_508
timestamp 1586547711
transform 1 0 7300 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_505
timestamp 1586547711
transform 1 0 6932 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_323
timestamp 1586547711
transform 1 0 7116 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL35420x54400
timestamp 1586547711
transform 1 0 7484 0 -1 11824
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILL41860x54400
timestamp 1586547711
transform 1 0 8772 0 -1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1109
timestamp 1586547711
transform 1 0 8036 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL39100x54400
timestamp 1586547711
transform 1 0 8220 0 -1 11824
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1586547711
transform 1 0 8864 0 -1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL40020x51680
timestamp 1586547711
transform 1 0 8404 0 1 10736
box 0 -48 736 592
use sky130_fd_sc_hd__a21o_4  _360_
timestamp 1586547711
transform 1 0 7300 0 1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_200
timestamp 1586547711
transform 1 0 9140 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_216
timestamp 1586547711
transform 1 0 9324 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_333
timestamp 1586547711
transform 1 0 9508 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_504
timestamp 1586547711
transform 1 0 9692 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL42780x54400
timestamp 1586547711
transform 1 0 8956 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _358_
timestamp 1586547711
transform 1 0 9140 0 -1 11824
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1147
timestamp 1586547711
transform 1 0 9876 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL48300x51680
timestamp 1586547711
transform 1 0 10060 0 1 10736
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL47840x54400
timestamp 1586547711
transform 1 0 9968 0 -1 11824
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL51060x51680
timestamp 1586547711
transform 1 0 10612 0 1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_170
timestamp 1586547711
transform 1 0 10704 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1144
timestamp 1586547711
transform 1 0 10888 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _261_
timestamp 1586547711
transform 1 0 10704 0 -1 11824
box 0 -48 460 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1133
timestamp 1586547711
transform 1 0 11440 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1586547711
transform 1 0 11624 0 1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL53360x51680
timestamp 1586547711
transform 1 0 11072 0 1 10736
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _307_
timestamp 1586547711
transform 1 0 11716 0 1 10736
box 0 -48 644 592
use sky130_fd_sc_hd__fill_1  FILL61180x54400
timestamp 1586547711
transform 1 0 12636 0 -1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_160
timestamp 1586547711
transform 1 0 12360 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_377
timestamp 1586547711
transform 1 0 12544 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_301
timestamp 1586547711
transform 1 0 12728 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_303
timestamp 1586547711
transform 1 0 12912 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL59340x54400
timestamp 1586547711
transform 1 0 12268 0 -1 11824
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _289_
timestamp 1586547711
transform 1 0 13096 0 1 10736
box 0 -48 644 592
use sky130_fd_sc_hd__inv_4  _290_
timestamp 1586547711
transform 1 0 12728 0 -1 11824
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL53820x54400
timestamp 1586547711
transform 1 0 11164 0 -1 11824
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1131
timestamp 1586547711
transform 1 0 13188 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1137
timestamp 1586547711
transform 1 0 13372 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_300
timestamp 1586547711
transform 1 0 13740 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1114
timestamp 1586547711
transform 1 0 13924 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL65780x54400
timestamp 1586547711
transform 1 0 13556 0 -1 11824
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1143
timestamp 1586547711
transform 1 0 14292 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1128
timestamp 1586547711
transform 1 0 14568 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_876
timestamp 1586547711
transform 1 0 14108 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_802
timestamp 1586547711
transform 1 0 14292 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1586547711
transform 1 0 14476 0 -1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL71760x54400
timestamp 1586547711
transform 1 0 14752 0 -1 11824
box 0 -48 368 592
use sky130_fd_sc_hd__or4_4  _515_
timestamp 1586547711
transform 1 0 14476 0 1 10736
box 0 -48 828 592
use sky130_fd_sc_hd__fill_1  FILL73600x54400
timestamp 1586547711
transform 1 0 15120 0 -1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_145
timestamp 1586547711
transform 1 0 15212 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL83720x51680
timestamp 1586547711
transform 1 0 17144 0 1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_912
timestamp 1586547711
transform 1 0 15396 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_302
timestamp 1586547711
transform 1 0 15304 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL80960x51680
timestamp 1586547711
transform 1 0 16592 0 1 10736
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1586547711
transform 1 0 17236 0 1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL75900x54400
timestamp 1586547711
transform 1 0 15580 0 -1 11824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL81420x54400
timestamp 1586547711
transform 1 0 16684 0 -1 11824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL75440x51680
timestamp 1586547711
transform 1 0 15488 0 1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL84640x51680
timestamp 1586547711
transform 1 0 17328 0 1 10736
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_837
timestamp 1586547711
transform 1 0 18064 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_835
timestamp 1586547711
transform 1 0 18248 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_830
timestamp 1586547711
transform 1 0 19260 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__nand2_4  _497_
timestamp 1586547711
transform 1 0 18432 0 1 10736
box 0 -48 828 592
use sky130_fd_sc_hd__decap_12  FILL86940x54400
timestamp 1586547711
transform 1 0 17788 0 -1 11824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL92460x54400
timestamp 1586547711
transform 1 0 18892 0 -1 11824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL95220x51680
timestamp 1586547711
transform 1 0 19444 0 1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL97980x54400
timestamp 1586547711
transform 1 0 19996 0 -1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL100740x51680
timestamp 1586547711
transform 1 0 20548 0 1 10736
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1586547711
transform 1 0 20088 0 -1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _531_
timestamp 1586547711
transform 1 0 21100 0 1 10736
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL98900x54400
timestamp 1586547711
transform 1 0 20180 0 -1 11824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL104420x54400
timestamp 1586547711
transform 1 0 21284 0 -1 11824
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_142
timestamp 1586547711
transform 1 0 21652 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_906
timestamp 1586547711
transform 1 0 21836 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL109940x54400
timestamp 1586547711
transform 1 0 22388 0 -1 11824
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL108100x51680
timestamp 1586547711
transform 1 0 22020 0 1 10736
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL112700x54400
timestamp 1586547711
transform 1 0 22940 0 -1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL115920x54400
timestamp 1586547711
transform 1 0 23584 0 -1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL111780x51680
timestamp 1586547711
transform 1 0 22756 0 1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_639
timestamp 1586547711
transform 1 0 23032 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_893
timestamp 1586547711
transform 1 0 23676 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1586547711
transform 1 0 22848 0 1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL114080x54400
timestamp 1586547711
transform 1 0 23216 0 -1 11824
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL112700x51680
timestamp 1586547711
transform 1 0 22940 0 1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1024
timestamp 1586547711
transform 1 0 23860 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1075
timestamp 1586547711
transform 1 0 24044 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_135
timestamp 1586547711
transform 1 0 24412 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_892
timestamp 1586547711
transform 1 0 24596 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL118220x51680
timestamp 1586547711
transform 1 0 24044 0 1 10736
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL119140x54400
timestamp 1586547711
transform 1 0 24228 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _524_
timestamp 1586547711
transform 1 0 24412 0 -1 11824
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1586547711
transform 1 0 25700 0 -1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL122820x54400
timestamp 1586547711
transform 1 0 24964 0 -1 11824
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILL126960x54400
timestamp 1586547711
transform 1 0 25792 0 -1 11824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL121900x51680
timestamp 1586547711
transform 1 0 24780 0 1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1586547711
transform 1 0 26988 0 -1 11824
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1586547711
transform 1 0 26988 0 1 10736
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL132480x54400
timestamp 1586547711
transform 1 0 26896 0 -1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL127420x51680
timestamp 1586547711
transform 1 0 25884 0 1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1586547711
transform 1 0 400 0 1 11824
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL7820x57120
timestamp 1586547711
transform 1 0 1964 0 1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_567
timestamp 1586547711
transform 1 0 1228 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_557
timestamp 1586547711
transform 1 0 1412 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_476
timestamp 1586547711
transform 1 0 1596 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_535
timestamp 1586547711
transform 1 0 1780 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL1380x57120
timestamp 1586547711
transform 1 0 676 0 1 11824
box 0 -48 552 592
use sky130_fd_sc_hd__or4_4  _402_
timestamp 1586547711
transform 1 0 2056 0 1 11824
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA_503
timestamp 1586547711
transform 1 0 2884 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_215
timestamp 1586547711
transform 1 0 3252 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_198
timestamp 1586547711
transform 1 0 3436 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_182
timestamp 1586547711
transform 1 0 4448 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_526
timestamp 1586547711
transform 1 0 4632 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL13340x57120
timestamp 1586547711
transform 1 0 3068 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _341_
timestamp 1586547711
transform 1 0 3620 0 1 11824
box 0 -48 828 592
use sky130_fd_sc_hd__fill_1  FILL23920x57120
timestamp 1586547711
transform 1 0 5184 0 1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_531
timestamp 1586547711
transform 1 0 4816 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_533
timestamp 1586547711
transform 1 0 5000 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_538
timestamp 1586547711
transform 1 0 5276 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_534
timestamp 1586547711
transform 1 0 5460 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_523
timestamp 1586547711
transform 1 0 5644 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_486
timestamp 1586547711
transform 1 0 5828 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1586547711
transform 1 0 6012 0 1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__or4_4  _368_
timestamp 1586547711
transform 1 0 6104 0 1 11824
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA_515
timestamp 1586547711
transform 1 0 6932 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_539
timestamp 1586547711
transform 1 0 7116 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_556
timestamp 1586547711
transform 1 0 7300 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_579
timestamp 1586547711
transform 1 0 7484 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_525
timestamp 1586547711
transform 1 0 7668 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_468
timestamp 1586547711
transform 1 0 7852 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_184
timestamp 1586547711
transform 1 0 8864 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _364_
timestamp 1586547711
transform 1 0 8036 0 1 11824
box 0 -48 828 592
use sky130_fd_sc_hd__fill_1  FILL52440x57120
timestamp 1586547711
transform 1 0 10888 0 1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_181
timestamp 1586547711
transform 1 0 10980 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL43240x57120
timestamp 1586547711
transform 1 0 9048 0 1 11824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL48760x57120
timestamp 1586547711
transform 1 0 10152 0 1 11824
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL55660x57120
timestamp 1586547711
transform 1 0 11532 0 1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_332
timestamp 1586547711
transform 1 0 11164 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_431
timestamp 1586547711
transform 1 0 11348 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_433
timestamp 1586547711
transform 1 0 11716 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1586547711
transform 1 0 11624 0 1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL57500x57120
timestamp 1586547711
transform 1 0 11900 0 1 11824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL63020x57120
timestamp 1586547711
transform 1 0 13004 0 1 11824
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_913
timestamp 1586547711
transform 1 0 13924 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_131
timestamp 1586547711
transform 1 0 14108 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL66700x57120
timestamp 1586547711
transform 1 0 13740 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _557_
timestamp 1586547711
transform 1 0 14292 0 1 11824
box 0 -48 2116 592
use sky130_fd_sc_hd__fill_1  FILL83720x57120
timestamp 1586547711
transform 1 0 17144 0 1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL84640x57120
timestamp 1586547711
transform 1 0 17328 0 1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1586547711
transform 1 0 17236 0 1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL80040x57120
timestamp 1586547711
transform 1 0 16408 0 1 11824
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_771
timestamp 1586547711
transform 1 0 17420 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_815
timestamp 1586547711
transform 1 0 17604 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_816
timestamp 1586547711
transform 1 0 17788 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL87860x57120
timestamp 1586547711
transform 1 0 17972 0 1 11824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL93380x57120
timestamp 1586547711
transform 1 0 19076 0 1 11824
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL104420x57120
timestamp 1586547711
transform 1 0 21284 0 1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_740
timestamp 1586547711
transform 1 0 20180 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_741
timestamp 1586547711
transform 1 0 20364 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_292
timestamp 1586547711
transform 1 0 21376 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_732
timestamp 1586547711
transform 1 0 21560 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL100740x57120
timestamp 1586547711
transform 1 0 20548 0 1 11824
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_734
timestamp 1586547711
transform 1 0 21744 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_648
timestamp 1586547711
transform 1 0 22480 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL107640x57120
timestamp 1586547711
transform 1 0 21928 0 1 11824
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILL112700x57120
timestamp 1586547711
transform 1 0 22940 0 1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL115000x57120
timestamp 1586547711
transform 1 0 23400 0 1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_265
timestamp 1586547711
transform 1 0 22664 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_110
timestamp 1586547711
transform 1 0 23032 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_249
timestamp 1586547711
transform 1 0 23216 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_111
timestamp 1586547711
transform 1 0 23492 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1586547711
transform 1 0 22848 0 1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _547_
timestamp 1586547711
transform 1 0 23676 0 1 11824
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_12  FILL126960x57120
timestamp 1586547711
transform 1 0 25792 0 1 11824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1586547711
transform 1 0 26988 0 1 11824
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL132480x57120
timestamp 1586547711
transform 1 0 26896 0 1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1586547711
transform 1 0 400 0 -1 12912
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_609
timestamp 1586547711
transform 1 0 2240 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _380_
timestamp 1586547711
transform 1 0 1596 0 -1 12912
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILL5060x59840
timestamp 1586547711
transform 1 0 1412 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL1380x59840
timestamp 1586547711
transform 1 0 676 0 -1 12912
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL10120x59840
timestamp 1586547711
transform 1 0 2424 0 -1 12912
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL14720x59840
timestamp 1586547711
transform 1 0 3344 0 -1 12912
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL13800x59840
timestamp 1586547711
transform 1 0 3160 0 -1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_466
timestamp 1586547711
transform 1 0 3620 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_493
timestamp 1586547711
transform 1 0 3988 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1586547711
transform 1 0 3252 0 -1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _366_
timestamp 1586547711
transform 1 0 4172 0 -1 12912
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILL17020x59840
timestamp 1586547711
transform 1 0 3804 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_580
timestamp 1586547711
transform 1 0 5736 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_543
timestamp 1586547711
transform 1 0 6748 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL25760x59840
timestamp 1586547711
transform 1 0 5552 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _387_
timestamp 1586547711
transform 1 0 5920 0 -1 12912
box 0 -48 828 592
use sky130_fd_sc_hd__decap_8  FILL22080x59840
timestamp 1586547711
transform 1 0 4816 0 -1 12912
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILL32660x59840
timestamp 1586547711
transform 1 0 6932 0 -1 12912
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_328
timestamp 1586547711
transform 1 0 7300 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_337
timestamp 1586547711
transform 1 0 7484 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_516
timestamp 1586547711
transform 1 0 7668 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_524
timestamp 1586547711
transform 1 0 7852 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_577
timestamp 1586547711
transform 1 0 8036 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1121
timestamp 1586547711
transform 1 0 8220 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL40020x59840
timestamp 1586547711
transform 1 0 8404 0 -1 12912
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILL41860x59840
timestamp 1586547711
transform 1 0 8772 0 -1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1586547711
transform 1 0 8864 0 -1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILL42780x59840
timestamp 1586547711
transform 1 0 8956 0 -1 12912
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL51520x59840
timestamp 1586547711
transform 1 0 10704 0 -1 12912
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_561
timestamp 1586547711
transform 1 0 9232 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1117
timestamp 1586547711
transform 1 0 9784 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL45080x59840
timestamp 1586547711
transform 1 0 9416 0 -1 12912
box 0 -48 368 592
use sky130_fd_sc_hd__a21o_4  _325_
timestamp 1586547711
transform 1 0 10980 0 -1 12912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL47840x59840
timestamp 1586547711
transform 1 0 9968 0 -1 12912
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_430
timestamp 1586547711
transform 1 0 12084 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL63020x59840
timestamp 1586547711
transform 1 0 13004 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL59340x59840
timestamp 1586547711
transform 1 0 12268 0 -1 12912
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL73600x59840
timestamp 1586547711
transform 1 0 15120 0 -1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_997
timestamp 1586547711
transform 1 0 13188 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1034
timestamp 1586547711
transform 1 0 14292 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL70840x59840
timestamp 1586547711
transform 1 0 14568 0 -1 12912
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1586547711
transform 1 0 14476 0 -1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL68540x59840
timestamp 1586547711
transform 1 0 14108 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _534_
timestamp 1586547711
transform 1 0 15212 0 -1 12912
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL64860x59840
timestamp 1586547711
transform 1 0 13372 0 -1 12912
box 0 -48 736 592
use sky130_fd_sc_hd__decap_6  FILL82340x59840
timestamp 1586547711
transform 1 0 16868 0 -1 12912
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL76820x59840
timestamp 1586547711
transform 1 0 15764 0 -1 12912
box 0 -48 1104 592
use sky130_fd_sc_hd__or2_4  _491_
timestamp 1586547711
transform 1 0 17420 0 -1 12912
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL88320x59840
timestamp 1586547711
transform 1 0 18064 0 -1 12912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL93840x59840
timestamp 1586547711
transform 1 0 19168 0 -1 12912
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_735
timestamp 1586547711
transform 1 0 20640 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_739
timestamp 1586547711
transform 1 0 20824 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1586547711
transform 1 0 20088 0 -1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL103040x59840
timestamp 1586547711
transform 1 0 21008 0 -1 12912
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL97520x59840
timestamp 1586547711
transform 1 0 19904 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _465_
timestamp 1586547711
transform 1 0 20180 0 -1 12912
box 0 -48 460 592
use sky130_fd_sc_hd__nor2_4  _462_
timestamp 1586547711
transform 1 0 21376 0 -1 12912
box 0 -48 828 592
use sky130_fd_sc_hd__fill_1  FILL112700x59840
timestamp 1586547711
transform 1 0 22940 0 -1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__o22ai_4  _440_
timestamp 1586547711
transform 1 0 23032 0 -1 12912
box 0 -48 1472 592
use sky130_fd_sc_hd__decap_8  FILL109020x59840
timestamp 1586547711
transform 1 0 22204 0 -1 12912
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL126040x59840
timestamp 1586547711
transform 1 0 25608 0 -1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1586547711
transform 1 0 25700 0 -1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL120520x59840
timestamp 1586547711
transform 1 0 24504 0 -1 12912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL126960x59840
timestamp 1586547711
transform 1 0 25792 0 -1 12912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1586547711
transform 1 0 26988 0 -1 12912
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL132480x59840
timestamp 1586547711
transform 1 0 26896 0 -1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1586547711
transform 1 0 400 0 1 12912
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_582
timestamp 1586547711
transform 1 0 1228 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_536
timestamp 1586547711
transform 1 0 1412 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_495
timestamp 1586547711
transform 1 0 1596 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_491
timestamp 1586547711
transform 1 0 1780 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL1380x62560
timestamp 1586547711
transform 1 0 676 0 1 12912
box 0 -48 552 592
use sky130_fd_sc_hd__or2_4  _353_
timestamp 1586547711
transform 1 0 1964 0 1 12912
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  FILL12880x62560
timestamp 1586547711
transform 1 0 2976 0 1 12912
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_473
timestamp 1586547711
transform 1 0 2608 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_488
timestamp 1586547711
transform 1 0 2792 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_550
timestamp 1586547711
transform 1 0 3252 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_547
timestamp 1586547711
transform 1 0 3436 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_487
timestamp 1586547711
transform 1 0 3620 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_467
timestamp 1586547711
transform 1 0 3804 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_199
timestamp 1586547711
transform 1 0 3988 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _352_
timestamp 1586547711
transform 1 0 4172 0 1 12912
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  FILL23920x62560
timestamp 1586547711
transform 1 0 5184 0 1 12912
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_183
timestamp 1586547711
transform 1 0 5000 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1151
timestamp 1586547711
transform 1 0 5460 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_546
timestamp 1586547711
transform 1 0 5644 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_335
timestamp 1586547711
transform 1 0 5828 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1586547711
transform 1 0 6012 0 1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _370_
timestamp 1586547711
transform 1 0 6104 0 1 12912
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA_218
timestamp 1586547711
transform 1 0 6932 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_210
timestamp 1586547711
transform 1 0 7116 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_173
timestamp 1586547711
transform 1 0 7300 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_193
timestamp 1586547711
transform 1 0 7484 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_429
timestamp 1586547711
transform 1 0 8496 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_506
timestamp 1586547711
transform 1 0 8864 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL41400x62560
timestamp 1586547711
transform 1 0 8680 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _386_
timestamp 1586547711
transform 1 0 7668 0 1 12912
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA_357
timestamp 1586547711
transform 1 0 9048 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_172
timestamp 1586547711
transform 1 0 10060 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_305
timestamp 1586547711
transform 1 0 10244 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_324
timestamp 1586547711
transform 1 0 10428 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1103
timestamp 1586547711
transform 1 0 10612 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_427
timestamp 1586547711
transform 1 0 10980 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL51980x62560
timestamp 1586547711
transform 1 0 10796 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__or3_4  _376_
timestamp 1586547711
transform 1 0 9232 0 1 12912
box 0 -48 828 592
use sky130_fd_sc_hd__fill_1  FILL55660x62560
timestamp 1586547711
transform 1 0 11532 0 1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_355
timestamp 1586547711
transform 1 0 11164 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_326
timestamp 1586547711
transform 1 0 11348 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1586547711
transform 1 0 11624 0 1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _324_
timestamp 1586547711
transform 1 0 11716 0 1 12912
box 0 -48 644 592
use sky130_fd_sc_hd__fill_1  FILL61640x62560
timestamp 1586547711
transform 1 0 12728 0 1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_363
timestamp 1586547711
transform 1 0 12360 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_428
timestamp 1586547711
transform 1 0 12544 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_90
timestamp 1586547711
transform 1 0 12820 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_44
timestamp 1586547711
transform 1 0 13004 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _327_
timestamp 1586547711
transform 1 0 13188 0 1 12912
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_12  FILL69920x62560
timestamp 1586547711
transform 1 0 14384 0 1 12912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL75440x62560
timestamp 1586547711
transform 1 0 15488 0 1 12912
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_207
timestamp 1586547711
transform 1 0 15764 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1102
timestamp 1586547711
transform 1 0 15948 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1586547711
transform 1 0 17236 0 1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _490_
timestamp 1586547711
transform 1 0 17328 0 1 12912
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL78660x62560
timestamp 1586547711
transform 1 0 16132 0 1 12912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL95220x62560
timestamp 1586547711
transform 1 0 19444 0 1 12912
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_813
timestamp 1586547711
transform 1 0 17788 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_814
timestamp 1586547711
transform 1 0 17972 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_726
timestamp 1586547711
transform 1 0 18524 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_745
timestamp 1586547711
transform 1 0 18708 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_766
timestamp 1586547711
transform 1 0 18892 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_770
timestamp 1586547711
transform 1 0 19076 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_772
timestamp 1586547711
transform 1 0 19260 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL88780x62560
timestamp 1586547711
transform 1 0 18156 0 1 12912
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_808
timestamp 1586547711
transform 1 0 19720 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_743
timestamp 1586547711
transform 1 0 19904 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_736
timestamp 1586547711
transform 1 0 20088 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_733
timestamp 1586547711
transform 1 0 20272 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_293
timestamp 1586547711
transform 1 0 20456 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__a211o_4  _464_
timestamp 1586547711
transform 1 0 20640 0 1 12912
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_3  FILL114540x62560
timestamp 1586547711
transform 1 0 23308 0 1 12912
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_295
timestamp 1586547711
transform 1 0 21928 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_729
timestamp 1586547711
transform 1 0 22112 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_737
timestamp 1586547711
transform 1 0 22296 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_702
timestamp 1586547711
transform 1 0 22940 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_706
timestamp 1586547711
transform 1 0 23124 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_701
timestamp 1586547711
transform 1 0 23584 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1586547711
transform 1 0 22848 0 1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL110400x62560
timestamp 1586547711
transform 1 0 22480 0 1 12912
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_250
timestamp 1586547711
transform 1 0 24412 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_266
timestamp 1586547711
transform 1 0 24596 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_264
timestamp 1586547711
transform 1 0 25608 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1073
timestamp 1586547711
transform 1 0 25792 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL121900x62560
timestamp 1586547711
transform 1 0 24780 0 1 12912
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _451_
timestamp 1586547711
transform 1 0 23768 0 1 12912
box 0 -48 644 592
use sky130_fd_sc_hd__inv_4  _276_
timestamp 1586547711
transform 1 0 25148 0 1 12912
box 0 -48 460 592
use sky130_fd_sc_hd__decap_3  FILL131560x62560
timestamp 1586547711
transform 1 0 26712 0 1 12912
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1586547711
transform 1 0 26988 0 1 12912
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL127880x62560
timestamp 1586547711
transform 1 0 25976 0 1 12912
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1586547711
transform 1 0 400 0 -1 14000
box 0 -48 276 592
use sky130_fd_sc_hd__or2_4  _389_
timestamp 1586547711
transform 1 0 1780 0 -1 14000
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL1380x65280
timestamp 1586547711
transform 1 0 676 0 -1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL10120x65280
timestamp 1586547711
transform 1 0 2424 0 -1 14000
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL13800x65280
timestamp 1586547711
transform 1 0 3160 0 -1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL17480x65280
timestamp 1586547711
transform 1 0 3896 0 -1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1107
timestamp 1586547711
transform 1 0 4632 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL14720x65280
timestamp 1586547711
transform 1 0 3344 0 -1 14000
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1586547711
transform 1 0 3252 0 -1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _371_
timestamp 1586547711
transform 1 0 3988 0 -1 14000
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1123
timestamp 1586547711
transform 1 0 6104 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL27600x65280
timestamp 1586547711
transform 1 0 5920 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL22080x65280
timestamp 1586547711
transform 1 0 4816 0 -1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL29440x65280
timestamp 1586547711
transform 1 0 6288 0 -1 14000
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL33120x65280
timestamp 1586547711
transform 1 0 7024 0 -1 14000
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_578
timestamp 1586547711
transform 1 0 8128 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL39560x65280
timestamp 1586547711
transform 1 0 8312 0 -1 14000
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1586547711
transform 1 0 8864 0 -1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _298_
timestamp 1586547711
transform 1 0 7300 0 -1 14000
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  FILL42780x65280
timestamp 1586547711
transform 1 0 8956 0 -1 14000
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_527
timestamp 1586547711
transform 1 0 9232 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL45080x65280
timestamp 1586547711
transform 1 0 9416 0 -1 14000
box 0 -48 368 592
use sky130_fd_sc_hd__and4_4  _296_
timestamp 1586547711
transform 1 0 9784 0 -1 14000
box 0 -48 828 592
use sky130_fd_sc_hd__decap_8  FILL51060x65280
timestamp 1586547711
transform 1 0 10612 0 -1 14000
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL63480x65280
timestamp 1586547711
transform 1 0 13096 0 -1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_385
timestamp 1586547711
transform 1 0 11992 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1106
timestamp 1586547711
transform 1 0 12176 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _323_
timestamp 1586547711
transform 1 0 11348 0 -1 14000
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL59800x65280
timestamp 1586547711
transform 1 0 12360 0 -1 14000
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_432
timestamp 1586547711
transform 1 0 13188 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1586547711
transform 1 0 14476 0 -1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL64860x65280
timestamp 1586547711
transform 1 0 13372 0 -1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL70840x65280
timestamp 1586547711
transform 1 0 14568 0 -1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL76360x65280
timestamp 1586547711
transform 1 0 15672 0 -1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL84640x65280
timestamp 1586547711
transform 1 0 17328 0 -1 14000
box 0 -48 368 592
use sky130_fd_sc_hd__inv_4  _264_
timestamp 1586547711
transform 1 0 15764 0 -1 14000
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL79120x65280
timestamp 1586547711
transform 1 0 16224 0 -1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL87400x65280
timestamp 1586547711
transform 1 0 17880 0 -1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_809
timestamp 1586547711
transform 1 0 17696 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_765
timestamp 1586547711
transform 1 0 17972 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL88780x65280
timestamp 1586547711
transform 1 0 18156 0 -1 14000
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILL94760x65280
timestamp 1586547711
transform 1 0 19352 0 -1 14000
box 0 -48 368 592
use sky130_fd_sc_hd__or4_4  _477_
timestamp 1586547711
transform 1 0 18524 0 -1 14000
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA_744
timestamp 1586547711
transform 1 0 19720 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_738
timestamp 1586547711
transform 1 0 20824 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL103040x65280
timestamp 1586547711
transform 1 0 21008 0 -1 14000
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1586547711
transform 1 0 20088 0 -1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _487_
timestamp 1586547711
transform 1 0 20180 0 -1 14000
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILL97520x65280
timestamp 1586547711
transform 1 0 19904 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _463_
timestamp 1586547711
transform 1 0 21560 0 -1 14000
box 0 -48 644 592
use sky130_fd_sc_hd__fill_1  FILL109020x65280
timestamp 1586547711
transform 1 0 22204 0 -1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL112240x65280
timestamp 1586547711
transform 1 0 22848 0 -1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_731
timestamp 1586547711
transform 1 0 22296 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_728
timestamp 1586547711
transform 1 0 23400 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1074
timestamp 1586547711
transform 1 0 23584 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL110400x65280
timestamp 1586547711
transform 1 0 22480 0 -1 14000
box 0 -48 368 592
use sky130_fd_sc_hd__inv_4  _452_
timestamp 1586547711
transform 1 0 22940 0 -1 14000
box 0 -48 460 592
use sky130_fd_sc_hd__fill_1  FILL126040x65280
timestamp 1586547711
transform 1 0 25608 0 -1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1586547711
transform 1 0 25700 0 -1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL116840x65280
timestamp 1586547711
transform 1 0 23768 0 -1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL126960x65280
timestamp 1586547711
transform 1 0 25792 0 -1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL122360x65280
timestamp 1586547711
transform 1 0 24872 0 -1 14000
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1586547711
transform 1 0 26988 0 -1 14000
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL132480x65280
timestamp 1586547711
transform 1 0 26896 0 -1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1586547711
transform 1 0 400 0 1 14000
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_588
timestamp 1586547711
transform 1 0 1228 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_586
timestamp 1586547711
transform 1 0 1412 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_583
timestamp 1586547711
transform 1 0 1596 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_544
timestamp 1586547711
transform 1 0 1780 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL1380x68000
timestamp 1586547711
transform 1 0 676 0 1 14000
box 0 -48 552 592
use sky130_fd_sc_hd__or4_4  _391_
timestamp 1586547711
transform 1 0 1964 0 1 14000
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA_502
timestamp 1586547711
transform 1 0 2792 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_585
timestamp 1586547711
transform 1 0 2976 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_551
timestamp 1586547711
transform 1 0 3160 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_203
timestamp 1586547711
transform 1 0 3344 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_511
timestamp 1586547711
transform 1 0 3528 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_540
timestamp 1586547711
transform 1 0 3712 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _372_
timestamp 1586547711
transform 1 0 3896 0 1 14000
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA_501
timestamp 1586547711
transform 1 0 4724 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL22540x68000
timestamp 1586547711
transform 1 0 4908 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_178
timestamp 1586547711
transform 1 0 5092 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_212
timestamp 1586547711
transform 1 0 5276 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_330
timestamp 1586547711
transform 1 0 5460 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_394
timestamp 1586547711
transform 1 0 5644 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1119
timestamp 1586547711
transform 1 0 5828 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1586547711
transform 1 0 6012 0 1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL28520x68000
timestamp 1586547711
transform 1 0 6104 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_528
timestamp 1586547711
transform 1 0 6288 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_510
timestamp 1586547711
transform 1 0 6472 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_408
timestamp 1586547711
transform 1 0 6656 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_383
timestamp 1586547711
transform 1 0 6840 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_366
timestamp 1586547711
transform 1 0 7024 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_339
timestamp 1586547711
transform 1 0 8036 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_548
timestamp 1586547711
transform 1 0 8220 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_562
timestamp 1586547711
transform 1 0 8404 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_563
timestamp 1586547711
transform 1 0 8588 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_576
timestamp 1586547711
transform 1 0 8772 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _385_
timestamp 1586547711
transform 1 0 7208 0 1 14000
box 0 -48 828 592
use sky130_fd_sc_hd__fill_1  FILL52440x68000
timestamp 1586547711
transform 1 0 10888 0 1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_325
timestamp 1586547711
transform 1 0 8956 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_338
timestamp 1586547711
transform 1 0 9140 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_340
timestamp 1586547711
transform 1 0 9324 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_306
timestamp 1586547711
transform 1 0 9508 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_211
timestamp 1586547711
transform 1 0 9692 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_175
timestamp 1586547711
transform 1 0 10704 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_379
timestamp 1586547711
transform 1 0 10980 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _302_
timestamp 1586547711
transform 1 0 9876 0 1 14000
box 0 -48 828 592
use sky130_fd_sc_hd__fill_1  FILL55660x68000
timestamp 1586547711
transform 1 0 11532 0 1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_378
timestamp 1586547711
transform 1 0 11164 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_213
timestamp 1586547711
transform 1 0 11348 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_196
timestamp 1586547711
transform 1 0 12544 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1120
timestamp 1586547711
transform 1 0 12728 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1146
timestamp 1586547711
transform 1 0 12912 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1586547711
transform 1 0 11624 0 1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL63480x68000
timestamp 1586547711
transform 1 0 13096 0 1 14000
box 0 -48 368 592
use sky130_fd_sc_hd__or4_4  _309_
timestamp 1586547711
transform 1 0 11716 0 1 14000
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1264
timestamp 1586547711
transform 1 0 13832 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1279
timestamp 1586547711
transform 1 0 14016 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[4\].id.delaybuf0
timestamp 1586547711
transform 1 0 13464 0 1 14000
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL69000x68000
timestamp 1586547711
transform 1 0 14200 0 1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL74520x68000
timestamp 1586547711
transform 1 0 15304 0 1 14000
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL78200x68000
timestamp 1586547711
transform 1 0 16040 0 1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1586547711
transform 1 0 16132 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_751
timestamp 1586547711
transform 1 0 16316 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_761
timestamp 1586547711
transform 1 0 16500 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_810
timestamp 1586547711
transform 1 0 16684 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_812
timestamp 1586547711
transform 1 0 16868 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_811
timestamp 1586547711
transform 1 0 17052 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_767
timestamp 1586547711
transform 1 0 17328 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1586547711
transform 1 0 17236 0 1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_727
timestamp 1586547711
transform 1 0 17512 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_730
timestamp 1586547711
transform 1 0 19352 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL92920x68000
timestamp 1586547711
transform 1 0 18984 0 1 14000
box 0 -48 368 592
use sky130_fd_sc_hd__a211o_4  _489_
timestamp 1586547711
transform 1 0 17696 0 1 14000
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA_296
timestamp 1586547711
transform 1 0 19536 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _466_
timestamp 1586547711
transform 1 0 19720 0 1 14000
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_8  FILL102580x68000
timestamp 1586547711
transform 1 0 20916 0 1 14000
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL106260x68000
timestamp 1586547711
transform 1 0 21652 0 1 14000
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_707
timestamp 1586547711
transform 1 0 21928 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_705
timestamp 1586547711
transform 1 0 22112 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_697
timestamp 1586547711
transform 1 0 22296 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_700
timestamp 1586547711
transform 1 0 22480 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_704
timestamp 1586547711
transform 1 0 22664 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1586547711
transform 1 0 22848 0 1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__o21a_4  _460_
timestamp 1586547711
transform 1 0 22940 0 1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL124660x68000
timestamp 1586547711
transform 1 0 25332 0 1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1052
timestamp 1586547711
transform 1 0 24044 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _525_
timestamp 1586547711
transform 1 0 25424 0 1 14000
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL119140x68000
timestamp 1586547711
transform 1 0 24228 0 1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1586547711
transform 1 0 26988 0 1 14000
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL132480x68000
timestamp 1586547711
transform 1 0 26896 0 1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_136
timestamp 1586547711
transform 1 0 25976 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_894
timestamp 1586547711
transform 1 0 26160 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL129720x68000
timestamp 1586547711
transform 1 0 26344 0 1 14000
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1586547711
transform 1 0 400 0 1 15088
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1586547711
transform 1 0 400 0 -1 15088
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1586547711
transform 1 0 1320 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL1380x73440
timestamp 1586547711
transform 1 0 676 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _283_
timestamp 1586547711
transform 1 0 860 0 1 15088
box 0 -48 460 592
use sky130_fd_sc_hd__fill_1  FILL6900x70720
timestamp 1586547711
transform 1 0 1780 0 -1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_288
timestamp 1586547711
transform 1 0 1504 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_485
timestamp 1586547711
transform 1 0 1688 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_481
timestamp 1586547711
transform 1 0 1872 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_500
timestamp 1586547711
transform 1 0 1872 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_490
timestamp 1586547711
transform 1 0 2056 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_587
timestamp 1586547711
transform 1 0 2240 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_603
timestamp 1586547711
transform 1 0 2424 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _405_
timestamp 1586547711
transform 1 0 2056 0 1 15088
box 0 -48 828 592
use sky130_fd_sc_hd__decap_12  FILL1380x70720
timestamp 1586547711
transform 1 0 676 0 -1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL13800x70720
timestamp 1586547711
transform 1 0 3160 0 -1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_457
timestamp 1586547711
transform 1 0 2884 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_612
timestamp 1586547711
transform 1 0 3068 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL11040x70720
timestamp 1586547711
transform 1 0 2608 0 -1 15088
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1586547711
transform 1 0 3252 0 -1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL14260x73440
timestamp 1586547711
transform 1 0 3252 0 1 15088
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL17940x73440
timestamp 1586547711
transform 1 0 3988 0 1 15088
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_542
timestamp 1586547711
transform 1 0 3988 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _390_
timestamp 1586547711
transform 1 0 3344 0 -1 15088
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_401
timestamp 1586547711
transform 1 0 4264 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_398
timestamp 1586547711
transform 1 0 4448 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_552
timestamp 1586547711
transform 1 0 4172 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _314_
timestamp 1586547711
transform 1 0 4632 0 1 15088
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL19780x70720
timestamp 1586547711
transform 1 0 4356 0 -1 15088
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_179
timestamp 1586547711
transform 1 0 5276 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_219
timestamp 1586547711
transform 1 0 5460 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _312_
timestamp 1586547711
transform 1 0 5092 0 -1 15088
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA_202
timestamp 1586547711
transform 1 0 5644 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_194
timestamp 1586547711
transform 1 0 5828 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_309
timestamp 1586547711
transform 1 0 5920 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_329
timestamp 1586547711
transform 1 0 6104 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_345
timestamp 1586547711
transform 1 0 6288 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1586547711
transform 1 0 6012 0 1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _300_
timestamp 1586547711
transform 1 0 6104 0 1 15088
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA_570
timestamp 1586547711
transform 1 0 6472 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1152
timestamp 1586547711
transform 1 0 6656 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL34040x70720
timestamp 1586547711
transform 1 0 7208 0 -1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_174
timestamp 1586547711
transform 1 0 6932 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_565
timestamp 1586547711
transform 1 0 7116 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_559
timestamp 1586547711
transform 1 0 7300 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_365
timestamp 1586547711
transform 1 0 7484 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL32200x70720
timestamp 1586547711
transform 1 0 6840 0 -1 15088
box 0 -48 368 592
use sky130_fd_sc_hd__or4_4  _377_
timestamp 1586547711
transform 1 0 7300 0 -1 15088
box 0 -48 828 592
use sky130_fd_sc_hd__or4_4  _378_
timestamp 1586547711
transform 1 0 7668 0 1 15088
box 0 -48 828 592
use sky130_fd_sc_hd__decap_8  FILL38640x70720
timestamp 1586547711
transform 1 0 8128 0 -1 15088
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_351
timestamp 1586547711
transform 1 0 8496 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1586547711
transform 1 0 8864 0 -1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL41400x73440
timestamp 1586547711
transform 1 0 8680 0 1 15088
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILL46000x70720
timestamp 1586547711
transform 1 0 9600 0 -1 15088
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL43240x73440
timestamp 1586547711
transform 1 0 9048 0 1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_176
timestamp 1586547711
transform 1 0 9140 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_195
timestamp 1586547711
transform 1 0 9324 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_307
timestamp 1586547711
transform 1 0 9508 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_358
timestamp 1586547711
transform 1 0 9692 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1105
timestamp 1586547711
transform 1 0 9876 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_353
timestamp 1586547711
transform 1 0 9876 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _299_
timestamp 1586547711
transform 1 0 8956 0 -1 15088
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1118
timestamp 1586547711
transform 1 0 10060 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL48300x73440
timestamp 1586547711
transform 1 0 10060 0 1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL49220x70720
timestamp 1586547711
transform 1 0 10244 0 -1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL53820x73440
timestamp 1586547711
transform 1 0 11164 0 1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_386
timestamp 1586547711
transform 1 0 11256 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_387
timestamp 1586547711
transform 1 0 11440 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL56580x73440
timestamp 1586547711
transform 1 0 11716 0 1 15088
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1586547711
transform 1 0 11624 0 1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__or4_4  _316_
timestamp 1586547711
transform 1 0 11348 0 -1 15088
box 0 -48 828 592
use sky130_fd_sc_hd__fill_1  FILL59340x73440
timestamp 1586547711
transform 1 0 12268 0 1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1267
timestamp 1586547711
transform 1 0 12360 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1262
timestamp 1586547711
transform 1 0 12544 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_999
timestamp 1586547711
transform 1 0 12728 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_998
timestamp 1586547711
transform 1 0 12912 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_410
timestamp 1586547711
transform 1 0 12176 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1145
timestamp 1586547711
transform 1 0 12360 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1260
timestamp 1586547711
transform 1 0 13096 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL60720x70720
timestamp 1586547711
transform 1 0 12544 0 -1 15088
box 0 -48 552 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[3\].id.delayenb0
timestamp 1586547711
transform 1 0 13096 0 1 15088
box 0 -48 1656 592
use sky130_fd_sc_hd__decap_3  FILL69000x70720
timestamp 1586547711
transform 1 0 14200 0 -1 15088
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_763
timestamp 1586547711
transform 1 0 15120 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1263
timestamp 1586547711
transform 1 0 13280 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1586547711
transform 1 0 14476 0 -1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL71760x73440
timestamp 1586547711
transform 1 0 14752 0 1 15088
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL70840x70720
timestamp 1586547711
transform 1 0 14568 0 -1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL65320x70720
timestamp 1586547711
transform 1 0 13464 0 -1 15088
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL78200x70720
timestamp 1586547711
transform 1 0 16040 0 -1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_760
timestamp 1586547711
transform 1 0 15304 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_756
timestamp 1586547711
transform 1 0 15488 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_755
timestamp 1586547711
transform 1 0 15672 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_757
timestamp 1586547711
transform 1 0 15856 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _471_
timestamp 1586547711
transform 1 0 15856 0 1 15088
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILL76360x70720
timestamp 1586547711
transform 1 0 15672 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_289
timestamp 1586547711
transform 1 0 16500 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_290
timestamp 1586547711
transform 1 0 16684 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_764
timestamp 1586547711
transform 1 0 16868 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1586547711
transform 1 0 17236 0 1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL84180x70720
timestamp 1586547711
transform 1 0 17236 0 -1 15088
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL83260x73440
timestamp 1586547711
transform 1 0 17052 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _488_
timestamp 1586547711
transform 1 0 16132 0 -1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL84640x73440
timestamp 1586547711
transform 1 0 17328 0 1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL86020x70720
timestamp 1586547711
transform 1 0 17604 0 -1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL87400x70720
timestamp 1586547711
transform 1 0 17880 0 -1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_768
timestamp 1586547711
transform 1 0 17696 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _475_
timestamp 1586547711
transform 1 0 17972 0 -1 15088
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL90160x73440
timestamp 1586547711
transform 1 0 18432 0 1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL90160x70720
timestamp 1586547711
transform 1 0 18432 0 -1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL98440x73440
timestamp 1586547711
transform 1 0 20088 0 1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1586547711
transform 1 0 20180 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_718
timestamp 1586547711
transform 1 0 20364 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_742
timestamp 1586547711
transform 1 0 19720 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL95680x73440
timestamp 1586547711
transform 1 0 19536 0 1 15088
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1586547711
transform 1 0 20088 0 -1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL95680x70720
timestamp 1586547711
transform 1 0 19536 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL97520x70720
timestamp 1586547711
transform 1 0 19904 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_724
timestamp 1586547711
transform 1 0 20548 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_725
timestamp 1586547711
transform 1 0 20732 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL104420x70720
timestamp 1586547711
transform 1 0 21284 0 -1 15088
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILL102580x73440
timestamp 1586547711
transform 1 0 20916 0 1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL98900x70720
timestamp 1586547711
transform 1 0 20180 0 -1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL108100x70720
timestamp 1586547711
transform 1 0 22020 0 -1 15088
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL109940x73440
timestamp 1586547711
transform 1 0 22388 0 1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_696
timestamp 1586547711
transform 1 0 22480 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL108100x73440
timestamp 1586547711
transform 1 0 22020 0 1 15088
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILL115000x73440
timestamp 1586547711
transform 1 0 23400 0 1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_649
timestamp 1586547711
transform 1 0 22664 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_112
timestamp 1586547711
transform 1 0 23492 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_242
timestamp 1586547711
transform 1 0 23676 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_268
timestamp 1586547711
transform 1 0 23584 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1586547711
transform 1 0 22848 0 1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _450_
timestamp 1586547711
transform 1 0 22940 0 1 15088
box 0 -48 460 592
use sky130_fd_sc_hd__o22a_4  _461_
timestamp 1586547711
transform 1 0 22296 0 -1 15088
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_1  FILL117300x73440
timestamp 1586547711
transform 1 0 23860 0 1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_113
timestamp 1586547711
transform 1 0 23952 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_640
timestamp 1586547711
transform 1 0 23768 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_895
timestamp 1586547711
transform 1 0 24136 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1025
timestamp 1586547711
transform 1 0 24320 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1078
timestamp 1586547711
transform 1 0 24504 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL117760x70720
timestamp 1586547711
transform 1 0 23952 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL121440x70720
timestamp 1586547711
transform 1 0 24688 0 -1 15088
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL125120x70720
timestamp 1586547711
transform 1 0 25424 0 -1 15088
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1586547711
transform 1 0 25700 0 -1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _548_
timestamp 1586547711
transform 1 0 24136 0 1 15088
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_12  FILL126960x70720
timestamp 1586547711
transform 1 0 25792 0 -1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1586547711
transform 1 0 26988 0 1 15088
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1586547711
transform 1 0 26988 0 -1 15088
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL132480x70720
timestamp 1586547711
transform 1 0 26896 0 -1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_267
timestamp 1586547711
transform 1 0 26252 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1076
timestamp 1586547711
transform 1 0 26436 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL131100x73440
timestamp 1586547711
transform 1 0 26620 0 1 15088
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1586547711
transform 1 0 400 0 -1 16176
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL5060x76160
timestamp 1586547711
transform 1 0 1412 0 -1 16176
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_613
timestamp 1586547711
transform 1 0 1688 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_596
timestamp 1586547711
transform 1 0 2516 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _357_
timestamp 1586547711
transform 1 0 1872 0 -1 16176
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL1380x76160
timestamp 1586547711
transform 1 0 676 0 -1 16176
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL17480x76160
timestamp 1586547711
transform 1 0 3896 0 -1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_571
timestamp 1586547711
transform 1 0 3988 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL11500x76160
timestamp 1586547711
transform 1 0 2700 0 -1 16176
box 0 -48 552 592
use sky130_fd_sc_hd__decap_6  FILL14720x76160
timestamp 1586547711
transform 1 0 3344 0 -1 16176
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1586547711
transform 1 0 3252 0 -1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL18860x76160
timestamp 1586547711
transform 1 0 4172 0 -1 16176
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1104
timestamp 1586547711
transform 1 0 6656 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL24380x76160
timestamp 1586547711
transform 1 0 5276 0 -1 16176
box 0 -48 552 592
use sky130_fd_sc_hd__and4_4  _381_
timestamp 1586547711
transform 1 0 5828 0 -1 16176
box 0 -48 828 592
use sky130_fd_sc_hd__fill_1  FILL35880x76160
timestamp 1586547711
transform 1 0 7576 0 -1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL39100x76160
timestamp 1586547711
transform 1 0 8220 0 -1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_564
timestamp 1586547711
transform 1 0 7668 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_311
timestamp 1586547711
transform 1 0 8312 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1586547711
transform 1 0 8864 0 -1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL37260x76160
timestamp 1586547711
transform 1 0 7852 0 -1 16176
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILL40480x76160
timestamp 1586547711
transform 1 0 8496 0 -1 16176
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILL32200x76160
timestamp 1586547711
transform 1 0 6840 0 -1 16176
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILL42780x76160
timestamp 1586547711
transform 1 0 8956 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _303_
timestamp 1586547711
transform 1 0 9140 0 -1 16176
box 0 -48 828 592
use sky130_fd_sc_hd__decap_12  FILL47840x76160
timestamp 1586547711
transform 1 0 9968 0 -1 16176
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL63020x76160
timestamp 1586547711
transform 1 0 13004 0 -1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_57
timestamp 1586547711
transform 1 0 11716 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_566
timestamp 1586547711
transform 1 0 11900 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_958
timestamp 1586547711
transform 1 0 12084 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen0
timestamp 1586547711
transform 1 0 13096 0 -1 16176
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILL53360x76160
timestamp 1586547711
transform 1 0 11072 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _310_
timestamp 1586547711
transform 1 0 11256 0 -1 16176
box 0 -48 460 592
use sky130_fd_sc_hd__decap_8  FILL59340x76160
timestamp 1586547711
transform 1 0 12268 0 -1 16176
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1586547711
transform 1 0 14476 0 -1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL66700x76160
timestamp 1586547711
transform 1 0 13740 0 -1 16176
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL70840x76160
timestamp 1586547711
transform 1 0 14568 0 -1 16176
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL75440x76160
timestamp 1586547711
transform 1 0 15488 0 -1 16176
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_759
timestamp 1586547711
transform 1 0 15304 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_750
timestamp 1586547711
transform 1 0 15764 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__a211o_4  _474_
timestamp 1586547711
transform 1 0 15948 0 -1 16176
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL84180x76160
timestamp 1586547711
transform 1 0 17236 0 -1 16176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILL95220x76160
timestamp 1586547711
transform 1 0 19444 0 -1 16176
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL89700x76160
timestamp 1586547711
transform 1 0 18340 0 -1 16176
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL97980x76160
timestamp 1586547711
transform 1 0 19996 0 -1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1586547711
transform 1 0 20088 0 -1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__o21a_4  _459_
timestamp 1586547711
transform 1 0 20180 0 -1 16176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL104420x76160
timestamp 1586547711
transform 1 0 21284 0 -1 16176
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_698
timestamp 1586547711
transform 1 0 22940 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL109940x76160
timestamp 1586547711
transform 1 0 22388 0 -1 16176
box 0 -48 552 592
use sky130_fd_sc_hd__decap_4  FILL113620x76160
timestamp 1586547711
transform 1 0 23124 0 -1 16176
box 0 -48 368 592
use sky130_fd_sc_hd__o22ai_4  _441_
timestamp 1586547711
transform 1 0 23492 0 -1 16176
box 0 -48 1472 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1057
timestamp 1586547711
transform 1 0 24964 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL123740x76160
timestamp 1586547711
transform 1 0 25148 0 -1 16176
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1586547711
transform 1 0 25700 0 -1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _277_
timestamp 1586547711
transform 1 0 25792 0 -1 16176
box 0 -48 460 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1586547711
transform 1 0 26988 0 -1 16176
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL129260x76160
timestamp 1586547711
transform 1 0 26252 0 -1 16176
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1586547711
transform 1 0 400 0 1 16176
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL3220x78880
timestamp 1586547711
transform 1 0 1044 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_614
timestamp 1586547711
transform 1 0 1136 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL1380x78880
timestamp 1586547711
transform 1 0 676 0 1 16176
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILL7360x78880
timestamp 1586547711
transform 1 0 1872 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_595
timestamp 1586547711
transform 1 0 1320 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_569
timestamp 1586547711
transform 1 0 1504 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_482
timestamp 1586547711
transform 1 0 1688 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_384
timestamp 1586547711
transform 1 0 1964 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_373
timestamp 1586547711
transform 1 0 2148 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _395_
timestamp 1586547711
transform 1 0 2332 0 1 16176
box 0 -48 828 592
use sky130_fd_sc_hd__fill_1  FILL14720x78880
timestamp 1586547711
transform 1 0 3344 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_344
timestamp 1586547711
transform 1 0 3160 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_572
timestamp 1586547711
transform 1 0 3436 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_489
timestamp 1586547711
transform 1 0 3620 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_456
timestamp 1586547711
transform 1 0 3804 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _382_
timestamp 1586547711
transform 1 0 3988 0 1 16176
box 0 -48 828 592
use sky130_fd_sc_hd__fill_1  FILL24840x78880
timestamp 1586547711
transform 1 0 5368 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_409
timestamp 1586547711
transform 1 0 4816 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_347
timestamp 1586547711
transform 1 0 5460 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_396
timestamp 1586547711
transform 1 0 5644 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_444
timestamp 1586547711
transform 1 0 5828 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1586547711
transform 1 0 6012 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL23000x78880
timestamp 1586547711
transform 1 0 5000 0 1 16176
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILL28520x78880
timestamp 1586547711
transform 1 0 6104 0 1 16176
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_395
timestamp 1586547711
transform 1 0 6840 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_402
timestamp 1586547711
transform 1 0 7024 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_405
timestamp 1586547711
transform 1 0 7208 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_208
timestamp 1586547711
transform 1 0 7944 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_191
timestamp 1586547711
transform 1 0 8128 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL34960x78880
timestamp 1586547711
transform 1 0 7392 0 1 16176
box 0 -48 552 592
use sky130_fd_sc_hd__and4_4  _291_
timestamp 1586547711
transform 1 0 8312 0 1 16176
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA_171
timestamp 1586547711
transform 1 0 9140 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1006
timestamp 1586547711
transform 1 0 10612 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_364
timestamp 1586547711
transform 1 0 10796 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_87
timestamp 1586547711
transform 1 0 10980 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL50140x78880
timestamp 1586547711
transform 1 0 10428 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL44620x78880
timestamp 1586547711
transform 1 0 9324 0 1 16176
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL55660x78880
timestamp 1586547711
transform 1 0 11532 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_78
timestamp 1586547711
transform 1 0 11164 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_48
timestamp 1586547711
transform 1 0 11348 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1586547711
transform 1 0 11624 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__a21bo_4  _379_
timestamp 1586547711
transform 1 0 11716 0 1 16176
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_12  FILL62560x78880
timestamp 1586547711
transform 1 0 12912 0 1 16176
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1259
timestamp 1586547711
transform 1 0 14568 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1261
timestamp 1586547711
transform 1 0 14752 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_749
timestamp 1586547711
transform 1 0 14936 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1586547711
transform 1 0 15120 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL68080x78880
timestamp 1586547711
transform 1 0 14016 0 1 16176
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1586547711
transform 1 0 16500 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_762
timestamp 1586547711
transform 1 0 16684 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_753
timestamp 1586547711
transform 1 0 17328 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1586547711
transform 1 0 17236 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL82340x78880
timestamp 1586547711
transform 1 0 16868 0 1 16176
box 0 -48 368 592
use sky130_fd_sc_hd__a21bo_4  _472_
timestamp 1586547711
transform 1 0 15304 0 1 16176
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA_710
timestamp 1586547711
transform 1 0 17512 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__xnor2_4  _470_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 17696 0 1 16176
box 0 -48 2024 592
use sky130_fd_sc_hd__decap_3  FILL96600x78880
timestamp 1586547711
transform 1 0 19720 0 1 16176
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_769
timestamp 1586547711
transform 1 0 19996 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_287
timestamp 1586547711
transform 1 0 20180 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_685
timestamp 1586547711
transform 1 0 20364 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_719
timestamp 1586547711
transform 1 0 20548 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_722
timestamp 1586547711
transform 1 0 20732 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1586547711
transform 1 0 21376 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_286
timestamp 1586547711
transform 1 0 21560 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _282_
timestamp 1586547711
transform 1 0 20916 0 1 16176
box 0 -48 460 592
use sky130_fd_sc_hd__diode_2  ANTENNA_703
timestamp 1586547711
transform 1 0 22296 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_270
timestamp 1586547711
transform 1 0 22480 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_244
timestamp 1586547711
transform 1 0 22664 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL106720x78880
timestamp 1586547711
transform 1 0 21744 0 1 16176
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1586547711
transform 1 0 22848 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _453_
timestamp 1586547711
transform 1 0 22940 0 1 16176
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1077
timestamp 1586547711
transform 1 0 24412 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_269
timestamp 1586547711
transform 1 0 24596 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_243
timestamp 1586547711
transform 1 0 24780 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL119140x78880
timestamp 1586547711
transform 1 0 24228 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _449_
timestamp 1586547711
transform 1 0 24964 0 1 16176
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1586547711
transform 1 0 26988 0 1 16176
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1586547711
transform 1 0 26252 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1023
timestamp 1586547711
transform 1 0 26436 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL131100x78880
timestamp 1586547711
transform 1 0 26620 0 1 16176
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1586547711
transform 1 0 400 0 -1 17264
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL5980x81600
timestamp 1586547711
transform 1 0 1596 0 -1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_71
timestamp 1586547711
transform 1 0 676 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_982
timestamp 1586547711
transform 1 0 860 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_594
timestamp 1586547711
transform 1 0 2516 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL3220x81600
timestamp 1586547711
transform 1 0 1044 0 -1 17264
box 0 -48 552 592
use sky130_fd_sc_hd__or4_4  _406_
timestamp 1586547711
transform 1 0 1688 0 -1 17264
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA_568
timestamp 1586547711
transform 1 0 4080 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_573
timestamp 1586547711
transform 1 0 4264 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_574
timestamp 1586547711
transform 1 0 4448 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL11500x81600
timestamp 1586547711
transform 1 0 2700 0 -1 17264
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1586547711
transform 1 0 3252 0 -1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL14720x81600
timestamp 1586547711
transform 1 0 3344 0 -1 17264
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL21160x81600
timestamp 1586547711
transform 1 0 4632 0 -1 17264
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL24840x81600
timestamp 1586547711
transform 1 0 5368 0 -1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_388
timestamp 1586547711
transform 1 0 6288 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL30360x81600
timestamp 1586547711
transform 1 0 6472 0 -1 17264
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _332_
timestamp 1586547711
transform 1 0 5460 0 -1 17264
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILL28520x81600
timestamp 1586547711
transform 1 0 6104 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL39100x81600
timestamp 1586547711
transform 1 0 8220 0 -1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_304
timestamp 1586547711
transform 1 0 8312 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1586547711
transform 1 0 8864 0 -1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL40480x81600
timestamp 1586547711
transform 1 0 8496 0 -1 17264
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _315_
timestamp 1586547711
transform 1 0 6840 0 -1 17264
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL35420x81600
timestamp 1586547711
transform 1 0 7484 0 -1 17264
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL42780x81600
timestamp 1586547711
transform 1 0 8956 0 -1 17264
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL45080x81600
timestamp 1586547711
transform 1 0 9416 0 -1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_441
timestamp 1586547711
transform 1 0 9232 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_361
timestamp 1586547711
transform 1 0 9508 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL51980x81600
timestamp 1586547711
transform 1 0 10796 0 -1 17264
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL46460x81600
timestamp 1586547711
transform 1 0 9692 0 -1 17264
box 0 -48 1104 592
use sky130_fd_sc_hd__a21bo_4  _336_
timestamp 1586547711
transform 1 0 11348 0 -1 17264
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_12  FILL60720x81600
timestamp 1586547711
transform 1 0 12544 0 -1 17264
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL69920x81600
timestamp 1586547711
transform 1 0 14384 0 -1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL74060x81600
timestamp 1586547711
transform 1 0 15212 0 -1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1586547711
transform 1 0 14476 0 -1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL72220x81600
timestamp 1586547711
transform 1 0 14844 0 -1 17264
box 0 -48 368 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[3\].id.delayint0
timestamp 1586547711
transform 1 0 14568 0 -1 17264
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL66240x81600
timestamp 1586547711
transform 1 0 13648 0 -1 17264
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL75440x81600
timestamp 1586547711
transform 1 0 15488 0 -1 17264
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_758
timestamp 1586547711
transform 1 0 15304 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _473_
timestamp 1586547711
transform 1 0 15764 0 -1 17264
box 0 -48 828 592
use sky130_fd_sc_hd__decap_12  FILL80960x81600
timestamp 1586547711
transform 1 0 16592 0 -1 17264
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_754
timestamp 1586547711
transform 1 0 17696 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL87400x81600
timestamp 1586547711
transform 1 0 17880 0 -1 17264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL92920x81600
timestamp 1586547711
transform 1 0 18984 0 -1 17264
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1586547711
transform 1 0 20088 0 -1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__a211o_4  _476_
timestamp 1586547711
transform 1 0 20180 0 -1 17264
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL105340x81600
timestamp 1586547711
transform 1 0 21468 0 -1 17264
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_699
timestamp 1586547711
transform 1 0 22940 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_708
timestamp 1586547711
transform 1 0 23124 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL110860x81600
timestamp 1586547711
transform 1 0 22572 0 -1 17264
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL114540x81600
timestamp 1586547711
transform 1 0 23308 0 -1 17264
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_695
timestamp 1586547711
transform 1 0 24964 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL120060x81600
timestamp 1586547711
transform 1 0 24412 0 -1 17264
box 0 -48 552 592
use sky130_fd_sc_hd__decap_6  FILL123740x81600
timestamp 1586547711
transform 1 0 25148 0 -1 17264
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1586547711
transform 1 0 25700 0 -1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__buf_2  _546_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 25792 0 -1 17264
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1586547711
transform 1 0 26988 0 -1 17264
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL132480x81600
timestamp 1586547711
transform 1 0 26896 0 -1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL128800x81600
timestamp 1586547711
transform 1 0 26160 0 -1 17264
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1586547711
transform 1 0 400 0 1 17264
box 0 -48 276 592
use sky130_fd_sc_hd__a21bo_4  _407_
timestamp 1586547711
transform 1 0 676 0 1 17264
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_8  FILL7360x84320
timestamp 1586547711
transform 1 0 1872 0 1 17264
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL11040x84320
timestamp 1586547711
transform 1 0 2608 0 1 17264
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_593
timestamp 1586547711
transform 1 0 2884 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_447
timestamp 1586547711
transform 1 0 3068 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_404
timestamp 1586547711
transform 1 0 3896 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_352
timestamp 1586547711
transform 1 0 4080 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_372
timestamp 1586547711
transform 1 0 4264 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_541
timestamp 1586547711
transform 1 0 4448 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _394_
timestamp 1586547711
transform 1 0 3252 0 1 17264
box 0 -48 644 592
use sky130_fd_sc_hd__or2_4  _369_
timestamp 1586547711
transform 1 0 4632 0 1 17264
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_393
timestamp 1586547711
transform 1 0 5276 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_446
timestamp 1586547711
transform 1 0 5460 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_390
timestamp 1586547711
transform 1 0 5644 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_348
timestamp 1586547711
transform 1 0 5828 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_341
timestamp 1586547711
transform 1 0 6748 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1586547711
transform 1 0 6012 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _301_
timestamp 1586547711
transform 1 0 6104 0 1 17264
box 0 -48 644 592
use sky130_fd_sc_hd__fill_1  FILL36340x84320
timestamp 1586547711
transform 1 0 7668 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_346
timestamp 1586547711
transform 1 0 6932 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_381
timestamp 1586547711
transform 1 0 7116 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_367
timestamp 1586547711
transform 1 0 7760 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_362
timestamp 1586547711
transform 1 0 7944 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_354
timestamp 1586547711
transform 1 0 8772 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL34500x84320
timestamp 1586547711
transform 1 0 7300 0 1 17264
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _305_
timestamp 1586547711
transform 1 0 8128 0 1 17264
box 0 -48 644 592
use sky130_fd_sc_hd__fill_1  FILL42780x84320
timestamp 1586547711
transform 1 0 8956 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL45080x84320
timestamp 1586547711
transform 1 0 9416 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_360
timestamp 1586547711
transform 1 0 9048 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_356
timestamp 1586547711
transform 1 0 9232 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _304_
timestamp 1586547711
transform 1 0 9508 0 1 17264
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_316
timestamp 1586547711
transform 1 0 10152 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_359
timestamp 1586547711
transform 1 0 10336 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp 1586547711
transform 1 0 10704 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL50600x84320
timestamp 1586547711
transform 1 0 10520 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_187
timestamp 1586547711
transform 1 0 10888 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILL62100x84320
timestamp 1586547711
transform 1 0 12820 0 1 17264
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_962
timestamp 1586547711
transform 1 0 13096 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL53360x84320
timestamp 1586547711
transform 1 0 11072 0 1 17264
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1586547711
transform 1 0 11624 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL56580x84320
timestamp 1586547711
transform 1 0 11716 0 1 17264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL66240x84320
timestamp 1586547711
transform 1 0 13648 0 1 17264
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1256
timestamp 1586547711
transform 1 0 13280 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1257
timestamp 1586547711
transform 1 0 13464 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1255
timestamp 1586547711
transform 1 0 14200 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1266
timestamp 1586547711
transform 1 0 14384 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1
timestamp 1586547711
transform 1 0 13924 0 1 17264
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL70840x84320
timestamp 1586547711
transform 1 0 14568 0 1 17264
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL82800x84320
timestamp 1586547711
transform 1 0 16960 0 1 17264
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_115
timestamp 1586547711
transform 1 0 15488 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_897
timestamp 1586547711
transform 1 0 15672 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1026
timestamp 1586547711
transform 1 0 15856 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1081
timestamp 1586547711
transform 1 0 16040 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1586547711
transform 1 0 17236 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL74520x84320
timestamp 1586547711
transform 1 0 15304 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL79120x84320
timestamp 1586547711
transform 1 0 16224 0 1 17264
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL84640x84320
timestamp 1586547711
transform 1 0 17328 0 1 17264
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL88320x84320
timestamp 1586547711
transform 1 0 18064 0 1 17264
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_271
timestamp 1586547711
transform 1 0 18340 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1079
timestamp 1586547711
transform 1 0 18524 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL91540x84320
timestamp 1586547711
transform 1 0 18708 0 1 17264
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL100740x84320
timestamp 1586547711
transform 1 0 20548 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_720
timestamp 1586547711
transform 1 0 19996 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_688
timestamp 1586547711
transform 1 0 20180 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_716
timestamp 1586547711
transform 1 0 20364 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_721
timestamp 1586547711
transform 1 0 21100 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_723
timestamp 1586547711
transform 1 0 21284 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL97060x84320
timestamp 1586547711
transform 1 0 19812 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _458_
timestamp 1586547711
transform 1 0 20640 0 1 17264
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL105340x84320
timestamp 1586547711
transform 1 0 21468 0 1 17264
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL110860x84320
timestamp 1586547711
transform 1 0 22572 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1048
timestamp 1586547711
transform 1 0 22664 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_102
timestamp 1586547711
transform 1 0 23400 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_245
timestamp 1586547711
transform 1 0 23584 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1586547711
transform 1 0 22848 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _272_
timestamp 1586547711
transform 1 0 22940 0 1 17264
box 0 -48 460 592
use sky130_fd_sc_hd__diode_2  ANTENNA_674
timestamp 1586547711
transform 1 0 23768 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_239
timestamp 1586547711
transform 1 0 24596 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1054
timestamp 1586547711
transform 1 0 24780 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL117760x84320
timestamp 1586547711
transform 1 0 23952 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _271_
timestamp 1586547711
transform 1 0 24136 0 1 17264
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL122820x84320
timestamp 1586547711
transform 1 0 24964 0 1 17264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1586547711
transform 1 0 26988 0 1 17264
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILL132020x84320
timestamp 1586547711
transform 1 0 26804 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL128340x84320
timestamp 1586547711
transform 1 0 26068 0 1 17264
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1586547711
transform 1 0 400 0 -1 18352
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_64
timestamp 1586547711
transform 1 0 676 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_615
timestamp 1586547711
transform 1 0 860 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_949
timestamp 1586547711
transform 1 0 1228 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL3220x87040
timestamp 1586547711
transform 1 0 1044 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL5060x87040
timestamp 1586547711
transform 1 0 1412 0 -1 18352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL10580x87040
timestamp 1586547711
transform 1 0 2516 0 -1 18352
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1586547711
transform 1 0 3252 0 -1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__or4_4  _383_
timestamp 1586547711
transform 1 0 4080 0 -1 18352
box 0 -48 828 592
use sky130_fd_sc_hd__decap_8  FILL14720x87040
timestamp 1586547711
transform 1 0 3344 0 -1 18352
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL28060x87040
timestamp 1586547711
transform 1 0 6012 0 -1 18352
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_453
timestamp 1586547711
transform 1 0 4908 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_483
timestamp 1586547711
transform 1 0 5092 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _311_
timestamp 1586547711
transform 1 0 6288 0 -1 18352
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL24380x87040
timestamp 1586547711
transform 1 0 5276 0 -1 18352
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL34500x87040
timestamp 1586547711
transform 1 0 7300 0 -1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_342
timestamp 1586547711
transform 1 0 7392 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_416
timestamp 1586547711
transform 1 0 7576 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_448
timestamp 1586547711
transform 1 0 7760 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1586547711
transform 1 0 8864 0 -1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL32660x87040
timestamp 1586547711
transform 1 0 6932 0 -1 18352
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL41400x87040
timestamp 1586547711
transform 1 0 8680 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL37720x87040
timestamp 1586547711
transform 1 0 7944 0 -1 18352
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL42780x87040
timestamp 1586547711
transform 1 0 8956 0 -1 18352
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL51060x87040
timestamp 1586547711
transform 1 0 10612 0 -1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_985
timestamp 1586547711
transform 1 0 10060 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL49220x87040
timestamp 1586547711
transform 1 0 10244 0 -1 18352
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _331_
timestamp 1586547711
transform 1 0 9232 0 -1 18352
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILL47380x87040
timestamp 1586547711
transform 1 0 9876 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _262_
timestamp 1586547711
transform 1 0 10704 0 -1 18352
box 0 -48 460 592
use sky130_fd_sc_hd__fill_1  FILL63020x87040
timestamp 1586547711
transform 1 0 13004 0 -1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen1
timestamp 1586547711
transform 1 0 13096 0 -1 18352
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL53820x87040
timestamp 1586547711
transform 1 0 11164 0 -1 18352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL59340x87040
timestamp 1586547711
transform 1 0 12268 0 -1 18352
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1268
timestamp 1586547711
transform 1 0 13740 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL67620x87040
timestamp 1586547711
transform 1 0 13924 0 -1 18352
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1586547711
transform 1 0 14476 0 -1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL70840x87040
timestamp 1586547711
transform 1 0 14568 0 -1 18352
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILL74520x87040
timestamp 1586547711
transform 1 0 15304 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _549_
timestamp 1586547711
transform 1 0 15488 0 -1 18352
box 0 -48 2116 592
use sky130_fd_sc_hd__fill_1  FILL86020x87040
timestamp 1586547711
transform 1 0 17604 0 -1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL89240x87040
timestamp 1586547711
transform 1 0 18248 0 -1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_259
timestamp 1586547711
transform 1 0 17696 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_274
timestamp 1586547711
transform 1 0 17880 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_693
timestamp 1586547711
transform 1 0 18064 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _278_
timestamp 1586547711
transform 1 0 18340 0 -1 18352
box 0 -48 460 592
use sky130_fd_sc_hd__decap_8  FILL92000x87040
timestamp 1586547711
transform 1 0 18800 0 -1 18352
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1080
timestamp 1586547711
transform 1 0 19536 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1586547711
transform 1 0 20088 0 -1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL96600x87040
timestamp 1586547711
transform 1 0 19720 0 -1 18352
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _457_
timestamp 1586547711
transform 1 0 20180 0 -1 18352
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL102120x87040
timestamp 1586547711
transform 1 0 20824 0 -1 18352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL111320x87040
timestamp 1586547711
transform 1 0 22664 0 -1 18352
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL113620x87040
timestamp 1586547711
transform 1 0 23124 0 -1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_672
timestamp 1586547711
transform 1 0 22940 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_667
timestamp 1586547711
transform 1 0 23216 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _432_
timestamp 1586547711
transform 1 0 23400 0 -1 18352
box 0 -48 460 592
use sky130_fd_sc_hd__decap_8  FILL107640x87040
timestamp 1586547711
transform 1 0 21928 0 -1 18352
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1056
timestamp 1586547711
transform 1 0 23860 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL123740x87040
timestamp 1586547711
transform 1 0 25148 0 -1 18352
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1586547711
transform 1 0 25700 0 -1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL118220x87040
timestamp 1586547711
transform 1 0 24044 0 -1 18352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL126960x87040
timestamp 1586547711
transform 1 0 25792 0 -1 18352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1586547711
transform 1 0 26988 0 -1 18352
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL132480x87040
timestamp 1586547711
transform 1 0 26896 0 -1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1586547711
transform 1 0 400 0 -1 19440
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1586547711
transform 1 0 400 0 1 18352
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_376
timestamp 1586547711
transform 1 0 1228 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_81
timestamp 1586547711
transform 1 0 860 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_54
timestamp 1586547711
transform 1 0 1044 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL1380x92480
timestamp 1586547711
transform 1 0 676 0 -1 19440
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILL1380x89760
timestamp 1586547711
transform 1 0 676 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL10120x89760
timestamp 1586547711
transform 1 0 2424 0 1 18352
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL10580x92480
timestamp 1586547711
transform 1 0 2516 0 -1 19440
box 0 -48 736 592
use sky130_fd_sc_hd__a21bo_4  _350_
timestamp 1586547711
transform 1 0 1228 0 1 18352
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_12  FILL5060x92480
timestamp 1586547711
transform 1 0 1412 0 -1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_479
timestamp 1586547711
transform 1 0 2976 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1586547711
transform 1 0 3252 0 -1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _345_
timestamp 1586547711
transform 1 0 3160 0 1 18352
box 0 -48 644 592
use sky130_fd_sc_hd__fill_1  FILL18860x89760
timestamp 1586547711
transform 1 0 4172 0 1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_343
timestamp 1586547711
transform 1 0 3804 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_370
timestamp 1586547711
transform 1 0 3988 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_424
timestamp 1586547711
transform 1 0 4264 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_423
timestamp 1586547711
transform 1 0 4448 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _351_
timestamp 1586547711
transform 1 0 4632 0 -1 19440
box 0 -48 644 592
use sky130_fd_sc_hd__or2_4  _337_
timestamp 1586547711
transform 1 0 4632 0 1 18352
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILL20240x92480
timestamp 1586547711
transform 1 0 4448 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL14720x92480
timestamp 1586547711
transform 1 0 3344 0 -1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_389
timestamp 1586547711
transform 1 0 5276 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_403
timestamp 1586547711
transform 1 0 5460 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_445
timestamp 1586547711
transform 1 0 6656 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL29900x92480
timestamp 1586547711
transform 1 0 6380 0 -1 19440
box 0 -48 552 592
use sky130_fd_sc_hd__decap_6  FILL28520x89760
timestamp 1586547711
transform 1 0 6104 0 1 18352
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1586547711
transform 1 0 6012 0 1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL26220x89760
timestamp 1586547711
transform 1 0 5644 0 1 18352
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL24380x92480
timestamp 1586547711
transform 1 0 5276 0 -1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL34040x92480
timestamp 1586547711
transform 1 0 7208 0 -1 19440
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL32660x92480
timestamp 1586547711
transform 1 0 6932 0 -1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_436
timestamp 1586547711
transform 1 0 7024 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_418
timestamp 1586547711
transform 1 0 6840 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_313
timestamp 1586547711
transform 1 0 7024 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_180
timestamp 1586547711
transform 1 0 7208 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _319_
timestamp 1586547711
transform 1 0 7484 0 -1 19440
box 0 -48 644 592
use sky130_fd_sc_hd__or4_4  _333_
timestamp 1586547711
transform 1 0 7392 0 1 18352
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA_46
timestamp 1586547711
transform 1 0 8220 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL40020x89760
timestamp 1586547711
transform 1 0 8404 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL38640x92480
timestamp 1586547711
transform 1 0 8128 0 -1 19440
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_314
timestamp 1586547711
transform 1 0 8588 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_312
timestamp 1586547711
transform 1 0 8772 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1586547711
transform 1 0 8864 0 -1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL46920x89760
timestamp 1586547711
transform 1 0 9784 0 1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_40
timestamp 1586547711
transform 1 0 9600 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_223
timestamp 1586547711
transform 1 0 9876 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _292_
timestamp 1586547711
transform 1 0 8956 0 1 18352
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_65
timestamp 1586547711
transform 1 0 10060 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_186
timestamp 1586547711
transform 1 0 10244 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_188
timestamp 1586547711
transform 1 0 10888 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _317_
timestamp 1586547711
transform 1 0 10428 0 1 18352
box 0 -48 460 592
use sky130_fd_sc_hd__o22ai_4  _408_
timestamp 1586547711
transform 1 0 10060 0 -1 19440
box 0 -48 1472 592
use sky130_fd_sc_hd__decap_12  FILL42780x92480
timestamp 1586547711
transform 1 0 8956 0 -1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_411
timestamp 1586547711
transform 1 0 11072 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_412
timestamp 1586547711
transform 1 0 11256 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL56580x89760
timestamp 1586547711
transform 1 0 11716 0 1 18352
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1586547711
transform 1 0 11624 0 1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL55200x89760
timestamp 1586547711
transform 1 0 11440 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL55660x92480
timestamp 1586547711
transform 1 0 11532 0 -1 19440
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL59340x92480
timestamp 1586547711
transform 1 0 12268 0 -1 19440
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL59340x89760
timestamp 1586547711
transform 1 0 12268 0 1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL63480x89760
timestamp 1586547711
transform 1 0 13096 0 1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_961
timestamp 1586547711
transform 1 0 12360 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_58
timestamp 1586547711
transform 1 0 12544 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_77
timestamp 1586547711
transform 1 0 12728 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_575
timestamp 1586547711
transform 1 0 12912 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _384_
timestamp 1586547711
transform 1 0 12544 0 -1 19440
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1258
timestamp 1586547711
transform 1 0 13740 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_963
timestamp 1586547711
transform 1 0 14200 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL67620x92480
timestamp 1586547711
transform 1 0 13924 0 -1 19440
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1586547711
transform 1 0 14476 0 -1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[3\].id.delayenb1
timestamp 1586547711
transform 1 0 13188 0 1 18352
box 0 -48 1012 592
use sky130_fd_sc_hd__decap_12  FILL70840x92480
timestamp 1586547711
transform 1 0 14568 0 -1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL69920x89760
timestamp 1586547711
transform 1 0 14384 0 1 18352
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL75440x89760
timestamp 1586547711
transform 1 0 15488 0 1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_137
timestamp 1586547711
transform 1 0 16132 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _526_
timestamp 1586547711
transform 1 0 15580 0 1 18352
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_272
timestamp 1586547711
transform 1 0 17328 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_896
timestamp 1586547711
transform 1 0 16316 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_641
timestamp 1586547711
transform 1 0 16684 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_257
timestamp 1586547711
transform 1 0 16868 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_114
timestamp 1586547711
transform 1 0 17052 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL81880x92480
timestamp 1586547711
transform 1 0 16776 0 -1 19440
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1586547711
transform 1 0 17236 0 1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL80500x89760
timestamp 1586547711
transform 1 0 16500 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__o22ai_4  _442_
timestamp 1586547711
transform 1 0 17328 0 1 18352
box 0 -48 1472 592
use sky130_fd_sc_hd__decap_12  FILL76360x92480
timestamp 1586547711
transform 1 0 15672 0 -1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_650
timestamp 1586547711
transform 1 0 17512 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_709
timestamp 1586547711
transform 1 0 18800 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_711
timestamp 1586547711
transform 1 0 18984 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_752
timestamp 1586547711
transform 1 0 19168 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_694
timestamp 1586547711
transform 1 0 19352 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL92920x92480
timestamp 1586547711
transform 1 0 18984 0 -1 19440
box 0 -48 552 592
use sky130_fd_sc_hd__o22a_4  _454_
timestamp 1586547711
transform 1 0 17696 0 -1 19440
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1061
timestamp 1586547711
transform 1 0 19536 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1059
timestamp 1586547711
transform 1 0 20180 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1586547711
transform 1 0 20088 0 -1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL96600x92480
timestamp 1586547711
transform 1 0 19720 0 -1 19440
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILL99820x92480
timestamp 1586547711
transform 1 0 20364 0 -1 19440
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL103500x92480
timestamp 1586547711
transform 1 0 21100 0 -1 19440
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL104420x89760
timestamp 1586547711
transform 1 0 21284 0 1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_241
timestamp 1586547711
transform 1 0 21376 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_248
timestamp 1586547711
transform 1 0 21560 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL101660x89760
timestamp 1586547711
transform 1 0 20732 0 1 18352
box 0 -48 552 592
use sky130_fd_sc_hd__o21a_4  _433_
timestamp 1586547711
transform 1 0 21376 0 -1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__a21oi_4  _469_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 19536 0 1 18352
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA_256
timestamp 1586547711
transform 1 0 21744 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_675
timestamp 1586547711
transform 1 0 21928 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_673
timestamp 1586547711
transform 1 0 22112 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_671
timestamp 1586547711
transform 1 0 22296 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_247
timestamp 1586547711
transform 1 0 22480 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL110400x92480
timestamp 1586547711
transform 1 0 22480 0 -1 19440
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILL112240x92480
timestamp 1586547711
transform 1 0 22848 0 -1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL113620x92480
timestamp 1586547711
transform 1 0 23124 0 -1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_636
timestamp 1586547711
transform 1 0 22940 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_240
timestamp 1586547711
transform 1 0 22664 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1586547711
transform 1 0 22848 0 1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__and3_4  _430_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 23216 0 -1 19440
box 0 -48 828 592
use sky130_fd_sc_hd__a211o_4  _431_
timestamp 1586547711
transform 1 0 22940 0 1 18352
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1051
timestamp 1586547711
transform 1 0 24228 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL120060x89760
timestamp 1586547711
transform 1 0 24412 0 1 18352
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILL126500x89760
timestamp 1586547711
transform 1 0 25700 0 1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_918
timestamp 1586547711
transform 1 0 24964 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_70
timestamp 1586547711
transform 1 0 25792 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL123740x92480
timestamp 1586547711
transform 1 0 25148 0 -1 19440
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1586547711
transform 1 0 25700 0 -1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _265_
timestamp 1586547711
transform 1 0 25792 0 -1 19440
box 0 -48 460 592
use sky130_fd_sc_hd__buf_4  _537_
timestamp 1586547711
transform 1 0 25148 0 1 18352
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL118220x92480
timestamp 1586547711
transform 1 0 24044 0 -1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1586547711
transform 1 0 26988 0 -1 19440
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1586547711
transform 1 0 26988 0 1 18352
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL132480x89760
timestamp 1586547711
transform 1 0 26896 0 1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_148
timestamp 1586547711
transform 1 0 25976 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_222
timestamp 1586547711
transform 1 0 26160 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL129720x89760
timestamp 1586547711
transform 1 0 26344 0 1 18352
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL129260x92480
timestamp 1586547711
transform 1 0 26252 0 -1 19440
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1586547711
transform 1 0 400 0 1 19440
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL5060x95200
timestamp 1586547711
transform 1 0 1412 0 1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_50
timestamp 1586547711
transform 1 0 676 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_85
timestamp 1586547711
transform 1 0 860 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_480
timestamp 1586547711
transform 1 0 1044 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1012
timestamp 1586547711
transform 1 0 1228 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1321
timestamp 1586547711
transform 1 0 1872 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1336
timestamp 1586547711
transform 1 0 2056 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[8\].id.delaybuf0
timestamp 1586547711
transform 1 0 1504 0 1 19440
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL9200x95200
timestamp 1586547711
transform 1 0 2240 0 1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_349
timestamp 1586547711
transform 1 0 4080 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_368
timestamp 1586547711
transform 1 0 4264 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_374
timestamp 1586547711
transform 1 0 4448 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL14720x95200
timestamp 1586547711
transform 1 0 3344 0 1 19440
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL21160x95200
timestamp 1586547711
transform 1 0 4632 0 1 19440
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL24840x95200
timestamp 1586547711
transform 1 0 5368 0 1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_375
timestamp 1586547711
transform 1 0 5460 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_391
timestamp 1586547711
transform 1 0 5644 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_406
timestamp 1586547711
transform 1 0 5828 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_422
timestamp 1586547711
transform 1 0 6104 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_425
timestamp 1586547711
transform 1 0 6288 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_484
timestamp 1586547711
transform 1 0 6472 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_420
timestamp 1586547711
transform 1 0 6656 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1586547711
transform 1 0 6012 0 1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_407
timestamp 1586547711
transform 1 0 6840 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_350
timestamp 1586547711
transform 1 0 7024 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_369
timestamp 1586547711
transform 1 0 7208 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_450
timestamp 1586547711
transform 1 0 8220 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_497
timestamp 1586547711
transform 1 0 8404 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_496
timestamp 1586547711
transform 1 0 8588 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_443
timestamp 1586547711
transform 1 0 8772 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _355_
timestamp 1586547711
transform 1 0 7392 0 1 19440
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA_392
timestamp 1586547711
transform 1 0 9600 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_442
timestamp 1586547711
transform 1 0 9784 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_449
timestamp 1586547711
transform 1 0 9968 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_451
timestamp 1586547711
transform 1 0 10152 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _354_
timestamp 1586547711
transform 1 0 8956 0 1 19440
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL49680x95200
timestamp 1586547711
transform 1 0 10336 0 1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILL62100x95200
timestamp 1586547711
transform 1 0 12820 0 1 19440
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1586547711
transform 1 0 11624 0 1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL55200x95200
timestamp 1586547711
transform 1 0 11440 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL56580x95200
timestamp 1586547711
transform 1 0 11716 0 1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1250
timestamp 1586547711
transform 1 0 13372 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1265
timestamp 1586547711
transform 1 0 13556 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL72220x95200
timestamp 1586547711
transform 1 0 14844 0 1 19440
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL66700x95200
timestamp 1586547711
transform 1 0 13740 0 1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_713
timestamp 1586547711
transform 1 0 15396 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_747
timestamp 1586547711
transform 1 0 15580 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_748
timestamp 1586547711
transform 1 0 15764 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1586547711
transform 1 0 17236 0 1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL83260x95200
timestamp 1586547711
transform 1 0 17052 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL77740x95200
timestamp 1586547711
transform 1 0 15948 0 1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL84640x95200
timestamp 1586547711
transform 1 0 17328 0 1 19440
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL88320x95200
timestamp 1586547711
transform 1 0 18064 0 1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_692
timestamp 1586547711
transform 1 0 18156 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_258
timestamp 1586547711
transform 1 0 18984 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_273
timestamp 1586547711
transform 1 0 19168 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL94760x95200
timestamp 1586547711
transform 1 0 19352 0 1 19440
box 0 -48 368 592
use sky130_fd_sc_hd__and2_4  _448_
timestamp 1586547711
transform 1 0 18340 0 1 19440
box 0 -48 644 592
use sky130_fd_sc_hd__fill_1  FILL96600x95200
timestamp 1586547711
transform 1 0 19720 0 1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_717
timestamp 1586547711
transform 1 0 19812 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_715
timestamp 1586547711
transform 1 0 19996 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_255
timestamp 1586547711
transform 1 0 20824 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_687
timestamp 1586547711
transform 1 0 21008 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_654
timestamp 1586547711
transform 1 0 21560 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL103960x95200
timestamp 1586547711
transform 1 0 21192 0 1 19440
box 0 -48 368 592
use sky130_fd_sc_hd__and2_4  _456_
timestamp 1586547711
transform 1 0 20180 0 1 19440
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  FILL112700x95200
timestamp 1586547711
transform 1 0 22940 0 1 19440
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1049
timestamp 1586547711
transform 1 0 21744 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1055
timestamp 1586547711
transform 1 0 21928 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1060
timestamp 1586547711
transform 1 0 22112 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1058
timestamp 1586547711
transform 1 0 23216 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_919
timestamp 1586547711
transform 1 0 23400 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_103
timestamp 1586547711
transform 1 0 23584 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL109480x95200
timestamp 1586547711
transform 1 0 22296 0 1 19440
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1586547711
transform 1 0 22848 0 1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _560_
timestamp 1586547711
transform 1 0 23768 0 1 19440
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1586547711
transform 1 0 26988 0 1 19440
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL127420x95200
timestamp 1586547711
transform 1 0 25884 0 1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1586547711
transform 1 0 400 0 -1 20528
box 0 -48 276 592
use sky130_fd_sc_hd__a21bo_4  _346_
timestamp 1586547711
transform 1 0 676 0 -1 20528
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_12  FILL7360x97920
timestamp 1586547711
transform 1 0 1872 0 -1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL12880x97920
timestamp 1586547711
transform 1 0 2976 0 -1 20528
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1586547711
transform 1 0 3252 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _306_
timestamp 1586547711
transform 1 0 4080 0 -1 20528
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL14720x97920
timestamp 1586547711
transform 1 0 3344 0 -1 20528
box 0 -48 736 592
use sky130_fd_sc_hd__or4_4  _321_
timestamp 1586547711
transform 1 0 5460 0 -1 20528
box 0 -48 828 592
use sky130_fd_sc_hd__decap_8  FILL21620x97920
timestamp 1586547711
transform 1 0 4724 0 -1 20528
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL29440x97920
timestamp 1586547711
transform 1 0 6288 0 -1 20528
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL41860x97920
timestamp 1586547711
transform 1 0 8772 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_492
timestamp 1586547711
transform 1 0 7852 0 -1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_498
timestamp 1586547711
transform 1 0 8036 0 -1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL39100x97920
timestamp 1586547711
transform 1 0 8220 0 -1 20528
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1586547711
transform 1 0 8864 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__or4_4  _328_
timestamp 1586547711
transform 1 0 7024 0 -1 20528
box 0 -48 828 592
use sky130_fd_sc_hd__fill_1  FILL44620x97920
timestamp 1586547711
transform 1 0 9324 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL42780x97920
timestamp 1586547711
transform 1 0 8956 0 -1 20528
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _334_
timestamp 1586547711
transform 1 0 9416 0 -1 20528
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL48300x97920
timestamp 1586547711
transform 1 0 10060 0 -1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL53820x97920
timestamp 1586547711
transform 1 0 11164 0 -1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL59340x97920
timestamp 1586547711
transform 1 0 12268 0 -1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1586547711
transform 1 0 14476 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[3\].id.delaybuf0
timestamp 1586547711
transform 1 0 13372 0 -1 20528
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILL66700x97920
timestamp 1586547711
transform 1 0 13740 0 -1 20528
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL70840x97920
timestamp 1586547711
transform 1 0 14568 0 -1 20528
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL74520x97920
timestamp 1586547711
transform 1 0 15304 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__xor2_4  _468_ /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 15396 0 -1 20528
box 0 -48 2024 592
use sky130_fd_sc_hd__decap_12  FILL85100x97920
timestamp 1586547711
transform 1 0 17420 0 -1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL90620x97920
timestamp 1586547711
transform 1 0 18524 0 -1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL97980x97920
timestamp 1586547711
transform 1 0 19996 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1586547711
transform 1 0 20088 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL96140x97920
timestamp 1586547711
transform 1 0 19628 0 -1 20528
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL104880x97920
timestamp 1586547711
transform 1 0 21376 0 -1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _274_
timestamp 1586547711
transform 1 0 20180 0 -1 20528
box 0 -48 460 592
use sky130_fd_sc_hd__and3_4  _424_
timestamp 1586547711
transform 1 0 21560 0 -1 20528
box 0 -48 828 592
use sky130_fd_sc_hd__decap_8  FILL101200x97920
timestamp 1586547711
transform 1 0 20640 0 -1 20528
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL115460x97920
timestamp 1586547711
transform 1 0 23492 0 -1 20528
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL109940x97920
timestamp 1586547711
transform 1 0 22388 0 -1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL126040x97920
timestamp 1586547711
transform 1 0 25608 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1037
timestamp 1586547711
transform 1 0 23768 0 -1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL123280x97920
timestamp 1586547711
transform 1 0 25056 0 -1 20528
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1586547711
transform 1 0 25700 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL117760x97920
timestamp 1586547711
transform 1 0 23952 0 -1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL126960x97920
timestamp 1586547711
transform 1 0 25792 0 -1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1586547711
transform 1 0 26988 0 -1 20528
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL132480x97920
timestamp 1586547711
transform 1 0 26896 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1586547711
transform 1 0 400 0 1 20528
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL6900x100640
timestamp 1586547711
transform 1 0 1780 0 1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1330
timestamp 1586547711
transform 1 0 1872 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1332
timestamp 1586547711
transform 1 0 2056 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL1380x100640
timestamp 1586547711
transform 1 0 676 0 1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL9200x100640
timestamp 1586547711
transform 1 0 2240 0 1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL20240x100640
timestamp 1586547711
transform 1 0 4448 0 1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_986
timestamp 1586547711
transform 1 0 4540 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL14720x100640
timestamp 1586547711
transform 1 0 3344 0 1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1195
timestamp 1586547711
transform 1 0 4724 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1196
timestamp 1586547711
transform 1 0 4908 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1586547711
transform 1 0 6012 0 1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL27140x100640
timestamp 1586547711
transform 1 0 5828 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL28520x100640
timestamp 1586547711
transform 1 0 6104 0 1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL23460x100640
timestamp 1586547711
transform 1 0 5092 0 1 20528
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_421
timestamp 1586547711
transform 1 0 7208 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_413
timestamp 1586547711
transform 1 0 8036 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_419
timestamp 1586547711
transform 1 0 8220 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _320_
timestamp 1586547711
transform 1 0 7392 0 1 20528
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL40020x100640
timestamp 1586547711
transform 1 0 8404 0 1 20528
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL43700x100640
timestamp 1586547711
transform 1 0 9140 0 1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_414
timestamp 1586547711
transform 1 0 9232 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_437
timestamp 1586547711
transform 1 0 9416 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_439
timestamp 1586547711
transform 1 0 9600 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL46920x100640
timestamp 1586547711
transform 1 0 9784 0 1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL52440x100640
timestamp 1586547711
transform 1 0 10888 0 1 20528
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL56580x100640
timestamp 1586547711
transform 1 0 11716 0 1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_45
timestamp 1586547711
transform 1 0 11808 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_89
timestamp 1586547711
transform 1 0 11992 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_440
timestamp 1586547711
transform 1 0 12176 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1000
timestamp 1586547711
transform 1 0 12360 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1003
timestamp 1586547711
transform 1 0 12912 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_88
timestamp 1586547711
transform 1 0 13096 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1586547711
transform 1 0 11624 0 1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL60720x100640
timestamp 1586547711
transform 1 0 12544 0 1 20528
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_47
timestamp 1586547711
transform 1 0 13280 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _335_
timestamp 1586547711
transform 1 0 13464 0 1 20528
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_12  FILL71300x100640
timestamp 1586547711
transform 1 0 14660 0 1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL78660x100640
timestamp 1586547711
transform 1 0 16132 0 1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_254
timestamp 1586547711
transform 1 0 16224 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL76820x100640
timestamp 1586547711
transform 1 0 15764 0 1 20528
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILL83720x100640
timestamp 1586547711
transform 1 0 17144 0 1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_278
timestamp 1586547711
transform 1 0 16408 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_690
timestamp 1586547711
transform 1 0 16592 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_712
timestamp 1586547711
transform 1 0 16776 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_714
timestamp 1586547711
transform 1 0 16960 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1586547711
transform 1 0 17236 0 1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL84640x100640
timestamp 1586547711
transform 1 0 17328 0 1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL90160x100640
timestamp 1586547711
transform 1 0 18432 0 1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL95680x100640
timestamp 1586547711
transform 1 0 19536 0 1 20528
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_104
timestamp 1586547711
transform 1 0 20272 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_678
timestamp 1586547711
transform 1 0 20456 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _435_
timestamp 1586547711
transform 1 0 19812 0 1 20528
box 0 -48 460 592
use sky130_fd_sc_hd__diode_2  ANTENNA_637
timestamp 1586547711
transform 1 0 20640 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_656
timestamp 1586547711
transform 1 0 20824 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_668
timestamp 1586547711
transform 1 0 21008 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_676
timestamp 1586547711
transform 1 0 21192 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_677
timestamp 1586547711
transform 1 0 21376 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL105800x100640
timestamp 1586547711
transform 1 0 21560 0 1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_100
timestamp 1586547711
transform 1 0 22664 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_246
timestamp 1586547711
transform 1 0 22940 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_635
timestamp 1586547711
transform 1 0 23124 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_666
timestamp 1586547711
transform 1 0 23308 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_670
timestamp 1586547711
transform 1 0 23492 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1586547711
transform 1 0 22848 0 1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL116380x100640
timestamp 1586547711
transform 1 0 23676 0 1 20528
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_147
timestamp 1586547711
transform 1 0 25148 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_916
timestamp 1586547711
transform 1 0 25332 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL120060x100640
timestamp 1586547711
transform 1 0 24412 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _536_
timestamp 1586547711
transform 1 0 24596 0 1 20528
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL125580x100640
timestamp 1586547711
transform 1 0 25516 0 1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1586547711
transform 1 0 26988 0 1 20528
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILL131100x100640
timestamp 1586547711
transform 1 0 26620 0 1 20528
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1586547711
transform 1 0 400 0 -1 21616
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL1380x103360
timestamp 1586547711
transform 1 0 676 0 -1 21616
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL3680x103360
timestamp 1586547711
transform 1 0 1136 0 -1 21616
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL6900x103360
timestamp 1586547711
transform 1 0 1780 0 -1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1338
timestamp 1586547711
transform 1 0 952 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1013
timestamp 1586547711
transform 1 0 1412 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1331
timestamp 1586547711
transform 1 0 1596 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[8\].id.delayint0
timestamp 1586547711
transform 1 0 1872 0 -1 21616
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL8740x103360
timestamp 1586547711
transform 1 0 2148 0 -1 21616
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL20240x103360
timestamp 1586547711
transform 1 0 4448 0 -1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1210
timestamp 1586547711
transform 1 0 4264 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen1
timestamp 1586547711
transform 1 0 4540 0 -1 21616
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1586547711
transform 1 0 3252 0 -1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL18400x103360
timestamp 1586547711
transform 1 0 4080 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL14720x103360
timestamp 1586547711
transform 1 0 3344 0 -1 21616
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILL23920x103360
timestamp 1586547711
transform 1 0 5184 0 -1 21616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL29440x103360
timestamp 1586547711
transform 1 0 6288 0 -1 21616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL34960x103360
timestamp 1586547711
transform 1 0 7392 0 -1 21616
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL40940x103360
timestamp 1586547711
transform 1 0 8588 0 -1 21616
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_973
timestamp 1586547711
transform 1 0 7668 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1586547711
transform 1 0 8864 0 -1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL37260x103360
timestamp 1586547711
transform 1 0 7852 0 -1 21616
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL42780x103360
timestamp 1586547711
transform 1 0 8956 0 -1 21616
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1252
timestamp 1586547711
transform 1 0 10796 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _329_
timestamp 1586547711
transform 1 0 9232 0 -1 21616
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILL51060x103360
timestamp 1586547711
transform 1 0 10612 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL47380x103360
timestamp 1586547711
transform 1 0 9876 0 -1 21616
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL52900x103360
timestamp 1586547711
transform 1 0 10980 0 -1 21616
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL56580x103360
timestamp 1586547711
transform 1 0 11716 0 -1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL63020x103360
timestamp 1586547711
transform 1 0 13004 0 -1 21616
box 0 -48 368 592
use sky130_fd_sc_hd__a21bo_4  _330_
timestamp 1586547711
transform 1 0 11808 0 -1 21616
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_1  FILL64860x103360
timestamp 1586547711
transform 1 0 13372 0 -1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL69920x103360
timestamp 1586547711
transform 1 0 14384 0 -1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_452
timestamp 1586547711
transform 1 0 13464 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1586547711
transform 1 0 14476 0 -1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL66240x103360
timestamp 1586547711
transform 1 0 13648 0 -1 21616
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL70840x103360
timestamp 1586547711
transform 1 0 14568 0 -1 21616
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1066
timestamp 1586547711
transform 1 0 15304 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_276
timestamp 1586547711
transform 1 0 15856 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_642
timestamp 1586547711
transform 1 0 16040 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL75440x103360
timestamp 1586547711
transform 1 0 15488 0 -1 21616
box 0 -48 368 592
use sky130_fd_sc_hd__o22ai_4  _455_
timestamp 1586547711
transform 1 0 16224 0 -1 21616
box 0 -48 1472 592
use sky130_fd_sc_hd__decap_3  FILL92000x103360
timestamp 1586547711
transform 1 0 18800 0 -1 21616
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1062
timestamp 1586547711
transform 1 0 19076 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL86480x103360
timestamp 1586547711
transform 1 0 17696 0 -1 21616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL94300x103360
timestamp 1586547711
transform 1 0 19260 0 -1 21616
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL97980x103360
timestamp 1586547711
transform 1 0 19996 0 -1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL100740x103360
timestamp 1586547711
transform 1 0 20548 0 -1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_149
timestamp 1586547711
transform 1 0 20180 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_920
timestamp 1586547711
transform 1 0 20364 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1586547711
transform 1 0 20088 0 -1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__a211o_4  _434_
timestamp 1586547711
transform 1 0 20640 0 -1 21616
box 0 -48 1288 592
use sky130_fd_sc_hd__a211o_4  _429_
timestamp 1586547711
transform 1 0 22664 0 -1 21616
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_8  FILL107640x103360
timestamp 1586547711
transform 1 0 21928 0 -1 21616
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL119600x103360
timestamp 1586547711
transform 1 0 24320 0 -1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_155
timestamp 1586547711
transform 1 0 24412 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_932
timestamp 1586547711
transform 1 0 24596 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1586547711
transform 1 0 25700 0 -1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL117760x103360
timestamp 1586547711
transform 1 0 23952 0 -1 21616
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL125580x103360
timestamp 1586547711
transform 1 0 25516 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL126960x103360
timestamp 1586547711
transform 1 0 25792 0 -1 21616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL121900x103360
timestamp 1586547711
transform 1 0 24780 0 -1 21616
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1586547711
transform 1 0 26988 0 -1 21616
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL132480x103360
timestamp 1586547711
transform 1 0 26896 0 -1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1586547711
transform 1 0 400 0 -1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL1380x108800
timestamp 1586547711
transform 1 0 676 0 -1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1586547711
transform 1 0 400 0 1 21616
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL3680x108800
timestamp 1586547711
transform 1 0 1136 0 -1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL1380x106080
timestamp 1586547711
transform 1 0 676 0 1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1334
timestamp 1586547711
transform 1 0 952 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1327
timestamp 1586547711
transform 1 0 1228 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1014
timestamp 1586547711
transform 1 0 768 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen0
timestamp 1586547711
transform 1 0 1412 0 -1 22704
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1333
timestamp 1586547711
transform 1 0 2056 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL9200x108800
timestamp 1586547711
transform 1 0 2240 0 -1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[8\].id.delayenb0
timestamp 1586547711
transform 1 0 952 0 1 21616
box 0 -48 1656 592
use sky130_fd_sc_hd__decap_3  FILL12880x108800
timestamp 1586547711
transform 1 0 2976 0 -1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILL14720x108800
timestamp 1586547711
transform 1 0 3344 0 -1 22704
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1586547711
transform 1 0 3252 0 -1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL17480x108800
timestamp 1586547711
transform 1 0 3896 0 -1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1197
timestamp 1586547711
transform 1 0 4264 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1208
timestamp 1586547711
transform 1 0 3712 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1194
timestamp 1586547711
transform 1 0 3896 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_987
timestamp 1586547711
transform 1 0 4080 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL20240x108800
timestamp 1586547711
transform 1 0 4448 0 -1 22704
box 0 -48 552 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp 1586547711
transform 1 0 3988 0 -1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[10\].id.delayenb1
timestamp 1586547711
transform 1 0 4264 0 1 21616
box 0 -48 1012 592
use sky130_fd_sc_hd__decap_12  FILL11040x106080
timestamp 1586547711
transform 1 0 2608 0 1 21616
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1198
timestamp 1586547711
transform 1 0 5276 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1200
timestamp 1586547711
transform 1 0 5460 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL26220x106080
timestamp 1586547711
transform 1 0 5644 0 1 21616
box 0 -48 368 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[10\].id.delayint0
timestamp 1586547711
transform 1 0 5000 0 -1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1206
timestamp 1586547711
transform 1 0 6472 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1223
timestamp 1586547711
transform 1 0 6656 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1586547711
transform 1 0 6012 0 1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[11\].id.delaybuf0
timestamp 1586547711
transform 1 0 6104 0 1 21616
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL24380x108800
timestamp 1586547711
transform 1 0 5276 0 -1 22704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL29900x108800
timestamp 1586547711
transform 1 0 6380 0 -1 22704
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL34040x106080
timestamp 1586547711
transform 1 0 7208 0 1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_426
timestamp 1586547711
transform 1 0 7668 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_92
timestamp 1586547711
transform 1 0 7300 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_42
timestamp 1586547711
transform 1 0 7484 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL32200x106080
timestamp 1586547711
transform 1 0 6840 0 1 21616
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL35420x108800
timestamp 1586547711
transform 1 0 7484 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILL40940x108800
timestamp 1586547711
transform 1 0 8588 0 -1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1586547711
transform 1 0 8864 0 -1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL37260x108800
timestamp 1586547711
transform 1 0 7852 0 -1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL42320x106080
timestamp 1586547711
transform 1 0 8864 0 1 21616
box 0 -48 736 592
use sky130_fd_sc_hd__a21bo_4  _322_
timestamp 1586547711
transform 1 0 7668 0 1 21616
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_3  FILL46000x106080
timestamp 1586547711
transform 1 0 9600 0 1 21616
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1243
timestamp 1586547711
transform 1 0 9876 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1242
timestamp 1586547711
transform 1 0 10060 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_959
timestamp 1586547711
transform 1 0 10888 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen1
timestamp 1586547711
transform 1 0 10244 0 1 21616
box 0 -48 644 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp 1586547711
transform 1 0 10796 0 -1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL42780x108800
timestamp 1586547711
transform 1 0 8956 0 -1 22704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL48300x108800
timestamp 1586547711
transform 1 0 10060 0 -1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1241
timestamp 1586547711
transform 1 0 11072 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_996
timestamp 1586547711
transform 1 0 11256 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_960
timestamp 1586547711
transform 1 0 11440 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1586547711
transform 1 0 11624 0 1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[2\].id.delayenb1
timestamp 1586547711
transform 1 0 11716 0 1 21616
box 0 -48 1012 592
use sky130_fd_sc_hd__decap_8  FILL53360x108800
timestamp 1586547711
transform 1 0 11072 0 -1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1244
timestamp 1586547711
transform 1 0 12728 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1249
timestamp 1586547711
transform 1 0 12912 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1253
timestamp 1586547711
transform 1 0 13096 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[2\].id.delayenb0
timestamp 1586547711
transform 1 0 11808 0 -1 22704
box 0 -48 1656 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1254
timestamp 1586547711
transform 1 0 13280 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1245
timestamp 1586547711
transform 1 0 13740 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[2\].id.delayint0
timestamp 1586547711
transform 1 0 13464 0 1 21616
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL65320x108800
timestamp 1586547711
transform 1 0 13464 0 -1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL69000x108800
timestamp 1586547711
transform 1 0 14200 0 -1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1247
timestamp 1586547711
transform 1 0 13924 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL68540x106080
timestamp 1586547711
transform 1 0 14108 0 1 21616
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1586547711
transform 1 0 14476 0 -1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL70840x108800
timestamp 1586547711
transform 1 0 14568 0 -1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL71300x106080
timestamp 1586547711
transform 1 0 14660 0 1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1083
timestamp 1586547711
transform 1 0 14752 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_691
timestamp 1586547711
transform 1 0 14936 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_651
timestamp 1586547711
transform 1 0 15120 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_746
timestamp 1586547711
transform 1 0 15304 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL75440x108800
timestamp 1586547711
transform 1 0 15488 0 -1 22704
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_116
timestamp 1586547711
transform 1 0 16500 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_252
timestamp 1586547711
transform 1 0 16684 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_689
timestamp 1586547711
transform 1 0 17052 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1586547711
transform 1 0 17236 0 1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL82340x106080
timestamp 1586547711
transform 1 0 16868 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _447_
timestamp 1586547711
transform 1 0 17328 0 1 21616
box 0 -48 644 592
use sky130_fd_sc_hd__o22ai_4  _443_
timestamp 1586547711
transform 1 0 15856 0 -1 22704
box 0 -48 1472 592
use sky130_fd_sc_hd__a21oi_4  _467_
timestamp 1586547711
transform 1 0 15304 0 1 21616
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_12  FILL84640x108800
timestamp 1586547711
transform 1 0 17328 0 -1 22704
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_253
timestamp 1586547711
transform 1 0 17972 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_277
timestamp 1586547711
transform 1 0 18156 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL89700x106080
timestamp 1586547711
transform 1 0 18340 0 1 21616
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILL90160x108800
timestamp 1586547711
transform 1 0 18432 0 -1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1064
timestamp 1586547711
transform 1 0 18524 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1038
timestamp 1586547711
transform 1 0 19076 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_921
timestamp 1586547711
transform 1 0 18708 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_105
timestamp 1586547711
transform 1 0 18892 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL91540x108800
timestamp 1586547711
transform 1 0 18708 0 -1 22704
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILL94300x108800
timestamp 1586547711
transform 1 0 19260 0 -1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__dfrtp_4  _561_
timestamp 1586547711
transform 1 0 19076 0 1 21616
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_3  FILL103960x106080
timestamp 1586547711
transform 1 0 21192 0 1 21616
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL97980x108800
timestamp 1586547711
transform 1 0 19996 0 -1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_663
timestamp 1586547711
transform 1 0 21468 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1586547711
transform 1 0 20088 0 -1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _427_
timestamp 1586547711
transform 1 0 21468 0 -1 22704
box 0 -48 460 592
use sky130_fd_sc_hd__buf_4  _538_
timestamp 1586547711
transform 1 0 20180 0 -1 22704
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL101660x108800
timestamp 1586547711
transform 1 0 20732 0 -1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL109020x106080
timestamp 1586547711
transform 1 0 22204 0 1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_665
timestamp 1586547711
transform 1 0 21652 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1050
timestamp 1586547711
transform 1 0 22296 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_669
timestamp 1586547711
transform 1 0 22480 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL107180x106080
timestamp 1586547711
transform 1 0 21836 0 1 21616
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILL107640x108800
timestamp 1586547711
transform 1 0 21928 0 -1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL112700x106080
timestamp 1586547711
transform 1 0 22940 0 1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_917
timestamp 1586547711
transform 1 0 23308 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1036
timestamp 1586547711
transform 1 0 23492 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1053
timestamp 1586547711
transform 1 0 23676 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_664
timestamp 1586547711
transform 1 0 22664 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_101
timestamp 1586547711
transform 1 0 23032 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1586547711
transform 1 0 22848 0 1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _428_
timestamp 1586547711
transform 1 0 22664 0 -1 22704
box 0 -48 644 592
use sky130_fd_sc_hd__dfrtp_4  _559_
timestamp 1586547711
transform 1 0 23216 0 1 21616
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_3  FILL117300x108800
timestamp 1586547711
transform 1 0 23860 0 -1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL119600x108800
timestamp 1586547711
transform 1 0 24320 0 -1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1088
timestamp 1586547711
transform 1 0 24136 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1586547711
transform 1 0 25700 0 -1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _544_
timestamp 1586547711
transform 1 0 24412 0 -1 22704
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL126960x108800
timestamp 1586547711
transform 1 0 25792 0 -1 22704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL124660x106080
timestamp 1586547711
transform 1 0 25332 0 1 21616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL122820x108800
timestamp 1586547711
transform 1 0 24964 0 -1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1586547711
transform 1 0 26988 0 -1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1586547711
transform 1 0 26988 0 1 21616
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL132480x108800
timestamp 1586547711
transform 1 0 26896 0 -1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL130180x106080
timestamp 1586547711
transform 1 0 26436 0 1 21616
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1586547711
transform 1 0 400 0 1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL1380x111520
timestamp 1586547711
transform 1 0 676 0 1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_981
timestamp 1586547711
transform 1 0 768 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_980
timestamp 1586547711
transform 1 0 952 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1328
timestamp 1586547711
transform 1 0 2148 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1329
timestamp 1586547711
transform 1 0 2332 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL10580x111520
timestamp 1586547711
transform 1 0 2516 0 1 22704
box 0 -48 368 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[8\].id.delayenb1
timestamp 1586547711
transform 1 0 1136 0 1 22704
box 0 -48 1012 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1326
timestamp 1586547711
transform 1 0 3160 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp 1586547711
transform 1 0 2884 0 1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL15640x111520
timestamp 1586547711
transform 1 0 3528 0 1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1337
timestamp 1586547711
transform 1 0 3344 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1209
timestamp 1586547711
transform 1 0 3804 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL19780x111520
timestamp 1586547711
transform 1 0 4356 0 1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1205
timestamp 1586547711
transform 1 0 3988 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_945
timestamp 1586547711
transform 1 0 4172 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1204
timestamp 1586547711
transform 1 0 4448 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen0
timestamp 1586547711
transform 1 0 4632 0 1 22704
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_944
timestamp 1586547711
transform 1 0 5276 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1199
timestamp 1586547711
transform 1 0 5460 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1586547711
transform 1 0 6012 0 1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL26220x111520
timestamp 1586547711
transform 1 0 5644 0 1 22704
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL28520x111520
timestamp 1586547711
transform 1 0 6104 0 1 22704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL34040x111520
timestamp 1586547711
transform 1 0 7208 0 1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_974
timestamp 1586547711
transform 1 0 7484 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1232
timestamp 1586547711
transform 1 0 7668 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1234
timestamp 1586547711
transform 1 0 7852 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL38180x111520
timestamp 1586547711
transform 1 0 8036 0 1 22704
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL43700x111520
timestamp 1586547711
transform 1 0 9140 0 1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1182
timestamp 1586547711
transform 1 0 9600 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1190
timestamp 1586547711
transform 1 0 9784 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1236
timestamp 1586547711
transform 1 0 10704 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1251
timestamp 1586547711
transform 1 0 10888 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL47840x111520
timestamp 1586547711
transform 1 0 9968 0 1 22704
box 0 -48 368 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[0\].id.delaybuf0
timestamp 1586547711
transform 1 0 9232 0 1 22704
box 0 -48 368 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[2\].id.delaybuf0
timestamp 1586547711
transform 1 0 10336 0 1 22704
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILL56580x111520
timestamp 1586547711
transform 1 0 11716 0 1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1246
timestamp 1586547711
transform 1 0 11808 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_994
timestamp 1586547711
transform 1 0 11992 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_434
timestamp 1586547711
transform 1 0 12176 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_43
timestamp 1586547711
transform 1 0 12360 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen0
timestamp 1586547711
transform 1 0 12544 0 1 22704
box 0 -48 644 592
use sky130_fd_sc_hd__decap_6  FILL53360x111520
timestamp 1586547711
transform 1 0 11072 0 1 22704
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1586547711
transform 1 0 11624 0 1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_91
timestamp 1586547711
transform 1 0 13188 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_995
timestamp 1586547711
transform 1 0 13372 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1248
timestamp 1586547711
transform 1 0 13556 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL66700x111520
timestamp 1586547711
transform 1 0 13740 0 1 22704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL72220x111520
timestamp 1586547711
transform 1 0 14844 0 1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL75900x111520
timestamp 1586547711
transform 1 0 15580 0 1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1082
timestamp 1586547711
transform 1 0 15856 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_251
timestamp 1586547711
transform 1 0 16500 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_275
timestamp 1586547711
transform 1 0 16684 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1063
timestamp 1586547711
transform 1 0 16868 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL84640x111520
timestamp 1586547711
transform 1 0 17328 0 1 22704
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1586547711
transform 1 0 17236 0 1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL83260x111520
timestamp 1586547711
transform 1 0 17052 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _273_
timestamp 1586547711
transform 1 0 16040 0 1 22704
box 0 -48 460 592
use sky130_fd_sc_hd__fill_1  FILL90160x111520
timestamp 1586547711
transform 1 0 18432 0 1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1065
timestamp 1586547711
transform 1 0 17880 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_657
timestamp 1586547711
transform 1 0 18064 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_679
timestamp 1586547711
transform 1 0 18248 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_655
timestamp 1586547711
transform 1 0 19168 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_658
timestamp 1586547711
transform 1 0 19352 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _425_
timestamp 1586547711
transform 1 0 18524 0 1 22704
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  FILL99360x111520
timestamp 1586547711
transform 1 0 20272 0 1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_659
timestamp 1586547711
transform 1 0 20548 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_662
timestamp 1586547711
transform 1 0 20732 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1069
timestamp 1586547711
transform 1 0 20916 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL103500x111520
timestamp 1586547711
transform 1 0 21100 0 1 22704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL95680x111520
timestamp 1586547711
transform 1 0 19536 0 1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL111780x111520
timestamp 1586547711
transform 1 0 22756 0 1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL116380x111520
timestamp 1586547711
transform 1 0 23676 0 1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL109020x111520
timestamp 1586547711
transform 1 0 22204 0 1 22704
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1586547711
transform 1 0 22848 0 1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL112700x111520
timestamp 1586547711
transform 1 0 22940 0 1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_933
timestamp 1586547711
transform 1 0 23768 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1586547711
transform 1 0 23952 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _567_
timestamp 1586547711
transform 1 0 24136 0 1 22704
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1586547711
transform 1 0 26988 0 1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL129260x111520
timestamp 1586547711
transform 1 0 26252 0 1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1586547711
transform 1 0 400 0 -1 23792
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_590
timestamp 1586547711
transform 1 0 860 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1339
timestamp 1586547711
transform 1 0 1872 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen1
timestamp 1586547711
transform 1 0 1228 0 -1 23792
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILL1380x114240
timestamp 1586547711
transform 1 0 676 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL3220x114240
timestamp 1586547711
transform 1 0 1044 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL8280x114240
timestamp 1586547711
transform 1 0 2056 0 -1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL13800x114240
timestamp 1586547711
transform 1 0 3160 0 -1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL18400x114240
timestamp 1586547711
transform 1 0 4080 0 -1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1586547711
transform 1 0 3252 0 -1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[10\].id.delayenb0
timestamp 1586547711
transform 1 0 4172 0 -1 23792
box 0 -48 1656 592
use sky130_fd_sc_hd__decap_8  FILL14720x114240
timestamp 1586547711
transform 1 0 3344 0 -1 23792
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILL27140x114240
timestamp 1586547711
transform 1 0 5828 0 -1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen0
timestamp 1586547711
transform 1 0 7484 0 -1 23792
box 0 -48 644 592
use sky130_fd_sc_hd__decap_6  FILL32660x114240
timestamp 1586547711
transform 1 0 6932 0 -1 23792
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1586547711
transform 1 0 8864 0 -1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL38640x114240
timestamp 1586547711
transform 1 0 8128 0 -1 23792
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILL42780x114240
timestamp 1586547711
transform 1 0 8956 0 -1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL48300x114240
timestamp 1586547711
transform 1 0 10060 0 -1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL59340x114240
timestamp 1586547711
transform 1 0 12268 0 -1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__a21bo_4  _326_
timestamp 1586547711
transform 1 0 12360 0 -1 23792
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_12  FILL53820x114240
timestamp 1586547711
transform 1 0 11164 0 -1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL70840x114240
timestamp 1586547711
transform 1 0 14568 0 -1 23792
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_138
timestamp 1586547711
transform 1 0 14844 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_898
timestamp 1586547711
transform 1 0 15028 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1586547711
transform 1 0 14476 0 -1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL69460x114240
timestamp 1586547711
transform 1 0 14292 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL65780x114240
timestamp 1586547711
transform 1 0 13556 0 -1 23792
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL74060x114240
timestamp 1586547711
transform 1 0 15212 0 -1 23792
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL77740x114240
timestamp 1586547711
transform 1 0 15948 0 -1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _279_
timestamp 1586547711
transform 1 0 16040 0 -1 23792
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL80500x114240
timestamp 1586547711
transform 1 0 16500 0 -1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL87860x114240
timestamp 1586547711
transform 1 0 17972 0 -1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL86020x114240
timestamp 1586547711
transform 1 0 17604 0 -1 23792
box 0 -48 368 592
use sky130_fd_sc_hd__nor2_4  _436_
timestamp 1586547711
transform 1 0 18064 0 -1 23792
box 0 -48 828 592
use sky130_fd_sc_hd__decap_12  FILL92460x114240
timestamp 1586547711
transform 1 0 18892 0 -1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL97980x114240
timestamp 1586547711
transform 1 0 19996 0 -1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1071
timestamp 1586547711
transform 1 0 21192 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1086
timestamp 1586547711
transform 1 0 21376 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1586547711
transform 1 0 20088 0 -1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL98900x114240
timestamp 1586547711
transform 1 0 20180 0 -1 23792
box 0 -48 368 592
use sky130_fd_sc_hd__and2_4  _426_
timestamp 1586547711
transform 1 0 20548 0 -1 23792
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL105800x114240
timestamp 1586547711
transform 1 0 21560 0 -1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL111320x114240
timestamp 1586547711
transform 1 0 22664 0 -1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL119600x114240
timestamp 1586547711
transform 1 0 24320 0 -1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1044
timestamp 1586547711
transform 1 0 24136 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_934
timestamp 1586547711
transform 1 0 24412 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1586547711
transform 1 0 25700 0 -1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL116840x114240
timestamp 1586547711
transform 1 0 23768 0 -1 23792
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL120980x114240
timestamp 1586547711
transform 1 0 24596 0 -1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL126960x114240
timestamp 1586547711
transform 1 0 25792 0 -1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1586547711
transform 1 0 26988 0 -1 23792
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL132480x114240
timestamp 1586547711
transform 1 0 26896 0 -1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1586547711
transform 1 0 400 0 1 23792
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_63
timestamp 1586547711
transform 1 0 676 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _404_
timestamp 1586547711
transform 1 0 860 0 1 23792
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_8  FILL8280x116960
timestamp 1586547711
transform 1 0 2056 0 1 23792
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1335
timestamp 1586547711
transform 1 0 3160 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1347
timestamp 1586547711
transform 1 0 3344 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1201
timestamp 1586547711
transform 1 0 4080 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1207
timestamp 1586547711
transform 1 0 4264 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL15640x116960
timestamp 1586547711
transform 1 0 3528 0 1 23792
box 0 -48 552 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[9\].id.delaybuf0
timestamp 1586547711
transform 1 0 2792 0 1 23792
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILL20240x116960
timestamp 1586547711
transform 1 0 4448 0 1 23792
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL23920x116960
timestamp 1586547711
transform 1 0 5184 0 1 23792
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL31280x116960
timestamp 1586547711
transform 1 0 6656 0 1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_52
timestamp 1586547711
transform 1 0 5460 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_83
timestamp 1586547711
transform 1 0 5644 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_371
timestamp 1586547711
transform 1 0 5828 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_943
timestamp 1586547711
transform 1 0 6104 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1239
timestamp 1586547711
transform 1 0 6748 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1586547711
transform 1 0 6012 0 1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL29440x116960
timestamp 1586547711
transform 1 0 6288 0 1 23792
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1233
timestamp 1586547711
transform 1 0 6932 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1231
timestamp 1586547711
transform 1 0 7116 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_975
timestamp 1586547711
transform 1 0 7300 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[1\].id.delayenb0
timestamp 1586547711
transform 1 0 7484 0 1 23792
box 0 -48 1656 592
use sky130_fd_sc_hd__fill_1  FILL47380x116960
timestamp 1586547711
transform 1 0 9876 0 1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_941
timestamp 1586547711
transform 1 0 9968 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1180
timestamp 1586547711
transform 1 0 10152 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1187
timestamp 1586547711
transform 1 0 10336 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL43700x116960
timestamp 1586547711
transform 1 0 9140 0 1 23792
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL50600x116960
timestamp 1586547711
transform 1 0 10520 0 1 23792
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL54280x116960
timestamp 1586547711
transform 1 0 11256 0 1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL55660x116960
timestamp 1586547711
transform 1 0 11532 0 1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1179
timestamp 1586547711
transform 1 0 11348 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1181
timestamp 1586547711
transform 1 0 11716 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1586547711
transform 1 0 11624 0 1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL57500x116960
timestamp 1586547711
transform 1 0 11900 0 1 23792
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILL59340x116960
timestamp 1586547711
transform 1 0 12268 0 1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1175
timestamp 1586547711
transform 1 0 12360 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1191
timestamp 1586547711
transform 1 0 12544 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL61640x116960
timestamp 1586547711
transform 1 0 12728 0 1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1027
timestamp 1586547711
transform 1 0 13832 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_899
timestamp 1586547711
transform 1 0 14016 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_117
timestamp 1586547711
transform 1 0 14200 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _550_
timestamp 1586547711
transform 1 0 14384 0 1 23792
box 0 -48 2116 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1586547711
transform 1 0 17236 0 1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL84640x116960
timestamp 1586547711
transform 1 0 17328 0 1 23792
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILL80500x116960
timestamp 1586547711
transform 1 0 16500 0 1 23792
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL86480x116960
timestamp 1586547711
transform 1 0 17696 0 1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_261
timestamp 1586547711
transform 1 0 17788 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_638
timestamp 1586547711
transform 1 0 17972 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_660
timestamp 1586547711
transform 1 0 18156 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_680
timestamp 1586547711
transform 1 0 18340 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_681
timestamp 1586547711
transform 1 0 18524 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL91540x116960
timestamp 1586547711
transform 1 0 18708 0 1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_684
timestamp 1586547711
transform 1 0 19996 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_281
timestamp 1586547711
transform 1 0 20180 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_263
timestamp 1586547711
transform 1 0 20364 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL97060x116960
timestamp 1586547711
transform 1 0 19812 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__a21oi_4  _446_
timestamp 1586547711
transform 1 0 20548 0 1 23792
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_1  FILL115460x116960
timestamp 1586547711
transform 1 0 23492 0 1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_683
timestamp 1586547711
transform 1 0 21744 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_279
timestamp 1586547711
transform 1 0 22296 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1085
timestamp 1586547711
transform 1 0 22480 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1093
timestamp 1586547711
transform 1 0 23584 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL112700x116960
timestamp 1586547711
transform 1 0 22940 0 1 23792
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1586547711
transform 1 0 22848 0 1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL107640x116960
timestamp 1586547711
transform 1 0 21928 0 1 23792
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL111320x116960
timestamp 1586547711
transform 1 0 22664 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_630
timestamp 1586547711
transform 1 0 23768 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_156
timestamp 1586547711
transform 1 0 23952 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__xor2_4  _419_
timestamp 1586547711
transform 1 0 24136 0 1 23792
box 0 -48 2024 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1586547711
transform 1 0 26988 0 1 23792
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL132480x116960
timestamp 1586547711
transform 1 0 26896 0 1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL128800x116960
timestamp 1586547711
transform 1 0 26160 0 1 23792
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1586547711
transform 1 0 400 0 -1 24880
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_72
timestamp 1586547711
transform 1 0 860 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_979
timestamp 1586547711
transform 1 0 1044 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1343
timestamp 1586547711
transform 1 0 1228 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1350
timestamp 1586547711
transform 1 0 1412 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL1380x119680
timestamp 1586547711
transform 1 0 676 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL5980x119680
timestamp 1586547711
transform 1 0 1596 0 -1 24880
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILL11500x119680
timestamp 1586547711
transform 1 0 2700 0 -1 24880
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1586547711
transform 1 0 3252 0 -1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[10\].id.delaybuf0
timestamp 1586547711
transform 1 0 4080 0 -1 24880
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILL14720x119680
timestamp 1586547711
transform 1 0 3344 0 -1 24880
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL20240x119680
timestamp 1586547711
transform 1 0 4448 0 -1 24880
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL23920x119680
timestamp 1586547711
transform 1 0 5184 0 -1 24880
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_957
timestamp 1586547711
transform 1 0 6656 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _348_
timestamp 1586547711
transform 1 0 5460 0 -1 24880
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_3  FILL40940x119680
timestamp 1586547711
transform 1 0 8588 0 -1 24880
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1240
timestamp 1586547711
transform 1 0 6840 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1235
timestamp 1586547711
transform 1 0 7668 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1586547711
transform 1 0 8864 0 -1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL33120x119680
timestamp 1586547711
transform 1 0 7024 0 -1 24880
box 0 -48 368 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[1\].id.delayint0
timestamp 1586547711
transform 1 0 7392 0 -1 24880
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL37260x119680
timestamp 1586547711
transform 1 0 7852 0 -1 24880
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL46460x119680
timestamp 1586547711
transform 1 0 9692 0 -1 24880
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_940
timestamp 1586547711
transform 1 0 9140 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_942
timestamp 1586547711
transform 1 0 9324 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1192
timestamp 1586547711
transform 1 0 9508 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen0
timestamp 1586547711
transform 1 0 9968 0 -1 24880
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILL42780x119680
timestamp 1586547711
transform 1 0 8956 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL51060x119680
timestamp 1586547711
transform 1 0 10612 0 -1 24880
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_952
timestamp 1586547711
transform 1 0 11624 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_954
timestamp 1586547711
transform 1 0 11808 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1178
timestamp 1586547711
transform 1 0 11992 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL58880x119680
timestamp 1586547711
transform 1 0 12176 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[0\].id.delayint0
timestamp 1586547711
transform 1 0 11348 0 -1 24880
box 0 -48 276 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1
timestamp 1586547711
transform 1 0 12360 0 -1 24880
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL61180x119680
timestamp 1586547711
transform 1 0 12636 0 -1 24880
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL71760x119680
timestamp 1586547711
transform 1 0 14752 0 -1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1084
timestamp 1586547711
transform 1 0 14568 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1586547711
transform 1 0 14476 0 -1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _527_
timestamp 1586547711
transform 1 0 14844 0 -1 24880
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL66700x119680
timestamp 1586547711
transform 1 0 13740 0 -1 24880
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL84180x119680
timestamp 1586547711
transform 1 0 17236 0 -1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1040
timestamp 1586547711
transform 1 0 17328 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL74980x119680
timestamp 1586547711
transform 1 0 15396 0 -1 24880
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL80500x119680
timestamp 1586547711
transform 1 0 16500 0 -1 24880
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL85560x119680
timestamp 1586547711
transform 1 0 17512 0 -1 24880
box 0 -48 276 592
use sky130_fd_sc_hd__a211o_4  _437_
timestamp 1586547711
transform 1 0 17788 0 -1 24880
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_8  FILL93380x119680
timestamp 1586547711
transform 1 0 19076 0 -1 24880
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL97060x119680
timestamp 1586547711
transform 1 0 19812 0 -1 24880
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL98900x119680
timestamp 1586547711
transform 1 0 20180 0 -1 24880
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL102120x119680
timestamp 1586547711
transform 1 0 20824 0 -1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_280
timestamp 1586547711
transform 1 0 20456 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_686
timestamp 1586547711
transform 1 0 20640 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1028
timestamp 1586547711
transform 1 0 21560 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1586547711
transform 1 0 20088 0 -1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _445_
timestamp 1586547711
transform 1 0 20916 0 -1 24880
box 0 -48 644 592
use sky130_fd_sc_hd__decap_6  FILL106720x119680
timestamp 1586547711
transform 1 0 21744 0 -1 24880
box 0 -48 552 592
use sky130_fd_sc_hd__inv_4  _280_
timestamp 1586547711
transform 1 0 22296 0 -1 24880
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL111780x119680
timestamp 1586547711
transform 1 0 22756 0 -1 24880
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL118220x119680
timestamp 1586547711
transform 1 0 24044 0 -1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL119600x119680
timestamp 1586547711
transform 1 0 24320 0 -1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1091
timestamp 1586547711
transform 1 0 23860 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1090
timestamp 1586547711
transform 1 0 24136 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1586547711
transform 1 0 25700 0 -1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _545_
timestamp 1586547711
transform 1 0 24412 0 -1 24880
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL126960x119680
timestamp 1586547711
transform 1 0 25792 0 -1 24880
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL122820x119680
timestamp 1586547711
transform 1 0 24964 0 -1 24880
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1586547711
transform 1 0 26988 0 -1 24880
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL132480x119680
timestamp 1586547711
transform 1 0 26896 0 -1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1586547711
transform 1 0 400 0 1 24880
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL1380x122400
timestamp 1586547711
transform 1 0 676 0 1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1342
timestamp 1586547711
transform 1 0 768 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1341
timestamp 1586547711
transform 1 0 952 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_983
timestamp 1586547711
transform 1 0 1780 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_984
timestamp 1586547711
transform 1 0 1964 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen1
timestamp 1586547711
transform 1 0 1136 0 1 24880
box 0 -48 644 592
use sky130_fd_sc_hd__decap_4  FILL8740x122400
timestamp 1586547711
transform 1 0 2148 0 1 24880
box 0 -48 368 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[9\].id.delayint0
timestamp 1586547711
transform 1 0 2516 0 1 24880
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1344
timestamp 1586547711
transform 1 0 2792 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1346
timestamp 1586547711
transform 1 0 2976 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1017
timestamp 1586547711
transform 1 0 3344 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1203
timestamp 1586547711
transform 1 0 3528 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1349
timestamp 1586547711
transform 1 0 3712 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL13800x122400
timestamp 1586547711
transform 1 0 3160 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL17480x122400
timestamp 1586547711
transform 1 0 3896 0 1 24880
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL27600x122400
timestamp 1586547711
transform 1 0 5920 0 1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL28520x122400
timestamp 1586547711
transform 1 0 6104 0 1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_955
timestamp 1586547711
transform 1 0 5184 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_553
timestamp 1586547711
transform 1 0 5368 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_79
timestamp 1586547711
transform 1 0 5552 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_56
timestamp 1586547711
transform 1 0 5736 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1586547711
transform 1 0 6012 0 1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL23000x122400
timestamp 1586547711
transform 1 0 5000 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[1\].id.delayenb1
timestamp 1586547711
transform 1 0 6196 0 1 24880
box 0 -48 1012 592
use sky130_fd_sc_hd__fill_1  FILL34960x122400
timestamp 1586547711
transform 1 0 7392 0 1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1230
timestamp 1586547711
transform 1 0 7208 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1238
timestamp 1586547711
transform 1 0 7484 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL37260x122400
timestamp 1586547711
transform 1 0 7852 0 1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1227
timestamp 1586547711
transform 1 0 7668 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1189
timestamp 1586547711
transform 1 0 7944 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[1\].id.delaybuf0
timestamp 1586547711
transform 1 0 8128 0 1 24880
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1188
timestamp 1586547711
transform 1 0 8496 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_315
timestamp 1586547711
transform 1 0 8680 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_93
timestamp 1586547711
transform 1 0 8864 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_41
timestamp 1586547711
transform 1 0 9048 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1193
timestamp 1586547711
transform 1 0 10888 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[0\].id.delayenb0
timestamp 1586547711
transform 1 0 9232 0 1 24880
box 0 -48 1656 592
use sky130_fd_sc_hd__diode_2  ANTENNA_499
timestamp 1586547711
transform 1 0 11072 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_80
timestamp 1586547711
transform 1 0 11256 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_55
timestamp 1586547711
transform 1 0 11440 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1586547711
transform 1 0 11624 0 1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[0\].id.delayenb1
timestamp 1586547711
transform 1 0 11716 0 1 24880
box 0 -48 1012 592
use sky130_fd_sc_hd__decap_12  FILL61640x122400
timestamp 1586547711
transform 1 0 12728 0 1 24880
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL72680x122400
timestamp 1586547711
transform 1 0 14936 0 1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1067
timestamp 1586547711
transform 1 0 14200 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1039
timestamp 1586547711
transform 1 0 14384 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_107
timestamp 1586547711
transform 1 0 14568 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_923
timestamp 1586547711
transform 1 0 14752 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL67160x122400
timestamp 1586547711
transform 1 0 13832 0 1 24880
box 0 -48 368 592
use sky130_fd_sc_hd__buf_4  _539_
timestamp 1586547711
transform 1 0 15028 0 1 24880
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_150
timestamp 1586547711
transform 1 0 15580 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_922
timestamp 1586547711
transform 1 0 15764 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1072
timestamp 1586547711
transform 1 0 16684 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_109
timestamp 1586547711
transform 1 0 16868 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_108
timestamp 1586547711
transform 1 0 17052 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1586547711
transform 1 0 17236 0 1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _563_
timestamp 1586547711
transform 1 0 17328 0 1 24880
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_8  FILL77740x122400
timestamp 1586547711
transform 1 0 15948 0 1 24880
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_647
timestamp 1586547711
transform 1 0 19444 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL97060x122400
timestamp 1586547711
transform 1 0 19812 0 1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_661
timestamp 1586547711
transform 1 0 19628 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_643
timestamp 1586547711
transform 1 0 19904 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_119
timestamp 1586547711
transform 1 0 20088 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_118
timestamp 1586547711
transform 1 0 20272 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__o22ai_4  _444_
timestamp 1586547711
transform 1 0 20456 0 1 24880
box 0 -48 1472 592
use sky130_fd_sc_hd__diode_2  ANTENNA_901
timestamp 1586547711
transform 1 0 21928 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1087
timestamp 1586547711
transform 1 0 22112 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1045
timestamp 1586547711
transform 1 0 23492 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_935
timestamp 1586547711
transform 1 0 23676 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL109480x122400
timestamp 1586547711
transform 1 0 22296 0 1 24880
box 0 -48 552 592
use sky130_fd_sc_hd__decap_6  FILL112700x122400
timestamp 1586547711
transform 1 0 22940 0 1 24880
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1586547711
transform 1 0 22848 0 1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _568_
timestamp 1586547711
transform 1 0 23860 0 1 24880
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_3  FILL131560x122400
timestamp 1586547711
transform 1 0 26712 0 1 24880
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1586547711
transform 1 0 26988 0 1 24880
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL127880x122400
timestamp 1586547711
transform 1 0 25976 0 1 24880
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1586547711
transform 1 0 400 0 1 25968
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1586547711
transform 1 0 400 0 -1 25968
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL3220x125120
timestamp 1586547711
transform 1 0 1044 0 -1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL1380x125120
timestamp 1586547711
transform 1 0 676 0 -1 25968
box 0 -48 368 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[9\].id.delayenb1
timestamp 1586547711
transform 1 0 1136 0 -1 25968
box 0 -48 1012 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1340
timestamp 1586547711
transform 1 0 2240 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1348
timestamp 1586547711
transform 1 0 2424 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL6900x127840
timestamp 1586547711
transform 1 0 1780 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp 1586547711
transform 1 0 1964 0 1 25968
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL1380x127840
timestamp 1586547711
transform 1 0 676 0 1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL8740x125120
timestamp 1586547711
transform 1 0 2148 0 -1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL11040x127840
timestamp 1586547711
transform 1 0 2608 0 1 25968
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1345
timestamp 1586547711
transform 1 0 2884 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1016
timestamp 1586547711
transform 1 0 3712 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1202
timestamp 1586547711
transform 1 0 3896 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen0
timestamp 1586547711
transform 1 0 3068 0 1 25968
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1586547711
transform 1 0 3252 0 -1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[9\].id.delayenb0
timestamp 1586547711
transform 1 0 3344 0 -1 25968
box 0 -48 1656 592
use sky130_fd_sc_hd__decap_12  FILL18400x127840
timestamp 1586547711
transform 1 0 4080 0 1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL23920x127840
timestamp 1586547711
transform 1 0 5184 0 1 25968
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL23000x125120
timestamp 1586547711
transform 1 0 5000 0 -1 25968
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL31740x127840
timestamp 1586547711
transform 1 0 6748 0 1 25968
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL27600x127840
timestamp 1586547711
transform 1 0 5920 0 1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL28520x127840
timestamp 1586547711
transform 1 0 6104 0 1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_956
timestamp 1586547711
transform 1 0 6196 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1228
timestamp 1586547711
transform 1 0 6380 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1229
timestamp 1586547711
transform 1 0 6564 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1586547711
transform 1 0 6012 0 1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__a21bo_4  _373_
timestamp 1586547711
transform 1 0 5736 0 -1 25968
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_1  FILL34500x125120
timestamp 1586547711
transform 1 0 7300 0 -1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL35880x125120
timestamp 1586547711
transform 1 0 7576 0 -1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_84
timestamp 1586547711
transform 1 0 7024 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_51
timestamp 1586547711
transform 1 0 7208 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1015
timestamp 1586547711
transform 1 0 7392 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL32660x125120
timestamp 1586547711
transform 1 0 6932 0 -1 25968
box 0 -48 368 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp 1586547711
transform 1 0 7668 0 -1 25968
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1237
timestamp 1586547711
transform 1 0 8128 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL39560x125120
timestamp 1586547711
transform 1 0 8312 0 -1 25968
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1586547711
transform 1 0 8864 0 -1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL37720x125120
timestamp 1586547711
transform 1 0 7944 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _347_
timestamp 1586547711
transform 1 0 7392 0 1 25968
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_12  FILL40940x127840
timestamp 1586547711
transform 1 0 8588 0 1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILL51980x127840
timestamp 1586547711
transform 1 0 10796 0 1 25968
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILL42780x125120
timestamp 1586547711
transform 1 0 8956 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _293_
timestamp 1586547711
transform 1 0 9140 0 -1 25968
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_12  FILL46460x127840
timestamp 1586547711
transform 1 0 9692 0 1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL49680x125120
timestamp 1586547711
transform 1 0 10336 0 -1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL54740x127840
timestamp 1586547711
transform 1 0 11348 0 1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL55200x125120
timestamp 1586547711
transform 1 0 11440 0 -1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1177
timestamp 1586547711
transform 1 0 11440 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen1
timestamp 1586547711
transform 1 0 11716 0 1 25968
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1586547711
transform 1 0 11624 0 1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_953
timestamp 1586547711
transform 1 0 12360 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1176
timestamp 1586547711
transform 1 0 12544 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _356_
timestamp 1586547711
transform 1 0 11532 0 -1 25968
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_12  FILL61640x127840
timestamp 1586547711
transform 1 0 12728 0 1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL61640x125120
timestamp 1586547711
transform 1 0 12728 0 -1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL67160x127840
timestamp 1586547711
transform 1 0 13832 0 1 25968
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL69920x125120
timestamp 1586547711
transform 1 0 14384 0 -1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1586547711
transform 1 0 14568 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_294
timestamp 1586547711
transform 1 0 14752 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL67160x125120
timestamp 1586547711
transform 1 0 13832 0 -1 25968
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1586547711
transform 1 0 14476 0 -1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _285_
timestamp 1586547711
transform 1 0 14108 0 1 25968
box 0 -48 460 592
use sky130_fd_sc_hd__dfrtp_4  _562_
timestamp 1586547711
transform 1 0 14568 0 -1 25968
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_8  FILL72680x127840
timestamp 1586547711
transform 1 0 14936 0 1 25968
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL84180x125120
timestamp 1586547711
transform 1 0 17236 0 -1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_106
timestamp 1586547711
transform 1 0 16132 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_682
timestamp 1586547711
transform 1 0 16316 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_925
timestamp 1586547711
transform 1 0 17328 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL81420x125120
timestamp 1586547711
transform 1 0 16684 0 -1 25968
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1586547711
transform 1 0 17236 0 1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL84640x127840
timestamp 1586547711
transform 1 0 17328 0 1 25968
box 0 -48 368 592
use sky130_fd_sc_hd__inv_4  _438_
timestamp 1586547711
transform 1 0 15672 0 1 25968
box 0 -48 460 592
use sky130_fd_sc_hd__decap_8  FILL80500x127840
timestamp 1586547711
transform 1 0 16500 0 1 25968
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL94760x127840
timestamp 1586547711
transform 1 0 19352 0 1 25968
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL85560x125120
timestamp 1586547711
transform 1 0 17512 0 -1 25968
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_151
timestamp 1586547711
transform 1 0 18248 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_924
timestamp 1586547711
transform 1 0 18432 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1070
timestamp 1586547711
transform 1 0 17788 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _439_
timestamp 1586547711
transform 1 0 17972 0 -1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__buf_4  _540_
timestamp 1586547711
transform 1 0 17696 0 1 25968
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL91080x127840
timestamp 1586547711
transform 1 0 18616 0 1 25968
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL93380x125120
timestamp 1586547711
transform 1 0 19076 0 -1 25968
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL97060x125120
timestamp 1586547711
transform 1 0 19812 0 -1 25968
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL98900x125120
timestamp 1586547711
transform 1 0 20180 0 -1 25968
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_260
timestamp 1586547711
transform 1 0 20088 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1068
timestamp 1586547711
transform 1 0 20272 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_262
timestamp 1586547711
transform 1 0 20456 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1586547711
transform 1 0 20088 0 -1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _275_
timestamp 1586547711
transform 1 0 19628 0 1 25968
box 0 -48 460 592
use sky130_fd_sc_hd__diode_2  ANTENNA_652
timestamp 1586547711
transform 1 0 20640 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _528_
timestamp 1586547711
transform 1 0 21560 0 1 25968
box 0 -48 552 592
use sky130_fd_sc_hd__dfrtp_4  _551_
timestamp 1586547711
transform 1 0 20824 0 -1 25968
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_12  FILL100280x127840
timestamp 1586547711
transform 1 0 20456 0 1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_139
timestamp 1586547711
transform 1 0 22112 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_900
timestamp 1586547711
transform 1 0 22296 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILL112700x127840
timestamp 1586547711
transform 1 0 22940 0 1 25968
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1586547711
transform 1 0 22848 0 1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL110400x127840
timestamp 1586547711
transform 1 0 22480 0 1 25968
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILL112700x125120
timestamp 1586547711
transform 1 0 22940 0 -1 25968
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1094
timestamp 1586547711
transform 1 0 23216 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1046
timestamp 1586547711
transform 1 0 23400 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_157
timestamp 1586547711
transform 1 0 23584 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL116380x125120
timestamp 1586547711
transform 1 0 23676 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1089
timestamp 1586547711
transform 1 0 23860 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL123740x125120
timestamp 1586547711
transform 1 0 25148 0 -1 25968
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1586547711
transform 1 0 25700 0 -1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _569_
timestamp 1586547711
transform 1 0 23768 0 1 25968
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_12  FILL118220x125120
timestamp 1586547711
transform 1 0 24044 0 -1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL126960x125120
timestamp 1586547711
transform 1 0 25792 0 -1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1586547711
transform 1 0 26988 0 1 25968
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1586547711
transform 1 0 26988 0 -1 25968
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL132480x125120
timestamp 1586547711
transform 1 0 26896 0 -1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL127420x127840
timestamp 1586547711
transform 1 0 25884 0 1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1586547711
transform 1 0 400 0 -1 27056
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL1380x130560
timestamp 1586547711
transform 1 0 676 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL6900x130560
timestamp 1586547711
transform 1 0 1780 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1586547711
transform 1 0 3252 0 -1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL12420x130560
timestamp 1586547711
transform 1 0 2884 0 -1 27056
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL14720x130560
timestamp 1586547711
transform 1 0 3344 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL20240x130560
timestamp 1586547711
transform 1 0 4448 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen1
timestamp 1586547711
transform 1 0 6196 0 -1 27056
box 0 -48 644 592
use sky130_fd_sc_hd__decap_6  FILL25760x130560
timestamp 1586547711
transform 1 0 5552 0 -1 27056
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1586547711
transform 1 0 6104 0 -1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILL41400x130560
timestamp 1586547711
transform 1 0 8680 0 -1 27056
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_438
timestamp 1586547711
transform 1 0 7392 0 -1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL32200x130560
timestamp 1586547711
transform 1 0 6840 0 -1 27056
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL35880x130560
timestamp 1586547711
transform 1 0 7576 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1586547711
transform 1 0 8956 0 -1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL43240x130560
timestamp 1586547711
transform 1 0 9048 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL48760x130560
timestamp 1586547711
transform 1 0 10152 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILL54280x130560
timestamp 1586547711
transform 1 0 11256 0 -1 27056
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1586547711
transform 1 0 11808 0 -1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL57500x130560
timestamp 1586547711
transform 1 0 11900 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL63020x130560
timestamp 1586547711
transform 1 0 13004 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILL68540x130560
timestamp 1586547711
transform 1 0 14108 0 -1 27056
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1586547711
transform 1 0 14660 0 -1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL71760x130560
timestamp 1586547711
transform 1 0 14752 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILL82800x130560
timestamp 1586547711
transform 1 0 16960 0 -1 27056
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL77280x130560
timestamp 1586547711
transform 1 0 15856 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1586547711
transform 1 0 17512 0 -1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL86020x130560
timestamp 1586547711
transform 1 0 17604 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL91540x130560
timestamp 1586547711
transform 1 0 18708 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILL97060x130560
timestamp 1586547711
transform 1 0 19812 0 -1 27056
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1586547711
transform 1 0 20364 0 -1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL100280x130560
timestamp 1586547711
transform 1 0 20456 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL105800x130560
timestamp 1586547711
transform 1 0 21560 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL116380x130560
timestamp 1586547711
transform 1 0 23676 0 -1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL111320x130560
timestamp 1586547711
transform 1 0 22664 0 -1 27056
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1586547711
transform 1 0 23216 0 -1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL114540x130560
timestamp 1586547711
transform 1 0 23308 0 -1 27056
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILL126960x130560
timestamp 1586547711
transform 1 0 25792 0 -1 27056
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1092
timestamp 1586547711
transform 1 0 23768 0 -1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL117760x130560
timestamp 1586547711
transform 1 0 23952 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL123280x130560
timestamp 1586547711
transform 1 0 25056 0 -1 27056
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1586547711
transform 1 0 26988 0 -1 27056
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL132480x130560
timestamp 1586547711
transform 1 0 26896 0 -1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1586547711
transform 1 0 26068 0 -1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL128800x130560
timestamp 1586547711
transform 1 0 26160 0 -1 27056
box 0 -48 736 592
<< labels >>
rlabel metal2 s 16384 0 16524 420 8 reset
port 0 nsew default input
rlabel metal2 s 376 0 516 420 8 extclk_sel
port 1 nsew default input
rlabel metal3 s 27303 22622 27735 22922 6 osc
port 2 nsew default input
rlabel metal3 s 0 23982 432 24282 4 clockc
port 3 nsew default tristate
rlabel metal2 s 24480 0 24620 420 8 clockp[1]
port 4 nsew default tristate
rlabel metal3 s 27303 16638 27735 16938 6 clockp[0]
port 5 nsew default tristate
rlabel metal2 s 6264 27315 6404 27735 6 clockd[3]
port 6 nsew default tristate
rlabel metal3 s 0 3038 432 3338 4 clockd[2]
port 7 nsew default tristate
rlabel metal3 s 27303 25614 27735 25914 6 clockd[1]
port 8 nsew default tristate
rlabel metal3 s 27303 10654 27735 10954 6 clockd[0]
port 9 nsew default tristate
rlabel metal3 s 27303 13646 27735 13946 6 div[4]
port 10 nsew default input
rlabel metal2 s 2216 27315 2356 27735 6 div[3]
port 11 nsew default input
rlabel metal3 s 0 15006 432 15306 4 div[2]
port 12 nsew default input
rlabel metal2 s 26504 0 26644 420 8 div[1]
port 13 nsew default input
rlabel metal2 s 4240 27315 4380 27735 6 div[0]
port 14 nsew default input
rlabel metal2 s 20432 0 20572 420 8 sel[2]
port 15 nsew default input
rlabel metal2 s 18408 0 18548 420 8 sel[1]
port 16 nsew default input
rlabel metal3 s 27303 1950 27735 2250 6 sel[0]
port 17 nsew default input
rlabel metal2 s 8288 0 8428 420 8 dco
port 18 nsew default input
rlabel metal3 s 0 9022 432 9322 4 ext_trim[25]
port 19 nsew default input
rlabel metal2 s 22456 0 22596 420 8 ext_trim[24]
port 20 nsew default input
rlabel metal3 s 27303 19630 27735 19930 6 ext_trim[23]
port 21 nsew default input
rlabel metal3 s 0 12014 432 12314 4 ext_trim[22]
port 22 nsew default input
rlabel metal3 s 0 26974 432 27274 4 ext_trim[21]
port 23 nsew default input
rlabel metal2 s 2216 0 2356 420 8 ext_trim[20]
port 24 nsew default input
rlabel metal2 s 4240 0 4380 420 8 ext_trim[19]
port 25 nsew default input
rlabel metal2 s 14360 0 14500 420 8 ext_trim[18]
port 26 nsew default input
rlabel metal2 s 10312 0 10452 420 8 ext_trim[17]
port 27 nsew default input
rlabel metal2 s 26320 27315 26460 27735 6 ext_trim[16]
port 28 nsew default input
rlabel metal2 s 12336 0 12476 420 8 ext_trim[15]
port 29 nsew default input
rlabel metal2 s 8288 27315 8428 27735 6 ext_trim[14]
port 30 nsew default input
rlabel metal2 s 14176 27315 14316 27735 6 ext_trim[13]
port 31 nsew default input
rlabel metal3 s 0 17998 432 18298 4 ext_trim[12]
port 32 nsew default input
rlabel metal2 s 6264 0 6404 420 8 ext_trim[11]
port 33 nsew default input
rlabel metal2 s 24296 27315 24436 27735 6 ext_trim[10]
port 34 nsew default input
rlabel metal2 s 12152 27315 12292 27735 6 ext_trim[9]
port 35 nsew default input
rlabel metal3 s 0 20990 432 21290 4 ext_trim[8]
port 36 nsew default input
rlabel metal3 s 0 6030 432 6330 4 ext_trim[7]
port 37 nsew default input
rlabel metal2 s 22272 27315 22412 27735 6 ext_trim[6]
port 38 nsew default input
rlabel metal2 s 20248 27315 20388 27735 6 ext_trim[5]
port 39 nsew default input
rlabel metal2 s 18224 27315 18364 27735 6 ext_trim[4]
port 40 nsew default input
rlabel metal3 s 27303 4942 27735 5242 6 ext_trim[3]
port 41 nsew default input
rlabel metal2 s 16200 27315 16340 27735 6 ext_trim[2]
port 42 nsew default input
rlabel metal3 s 27303 7662 27735 7962 6 ext_trim[1]
port 43 nsew default input
rlabel metal2 s 10312 27315 10452 27735 6 ext_trim[0]
port 44 nsew default input
flabel metal4 s 3526 464 3804 714 0 FreeSans 1600 0 0 0 vdd
port 45 nsew
flabel metal4 s 18884 474 19162 724 0 FreeSans 1600 0 0 0 vss
port 46 nsew
<< properties >>
string FIXED_BBOX 0 0 27735 27735
<< end >>
