magic
tech sky130A
magscale 1 2
timestamp 1587660775
<< checkpaint >>
rect -1260 -1260 887260 990260
<< viali >>
rect 342277 667569 342311 667603
rect 341081 667399 341115 667433
rect 228197 667297 228231 667331
rect 248437 667297 248471 667331
rect 268769 667297 268803 667331
rect 639529 280717 639563 280751
<< obsli1 >>
rect 519318 259446 519378 259454
<< metal1 >>
rect 351820 729372 351826 729424
rect 351878 729412 351884 729424
rect 353854 729412 353860 729424
rect 351878 729384 353860 729412
rect 351878 729372 351884 729384
rect 353854 729372 353860 729384
rect 353912 729412 353918 729424
rect 355914 729412 355920 729424
rect 353912 729384 355920 729412
rect 353912 729372 353918 729384
rect 355914 729372 355920 729384
rect 355972 729412 355978 729424
rect 356744 729412 356750 729424
rect 355972 729384 356750 729412
rect 355972 729372 355978 729384
rect 356744 729372 356750 729384
rect 356802 729372 356808 729424
rect 361030 729372 361036 729424
rect 361088 729412 361094 729424
rect 363098 729412 363126 729514
rect 366116 729412 366122 729424
rect 361088 729384 366122 729412
rect 361088 729372 361094 729384
rect 366116 729372 366122 729384
rect 366174 729372 366180 729424
rect 379016 729372 379022 729424
rect 379074 729412 379080 729424
rect 381056 729412 381062 729424
rect 379074 729384 381062 729412
rect 379074 729372 379080 729384
rect 381056 729372 381062 729384
rect 381114 729412 381120 729424
rect 383114 729412 383120 729424
rect 381114 729384 383120 729412
rect 381114 729372 381120 729384
rect 383114 729372 383120 729384
rect 383172 729412 383178 729424
rect 383944 729412 383950 729424
rect 383172 729384 383950 729412
rect 383172 729372 383178 729384
rect 383944 729372 383950 729384
rect 384002 729412 384008 729424
rect 386974 729412 386980 729424
rect 384002 729384 386980 729412
rect 384002 729372 384008 729384
rect 386974 729372 386980 729384
rect 387032 729412 387038 729424
rect 390304 729412 390332 729514
rect 393322 729412 393328 729424
rect 387032 729384 393328 729412
rect 387032 729372 387038 729384
rect 393322 729372 393328 729384
rect 393380 729372 393386 729424
rect 406386 729372 406392 729424
rect 406444 729412 406450 729424
rect 408042 729412 408048 729424
rect 406444 729384 408048 729412
rect 406444 729372 406450 729384
rect 408042 729372 408048 729384
rect 408100 729412 408106 729424
rect 410112 729412 410118 729424
rect 408100 729384 410118 729412
rect 408100 729372 408106 729384
rect 410112 729372 410118 729384
rect 410170 729372 410176 729424
rect 414298 729372 414304 729424
rect 414356 729412 414362 729424
rect 417306 729412 417334 729514
rect 420278 729412 420284 729424
rect 414356 729384 420284 729412
rect 414356 729372 414362 729384
rect 420278 729372 420284 729384
rect 420336 729372 420342 729424
rect 433220 729372 433226 729424
rect 433278 729412 433284 729424
rect 435256 729412 435262 729424
rect 433278 729384 435262 729412
rect 433278 729372 433284 729384
rect 435256 729372 435262 729384
rect 435314 729412 435320 729424
rect 437314 729412 437320 729424
rect 435314 729384 437320 729412
rect 435314 729372 435320 729384
rect 437314 729372 437320 729384
rect 437372 729412 437378 729424
rect 438144 729412 438150 729424
rect 437372 729384 438150 729412
rect 437372 729372 437378 729384
rect 438144 729372 438150 729384
rect 438202 729372 438208 729424
rect 441254 729372 441260 729424
rect 441312 729412 441318 729424
rect 444498 729412 444526 729514
rect 447510 729412 447516 729424
rect 441312 729384 447516 729412
rect 441312 729372 441318 729384
rect 447510 729372 447516 729384
rect 447568 729372 447574 729424
rect 460420 729372 460426 729424
rect 460478 729412 460484 729424
rect 462460 729412 462466 729424
rect 460478 729384 462466 729412
rect 460478 729372 460484 729384
rect 462460 729372 462466 729384
rect 462518 729412 462524 729424
rect 464514 729412 464520 729424
rect 462518 729384 464520 729412
rect 462518 729372 462524 729384
rect 464514 729372 464520 729384
rect 464572 729412 464578 729424
rect 465358 729412 465364 729424
rect 464572 729384 465364 729412
rect 464572 729372 464578 729384
rect 465358 729372 465364 729384
rect 465416 729412 465422 729424
rect 468578 729412 468584 729424
rect 465416 729384 468584 729412
rect 465416 729372 465422 729384
rect 468578 729372 468584 729384
rect 468636 729412 468642 729424
rect 471698 729412 471726 729514
rect 474742 729412 474748 729424
rect 468636 729384 474748 729412
rect 468636 729372 468642 729384
rect 474742 729372 474748 729384
rect 474800 729372 474806 729424
rect 487346 729372 487352 729424
rect 487404 729412 487410 729424
rect 489456 729412 489462 729424
rect 487404 729384 489462 729412
rect 487404 729372 487410 729384
rect 489456 729372 489462 729384
rect 489514 729412 489520 729424
rect 491514 729412 491520 729424
rect 489514 729384 491520 729412
rect 489514 729372 489520 729384
rect 491514 729372 491520 729384
rect 491572 729412 491578 729424
rect 492344 729412 492350 729424
rect 491572 729384 492350 729412
rect 491572 729372 491578 729384
rect 492344 729372 492350 729384
rect 492402 729412 492408 729424
rect 495442 729412 495448 729424
rect 492402 729384 495448 729412
rect 492402 729372 492408 729384
rect 495442 729372 495448 729384
rect 495500 729412 495506 729424
rect 498698 729412 498726 729514
rect 501716 729412 501722 729424
rect 495500 729384 501722 729412
rect 495500 729372 495506 729384
rect 501716 729372 501722 729384
rect 501774 729372 501780 729424
rect 514620 729372 514626 729424
rect 514678 729412 514684 729424
rect 516656 729412 516662 729424
rect 514678 729384 516662 729412
rect 514678 729372 514684 729384
rect 516656 729372 516662 729384
rect 516714 729412 516720 729424
rect 518718 729412 518724 729424
rect 516714 729384 518724 729412
rect 516714 729372 516720 729384
rect 518718 729372 518724 729384
rect 518776 729412 518782 729424
rect 519546 729412 519552 729424
rect 518776 729384 519552 729412
rect 518776 729372 518782 729384
rect 519546 729372 519552 729384
rect 519604 729412 519610 729424
rect 522674 729412 522680 729424
rect 519604 729384 522680 729412
rect 519604 729372 519610 729384
rect 522674 729372 522680 729384
rect 522732 729412 522738 729424
rect 525912 729412 525940 729514
rect 553098 729424 553126 729514
rect 575022 729480 575028 729492
rect 573154 729452 575028 729480
rect 528930 729412 528936 729424
rect 522732 729384 528936 729412
rect 522732 729372 522738 729384
rect 528930 729372 528936 729384
rect 528988 729372 528994 729424
rect 541902 729372 541908 729424
rect 541960 729412 541966 729424
rect 543856 729412 543862 729424
rect 541960 729384 543862 729412
rect 541960 729372 541966 729384
rect 543856 729372 543862 729384
rect 543914 729412 543920 729424
rect 545904 729412 545910 729424
rect 543914 729384 545910 729412
rect 543914 729372 543920 729384
rect 545904 729372 545910 729384
rect 545962 729412 545968 729424
rect 546732 729412 546738 729424
rect 545962 729384 546738 729412
rect 545962 729372 545968 729384
rect 546732 729372 546738 729384
rect 546790 729372 546796 729424
rect 553034 729372 553040 729424
rect 553092 729412 553126 729424
rect 556116 729412 556122 729424
rect 553092 729384 556122 729412
rect 553092 729372 553098 729384
rect 556116 729372 556122 729384
rect 556174 729372 556180 729424
rect 570330 729372 570336 729424
rect 570388 729412 570394 729424
rect 573154 729412 573182 729452
rect 575022 729440 575028 729452
rect 575080 729440 575086 729492
rect 570388 729384 573182 729412
rect 570388 729372 570394 729384
rect 573504 729372 573510 729424
rect 573562 729412 573568 729424
rect 573944 729412 573950 729424
rect 573562 729384 573950 729412
rect 573562 729372 573568 729384
rect 573944 729372 573950 729384
rect 574002 729412 574008 729424
rect 577046 729412 577052 729424
rect 574002 729384 577052 729412
rect 574002 729372 574008 729384
rect 577046 729372 577052 729384
rect 577104 729412 577110 729424
rect 580298 729412 580326 729514
rect 581161 729412 581167 729424
rect 577104 729384 581167 729412
rect 577104 729372 577110 729384
rect 581161 729372 581167 729384
rect 581219 729412 581225 729424
rect 583302 729412 583308 729424
rect 581219 729384 583308 729412
rect 581219 729372 581225 729384
rect 583302 729372 583308 729384
rect 583360 729372 583366 729424
rect 594158 729372 594164 729424
rect 594216 729412 594222 729424
rect 595875 729412 595881 729424
rect 594216 729384 595881 729412
rect 594216 729372 594222 729384
rect 595875 729372 595881 729384
rect 595933 729412 595939 729424
rect 595933 729384 596366 729412
rect 595933 729372 595939 729384
rect 380350 729304 380356 729356
rect 380408 729344 380414 729356
rect 384858 729344 384864 729356
rect 380408 729316 384864 729344
rect 380408 729304 380414 729316
rect 384858 729304 384864 729316
rect 384916 729304 384922 729356
rect 434545 729304 434551 729356
rect 434603 729344 434609 729356
rect 439138 729344 439144 729356
rect 434603 729316 439144 729344
rect 434603 729304 434609 729316
rect 439138 729304 439144 729316
rect 439196 729304 439202 729356
rect 488745 729304 488751 729356
rect 488803 729344 488809 729356
rect 493418 729344 493424 729356
rect 488803 729316 493424 729344
rect 488803 729304 488809 729316
rect 493418 729304 493424 729316
rect 493476 729304 493482 729356
rect 515958 729304 515964 729356
rect 516016 729344 516022 729356
rect 520466 729344 520472 729356
rect 516016 729316 520472 729344
rect 516016 729304 516022 729316
rect 520466 729304 520472 729316
rect 520524 729304 520530 729356
rect 522582 729304 522588 729356
rect 522640 729344 522646 729356
rect 523364 729344 523370 729356
rect 522640 729316 523370 729344
rect 522640 729304 522646 729316
rect 523364 729304 523370 729316
rect 523422 729304 523428 729356
rect 526761 729344 526767 729356
rect 523474 729316 526767 729344
rect 352382 729236 352388 729288
rect 352440 729276 352446 729288
rect 353145 729276 353151 729288
rect 352440 729248 353151 729276
rect 352440 729236 352446 729248
rect 353145 729236 353151 729248
rect 353203 729236 353209 729288
rect 431870 729236 431876 729288
rect 431928 729276 431934 729288
rect 432666 729276 432672 729288
rect 431928 729248 432672 729276
rect 431928 729236 431934 729248
rect 432666 729236 432672 729248
rect 432724 729236 432730 729288
rect 516878 729236 516884 729288
rect 516936 729276 516942 729288
rect 517865 729276 517871 729288
rect 516936 729248 517871 729276
rect 516936 729236 516942 729248
rect 517865 729236 517871 729248
rect 517923 729236 517929 729288
rect 519178 729236 519184 729288
rect 519236 729276 519242 729288
rect 523474 729276 523502 729316
rect 526761 729304 526767 729316
rect 526819 729304 526825 729356
rect 543145 729304 543151 729356
rect 543203 729344 543209 729356
rect 547698 729344 547704 729356
rect 543203 729316 547704 729344
rect 543203 729304 543209 729316
rect 547698 729304 547704 729316
rect 547756 729304 547762 729356
rect 568950 729304 568956 729356
rect 569008 729344 569014 729356
rect 571056 729344 571062 729356
rect 569008 729316 571062 729344
rect 569008 729304 569014 729316
rect 571056 729304 571062 729316
rect 571114 729344 571120 729356
rect 572262 729344 572268 729356
rect 571114 729316 572268 729344
rect 571114 729304 571120 729316
rect 572262 729304 572268 729316
rect 572320 729344 572326 729356
rect 573114 729344 573120 729356
rect 572320 729316 573120 729344
rect 572320 729304 572326 729316
rect 573114 729304 573120 729316
rect 573172 729304 573178 729356
rect 596338 729344 596366 729384
rect 597345 729372 597351 729424
rect 597403 729412 597409 729424
rect 601886 729412 601892 729424
rect 597403 729384 601892 729412
rect 597403 729372 597409 729384
rect 601886 729372 601892 729384
rect 601944 729372 601950 729424
rect 604765 729372 604771 729424
rect 604823 729412 604829 729424
rect 607298 729412 607326 729514
rect 624426 729430 624432 729482
rect 624484 729480 624490 729482
rect 629210 729480 629216 729492
rect 624484 729452 629216 729480
rect 624484 729430 624490 729452
rect 629210 729440 629216 729452
rect 629268 729440 629274 729492
rect 610442 729412 610448 729424
rect 604823 729384 610448 729412
rect 604823 729372 604829 729384
rect 610442 729372 610448 729384
rect 610500 729372 610506 729424
rect 623220 729372 623226 729424
rect 623278 729412 623284 729424
rect 625256 729412 625262 729424
rect 623278 729402 624137 729412
rect 624991 729402 625262 729412
rect 623278 729384 625262 729402
rect 623278 729372 623284 729384
rect 624095 729374 625027 729384
rect 625256 729372 625262 729384
rect 625314 729412 625320 729424
rect 626465 729412 626471 729424
rect 625314 729384 626471 729412
rect 625314 729372 625320 729384
rect 626465 729372 626471 729384
rect 626523 729412 626529 729424
rect 627324 729412 627330 729424
rect 626523 729384 627330 729412
rect 626523 729372 626529 729384
rect 627324 729372 627330 729384
rect 627382 729412 627388 729424
rect 627692 729412 627698 729424
rect 627382 729384 627698 729412
rect 627382 729372 627388 729384
rect 627692 729372 627698 729384
rect 627750 729412 627756 729424
rect 628152 729412 628158 729424
rect 627750 729384 628158 729412
rect 627750 729372 627756 729384
rect 628152 729372 628158 729384
rect 628210 729412 628216 729424
rect 631234 729412 631240 729424
rect 628210 729384 631240 729412
rect 628210 729372 628216 729384
rect 631234 729372 631240 729384
rect 631292 729412 631298 729424
rect 634498 729412 634526 729514
rect 635374 729412 635380 729424
rect 631292 729384 635380 729412
rect 631292 729372 631298 729384
rect 635374 729372 635380 729384
rect 635432 729412 635438 729424
rect 637490 729412 637496 729424
rect 635432 729384 637496 729412
rect 635432 729372 635438 729384
rect 637490 729372 637496 729384
rect 637548 729372 637554 729424
rect 650186 729372 650192 729424
rect 650244 729412 650250 729424
rect 650416 729412 650422 729424
rect 650244 729384 650422 729412
rect 650244 729372 650250 729384
rect 650416 729372 650422 729384
rect 650474 729412 650480 729424
rect 652456 729412 652462 729424
rect 650474 729384 652462 729412
rect 650474 729372 650480 729384
rect 652456 729372 652462 729384
rect 652514 729372 652520 729424
rect 654878 729372 654884 729424
rect 654936 729412 654942 729424
rect 654936 729384 658190 729412
rect 654936 729372 654942 729384
rect 598056 729344 598062 729356
rect 596338 729316 598062 729344
rect 598056 729304 598062 729316
rect 598114 729344 598120 729356
rect 600114 729344 600120 729356
rect 598114 729316 600120 729344
rect 598114 729304 598120 729316
rect 600114 729304 600120 729316
rect 600172 729304 600178 729356
rect 600506 729304 600512 729356
rect 600564 729344 600570 729356
rect 603843 729344 603849 729356
rect 600564 729316 603849 729344
rect 600564 729304 600570 729316
rect 603843 729304 603849 729316
rect 603901 729344 603907 729356
rect 608161 729344 608167 729356
rect 603901 729316 608167 729344
rect 603901 729304 603907 729316
rect 608161 729304 608167 729316
rect 608219 729304 608225 729356
rect 651750 729304 651756 729356
rect 651808 729344 651814 729356
rect 656258 729344 656264 729356
rect 651808 729316 656264 729344
rect 651808 729304 651814 729316
rect 656258 729304 656264 729316
rect 656316 729304 656322 729356
rect 658162 729344 658190 729384
rect 659165 729372 659171 729424
rect 659223 729412 659229 729424
rect 661704 729412 661732 729514
rect 664722 729412 664728 729424
rect 659223 729384 664728 729412
rect 659223 729372 659229 729384
rect 664722 729372 664728 729384
rect 664780 729372 664786 729424
rect 662561 729344 662567 729356
rect 658162 729316 662567 729344
rect 662561 729304 662567 729316
rect 662619 729304 662625 729356
rect 519236 729248 523502 729276
rect 519236 729236 519242 729248
rect 598574 729236 598580 729288
rect 598632 729276 598638 729288
rect 599264 729276 599270 729288
rect 598632 729248 599270 729276
rect 598632 729236 598638 729248
rect 599264 729236 599270 729248
rect 599322 729236 599328 729288
rect 600132 729276 600160 729304
rect 600944 729276 600950 729288
rect 600132 729248 600950 729276
rect 600944 729236 600950 729248
rect 601002 729236 601008 729288
rect 553310 729100 553316 729152
rect 553368 729140 553374 729152
rect 553954 729140 553960 729152
rect 553368 729112 553960 729140
rect 553368 729100 553374 729112
rect 553954 729100 553960 729112
rect 554012 729100 554018 729152
rect 465542 729032 465548 729084
rect 465600 729072 465606 729084
rect 492682 729072 492688 729084
rect 465600 729044 492688 729072
rect 465600 729032 465606 729044
rect 492682 729032 492688 729044
rect 492740 729032 492746 729084
rect 529114 729032 529120 729084
rect 529172 729072 529178 729084
rect 554690 729072 554696 729084
rect 529172 729044 554696 729072
rect 529172 729032 529178 729044
rect 554690 729032 554696 729044
rect 554748 729032 554754 729084
rect 555518 729032 555524 729084
rect 555576 729072 555582 729084
rect 556530 729072 556536 729084
rect 555576 729044 556536 729072
rect 555576 729032 555582 729044
rect 556530 729032 556536 729044
rect 556588 729072 556594 729084
rect 557082 729072 557088 729084
rect 556588 729044 557088 729072
rect 556588 729032 556594 729044
rect 557082 729032 557088 729044
rect 557140 729032 557146 729084
rect 602530 729032 602536 729084
rect 602588 729072 602594 729084
rect 610718 729072 610724 729084
rect 602588 729044 610724 729072
rect 602588 729032 602594 729044
rect 610718 729032 610724 729044
rect 610776 729032 610782 729084
rect 250906 728964 250912 729016
rect 250964 729004 250970 729016
rect 463610 729004 463616 729016
rect 250964 728976 463616 729004
rect 250964 728964 250970 728976
rect 463610 728964 463616 728976
rect 463668 728964 463674 729016
rect 474926 728964 474932 729016
rect 474984 729004 474990 729016
rect 500410 729004 500416 729016
rect 474984 728976 500416 729004
rect 474984 728964 474990 728976
rect 500410 728964 500416 728976
rect 500468 728964 500474 729016
rect 522490 728964 522496 729016
rect 522548 729004 522554 729016
rect 619550 729004 619556 729016
rect 522548 728976 619556 729004
rect 522548 728964 522554 728976
rect 619550 728964 619556 728976
rect 619608 728964 619614 729016
rect 360938 728896 360944 728948
rect 360996 728936 361002 728948
rect 568858 728936 568864 728948
rect 360996 728908 568864 728936
rect 360996 728896 361002 728908
rect 568858 728896 568864 728908
rect 568916 728896 568922 728948
rect 576494 728896 576500 728948
rect 576552 728936 576558 728948
rect 631142 728936 631148 728948
rect 576552 728908 631148 728936
rect 576552 728896 576558 728908
rect 631142 728896 631148 728908
rect 631200 728896 631206 728948
rect 356338 728828 356344 728880
rect 356396 728868 356402 728880
rect 363422 728868 363428 728880
rect 356396 728840 363428 728868
rect 356396 728828 356402 728840
rect 363422 728828 363428 728840
rect 363480 728868 363486 728880
rect 363974 728868 363980 728880
rect 363480 728840 363980 728868
rect 363480 728828 363486 728840
rect 363974 728828 363980 728840
rect 364032 728828 364038 728880
rect 366090 728828 366096 728880
rect 366148 728868 366154 728880
rect 378878 728868 378884 728880
rect 366148 728840 378884 728868
rect 366148 728828 366154 728840
rect 378878 728828 378884 728840
rect 378936 728828 378942 728880
rect 393322 728828 393328 728880
rect 393380 728868 393386 728880
rect 405742 728868 405748 728880
rect 393380 728840 405748 728868
rect 393380 728828 393386 728840
rect 405742 728828 405748 728840
rect 405800 728828 405806 728880
rect 420278 728828 420284 728880
rect 420336 728868 420342 728880
rect 433066 728868 433072 728880
rect 420336 728840 433072 728868
rect 420336 728828 420342 728840
rect 433066 728828 433072 728840
rect 433124 728828 433130 728880
rect 447510 728828 447516 728880
rect 447568 728868 447574 728880
rect 460298 728868 460304 728880
rect 447568 728840 460304 728868
rect 447568 728828 447574 728840
rect 460298 728828 460304 728840
rect 460356 728828 460362 728880
rect 463978 728828 463984 728880
rect 464036 728868 464042 728880
rect 464898 728868 464904 728880
rect 464036 728840 464904 728868
rect 464036 728828 464042 728840
rect 464898 728828 464904 728840
rect 464956 728868 464962 728880
rect 472258 728868 472264 728880
rect 464956 728840 472264 728868
rect 464956 728828 464962 728840
rect 472258 728828 472264 728840
rect 472316 728828 472322 728880
rect 474742 728828 474748 728880
rect 474800 728868 474806 728880
rect 487346 728868 487352 728880
rect 474800 728840 487352 728868
rect 474800 728828 474806 728840
rect 487346 728828 487352 728840
rect 487404 728828 487410 728880
rect 501698 728828 501704 728880
rect 501756 728868 501762 728880
rect 514486 728868 514492 728880
rect 501756 728840 514492 728868
rect 501756 728828 501762 728840
rect 514486 728828 514492 728840
rect 514544 728828 514550 728880
rect 521386 728868 521392 728880
rect 519058 728840 521392 728868
rect 358178 728760 358184 728812
rect 358236 728800 358242 728812
rect 366458 728800 366464 728812
rect 358236 728772 366464 728800
rect 358236 728760 358242 728772
rect 366458 728760 366464 728772
rect 366516 728800 366522 728812
rect 385502 728800 385508 728812
rect 366516 728772 385508 728800
rect 366516 728760 366522 728772
rect 385502 728760 385508 728772
rect 385560 728800 385566 728812
rect 393598 728800 393604 728812
rect 385560 728772 393604 728800
rect 385560 728760 385566 728772
rect 393598 728760 393604 728772
rect 393656 728800 393662 728812
rect 412458 728800 412464 728812
rect 393656 728772 412464 728800
rect 393656 728760 393662 728772
rect 412458 728760 412464 728772
rect 412516 728800 412522 728812
rect 420738 728800 420744 728812
rect 412516 728772 420744 728800
rect 412516 728760 412522 728772
rect 420738 728760 420744 728772
rect 420796 728800 420802 728812
rect 439598 728800 439604 728812
rect 420796 728772 439604 728800
rect 420796 728760 420802 728772
rect 439598 728760 439604 728772
rect 439656 728800 439662 728812
rect 447786 728800 447792 728812
rect 439656 728772 447792 728800
rect 439656 728760 439662 728772
rect 447786 728760 447792 728772
rect 447844 728800 447850 728812
rect 466922 728800 466928 728812
rect 447844 728772 466928 728800
rect 447844 728760 447850 728772
rect 466922 728760 466928 728772
rect 466980 728800 466986 728812
rect 475202 728800 475208 728812
rect 466980 728772 475208 728800
rect 466980 728760 466986 728772
rect 475202 728760 475208 728772
rect 475260 728800 475266 728812
rect 493878 728800 493884 728812
rect 475260 728772 493884 728800
rect 475260 728760 475266 728772
rect 493878 728760 493884 728772
rect 493936 728800 493942 728812
rect 502158 728800 502164 728812
rect 493936 728772 502164 728800
rect 493936 728760 493942 728772
rect 502158 728760 502164 728772
rect 502216 728800 502222 728812
rect 519058 728800 519086 728840
rect 521386 728828 521392 728840
rect 521444 728868 521450 728880
rect 529298 728868 529304 728880
rect 521444 728840 529304 728868
rect 521444 728828 521450 728840
rect 529298 728828 529304 728840
rect 529356 728868 529362 728880
rect 548250 728868 548256 728880
rect 529356 728840 548256 728868
rect 529356 728828 529362 728840
rect 548250 728828 548256 728840
rect 548308 728868 548314 728880
rect 555518 728868 555524 728880
rect 548308 728840 555524 728868
rect 548308 728828 548314 728840
rect 555518 728828 555524 728840
rect 555576 728828 555582 728880
rect 556254 728828 556260 728880
rect 556312 728868 556318 728880
rect 568490 728868 568496 728880
rect 556312 728840 568496 728868
rect 556312 728828 556318 728840
rect 568490 728828 568496 728840
rect 568548 728868 568554 728880
rect 577414 728868 577420 728880
rect 568548 728840 577420 728868
rect 568548 728828 568554 728840
rect 577414 728828 577420 728840
rect 577472 728828 577478 728880
rect 583302 728828 583308 728880
rect 583360 728868 583366 728880
rect 594158 728868 594164 728880
rect 583360 728840 594164 728868
rect 583360 728828 583366 728840
rect 594158 728828 594164 728840
rect 594216 728828 594222 728880
rect 611454 728828 611460 728880
rect 611512 728868 611518 728880
rect 622678 728868 622684 728880
rect 611512 728840 622684 728868
rect 611512 728828 611518 728840
rect 622678 728828 622684 728840
rect 622736 728868 622742 728880
rect 631970 728868 631976 728880
rect 622736 728840 631976 728868
rect 622736 728828 622742 728840
rect 631970 728828 631976 728840
rect 632028 728828 632034 728880
rect 502216 728772 519086 728800
rect 502216 728760 502222 728772
rect 528930 728760 528936 728812
rect 528988 728800 528994 728812
rect 541350 728800 541356 728812
rect 528988 728772 541356 728800
rect 528988 728760 528994 728772
rect 541350 728760 541356 728772
rect 541408 728760 541414 728812
rect 547698 728760 547704 728812
rect 547756 728800 547762 728812
rect 570330 728800 570336 728812
rect 547756 728772 570336 728800
rect 547756 728760 547762 728772
rect 570330 728760 570336 728772
rect 570388 728760 570394 728812
rect 577598 728760 577604 728812
rect 577656 728800 577662 728812
rect 583578 728800 583584 728812
rect 577656 728772 583584 728800
rect 577656 728760 577662 728772
rect 583578 728760 583584 728772
rect 583636 728800 583642 728812
rect 600506 728800 600512 728812
rect 583636 728772 600512 728800
rect 583636 728760 583642 728772
rect 600506 728760 600512 728772
rect 600564 728760 600570 728812
rect 610442 728760 610448 728812
rect 610500 728800 610506 728812
rect 623046 728800 623052 728812
rect 610500 728772 623052 728800
rect 610500 728760 610506 728772
rect 623046 728760 623052 728772
rect 623104 728760 623110 728812
rect 637674 728760 637680 728812
rect 637732 728800 637738 728812
rect 654878 728800 654884 728812
rect 637732 728772 654884 728800
rect 637732 728760 637738 728772
rect 654878 728760 654884 728772
rect 654936 728760 654942 728812
rect 353118 728692 353124 728744
rect 353176 728732 353182 728744
rect 357626 728732 357632 728744
rect 353176 728704 357632 728732
rect 353176 728692 353182 728704
rect 357626 728692 357632 728704
rect 357684 728732 357690 728744
rect 380350 728732 380356 728744
rect 357684 728704 380356 728732
rect 357684 728692 357690 728704
rect 380350 728692 380356 728704
rect 380408 728692 380414 728744
rect 384858 728692 384864 728744
rect 384916 728732 384922 728744
rect 407030 728732 407036 728744
rect 384916 728704 407036 728732
rect 384916 728692 384922 728704
rect 407030 728692 407036 728704
rect 407088 728732 407094 728744
rect 411906 728732 411912 728744
rect 407088 728704 411912 728732
rect 407088 728692 407094 728704
rect 411906 728692 411912 728704
rect 411964 728732 411970 728744
rect 434538 728732 434544 728744
rect 411964 728704 434544 728732
rect 411964 728692 411970 728704
rect 434538 728692 434544 728704
rect 434596 728692 434602 728744
rect 439138 728692 439144 728744
rect 439196 728732 439202 728744
rect 461770 728732 461776 728744
rect 439196 728704 461776 728732
rect 439196 728692 439202 728704
rect 461770 728692 461776 728704
rect 461828 728732 461834 728744
rect 466278 728732 466284 728744
rect 461828 728704 466284 728732
rect 461828 728692 461834 728704
rect 466278 728692 466284 728704
rect 466336 728732 466342 728744
rect 488726 728732 488732 728744
rect 466336 728704 488732 728732
rect 466336 728692 466342 728704
rect 488726 728692 488732 728704
rect 488784 728692 488790 728744
rect 493418 728692 493424 728744
rect 493476 728732 493482 728744
rect 515958 728732 515964 728744
rect 493476 728704 515964 728732
rect 493476 728692 493482 728704
rect 515958 728692 515964 728704
rect 516016 728692 516022 728744
rect 520466 728692 520472 728744
rect 520524 728732 520530 728744
rect 543098 728732 543104 728744
rect 520524 728704 543104 728732
rect 520524 728692 520530 728704
rect 543098 728692 543104 728704
rect 543156 728692 543162 728744
rect 546962 728692 546968 728744
rect 547020 728732 547026 728744
rect 547020 728704 573182 728732
rect 547020 728692 547026 728704
rect 356982 728664 356988 728676
rect 356770 728636 356988 728664
rect 287706 728420 287712 728472
rect 287764 728460 287770 728472
rect 356770 728460 356798 728636
rect 356982 728624 356988 728636
rect 357040 728664 357046 728676
rect 384030 728664 384036 728676
rect 357040 728636 384036 728664
rect 357040 728624 357046 728636
rect 384030 728624 384036 728636
rect 384088 728664 384094 728676
rect 411170 728664 411176 728676
rect 384088 728636 411176 728664
rect 384088 728624 384094 728636
rect 411170 728624 411176 728636
rect 411228 728664 411234 728676
rect 438310 728664 438316 728676
rect 411228 728636 438316 728664
rect 411228 728624 411234 728636
rect 438310 728624 438316 728636
rect 438368 728664 438374 728676
rect 465542 728664 465548 728676
rect 438368 728636 465548 728664
rect 438368 728624 438374 728636
rect 465542 728624 465548 728636
rect 465600 728624 465606 728676
rect 500410 728624 500416 728676
rect 500468 728664 500474 728676
rect 501606 728664 501612 728676
rect 500468 728636 501612 728664
rect 500468 728624 500474 728636
rect 501606 728624 501612 728636
rect 501664 728664 501670 728676
rect 529114 728664 529120 728676
rect 501664 728636 529120 728664
rect 501664 728624 501670 728636
rect 529114 728624 529120 728636
rect 529172 728624 529178 728676
rect 556162 728624 556168 728676
rect 556220 728664 556226 728676
rect 568950 728664 568956 728676
rect 556220 728636 568956 728664
rect 556220 728624 556226 728636
rect 568950 728624 568956 728636
rect 569008 728624 569014 728676
rect 573154 728664 573182 728704
rect 574930 728692 574936 728744
rect 574988 728732 574994 728744
rect 597286 728732 597292 728744
rect 574988 728704 597292 728732
rect 574988 728692 574994 728704
rect 597286 728692 597292 728704
rect 597344 728692 597350 728744
rect 601886 728692 601892 728744
rect 601944 728732 601950 728744
rect 624518 728732 624524 728744
rect 601944 728704 624524 728732
rect 601944 728692 601950 728704
rect 624518 728692 624524 728704
rect 624576 728692 624582 728744
rect 628382 728732 628388 728744
rect 627250 728704 628388 728732
rect 574194 728664 574200 728676
rect 573154 728636 574200 728664
rect 574194 728624 574200 728636
rect 574252 728664 574258 728676
rect 601150 728664 601156 728676
rect 574252 728636 601156 728664
rect 574252 728624 574258 728636
rect 601150 728624 601156 728636
rect 601208 728664 601214 728676
rect 627250 728664 627278 728704
rect 628382 728692 628388 728704
rect 628440 728732 628446 728744
rect 655430 728732 655436 728744
rect 628440 728704 655436 728732
rect 628440 728692 628446 728704
rect 654896 728676 654924 728704
rect 655430 728692 655436 728704
rect 655488 728692 655494 728744
rect 601208 728636 627278 728664
rect 601208 728624 601214 728636
rect 637490 728624 637496 728676
rect 637548 728664 637554 728676
rect 649542 728664 649548 728676
rect 637548 728636 649548 728664
rect 637548 728624 637554 728636
rect 649542 728624 649548 728636
rect 649600 728624 649606 728676
rect 654878 728624 654884 728676
rect 654936 728624 654942 728676
rect 368022 728556 368028 728608
rect 368080 728596 368086 728608
rect 392218 728596 392224 728608
rect 368080 728568 392224 728596
rect 368080 728556 368086 728568
rect 392218 728556 392224 728568
rect 392276 728596 392282 728608
rect 420186 728596 420192 728608
rect 392276 728568 420192 728596
rect 392276 728556 392282 728568
rect 420186 728556 420192 728568
rect 420244 728596 420250 728608
rect 447694 728596 447700 728608
rect 420244 728568 447700 728596
rect 420244 728556 420250 728568
rect 447694 728556 447700 728568
rect 447752 728596 447758 728608
rect 474926 728596 474932 728608
rect 447752 728568 474932 728596
rect 447752 728556 447758 728568
rect 474926 728556 474932 728568
rect 474984 728556 474990 728608
rect 492682 728556 492688 728608
rect 492740 728596 492746 728608
rect 519638 728596 519644 728608
rect 492740 728568 519644 728596
rect 492740 728556 492746 728568
rect 519638 728556 519644 728568
rect 519696 728596 519702 728608
rect 546962 728596 546968 728608
rect 519696 728568 546968 728596
rect 519696 728556 519702 728568
rect 546962 728556 546968 728568
rect 547020 728556 547026 728608
rect 550458 728556 550464 728608
rect 550516 728596 550522 728608
rect 621758 728596 621764 728608
rect 550516 728568 621764 728596
rect 550516 728556 550522 728568
rect 621758 728556 621764 728568
rect 621816 728556 621822 728608
rect 664722 728556 664728 728608
rect 664780 728596 664786 728608
rect 675946 728596 675952 728608
rect 664780 728568 675952 728596
rect 664780 728556 664786 728568
rect 675946 728556 675952 728568
rect 676004 728556 676010 728608
rect 468302 728488 468308 728540
rect 468360 728528 468366 728540
rect 468360 728500 511358 728528
rect 468360 728488 468366 728500
rect 287764 728432 356798 728460
rect 287764 728420 287770 728432
rect 383386 728420 383392 728472
rect 383444 728460 383450 728472
rect 391114 728460 391120 728472
rect 383444 728432 391120 728460
rect 383444 728420 383450 728432
rect 391114 728420 391120 728432
rect 391172 728420 391178 728472
rect 410710 728420 410716 728472
rect 410768 728460 410774 728472
rect 417518 728460 417524 728472
rect 410768 728432 417524 728460
rect 410768 728420 410774 728432
rect 417518 728420 417524 728432
rect 417576 728460 417582 728472
rect 418162 728460 418168 728472
rect 417576 728432 418168 728460
rect 417576 728420 417582 728432
rect 418162 728420 418168 728432
rect 418220 728420 418226 728472
rect 437482 728420 437488 728472
rect 437540 728460 437546 728472
rect 445302 728460 445308 728472
rect 437540 728432 445308 728460
rect 437540 728420 437546 728432
rect 445302 728420 445308 728432
rect 445360 728420 445366 728472
rect 491946 728420 491952 728472
rect 492004 728460 492010 728472
rect 499582 728460 499588 728472
rect 492004 728432 499588 728460
rect 492004 728420 492010 728432
rect 499582 728420 499588 728432
rect 499640 728420 499646 728472
rect 511330 728392 511358 728500
rect 629394 728488 629400 728540
rect 629452 728528 629458 728540
rect 651750 728528 651756 728540
rect 629452 728500 651756 728528
rect 629452 728488 629458 728500
rect 651750 728488 651756 728500
rect 651808 728488 651814 728540
rect 546318 728420 546324 728472
rect 546376 728460 546382 728472
rect 553310 728460 553316 728472
rect 546376 728432 553316 728460
rect 546376 728420 546382 728432
rect 553310 728420 553316 728432
rect 553368 728420 553374 728472
rect 575850 728420 575856 728472
rect 575908 728460 575914 728472
rect 583670 728460 583676 728472
rect 575908 728432 583676 728460
rect 575908 728420 575914 728432
rect 583670 728420 583676 728432
rect 583728 728420 583734 728472
rect 656258 728420 656264 728472
rect 656316 728460 656322 728472
rect 675854 728460 675860 728472
rect 656316 728432 675860 728460
rect 656316 728420 656322 728432
rect 675854 728420 675860 728432
rect 675912 728420 675918 728472
rect 597930 728392 597936 728404
rect 511330 728364 597936 728392
rect 597930 728352 597936 728364
rect 597988 728352 597994 728404
rect 335822 728284 335828 728336
rect 335880 728324 335886 728336
rect 441990 728324 441996 728336
rect 335880 728296 441996 728324
rect 335880 728284 335886 728296
rect 441990 728284 441996 728296
rect 442048 728284 442054 728336
rect 476398 728284 476404 728336
rect 476456 728324 476462 728336
rect 610074 728324 610080 728336
rect 476456 728296 610080 728324
rect 476456 728284 476462 728296
rect 610074 728284 610080 728296
rect 610132 728284 610138 728336
rect 436378 728216 436384 728268
rect 436436 728256 436442 728268
rect 600138 728256 600144 728268
rect 436436 728228 600144 728256
rect 436436 728216 436442 728228
rect 600138 728216 600144 728228
rect 600196 728216 600202 728268
rect 658248 728246 658300 728252
rect 414666 728148 414672 728200
rect 414724 728188 414730 728200
rect 584682 728188 584688 728200
rect 414724 728160 584688 728188
rect 414724 728148 414730 728160
rect 584682 728148 584688 728160
rect 584740 728148 584746 728200
rect 673124 728244 673176 728250
rect 658300 728205 673124 728233
rect 658248 728188 658300 728194
rect 673124 728185 673176 728192
rect 409238 728080 409244 728132
rect 409296 728120 409302 728132
rect 600230 728120 600236 728132
rect 409296 728092 600236 728120
rect 409296 728080 409302 728092
rect 600230 728080 600236 728092
rect 600288 728080 600294 728132
rect 394518 728012 394524 728064
rect 394576 728052 394582 728064
rect 589098 728052 589104 728064
rect 394576 728024 589104 728052
rect 394576 728012 394582 728024
rect 589098 728012 589104 728024
rect 589156 728012 589162 728064
rect 388078 727944 388084 727996
rect 388136 727984 388142 727996
rect 600322 727984 600328 727996
rect 388136 727956 600328 727984
rect 388136 727944 388142 727956
rect 600322 727944 600328 727956
rect 600380 727944 600386 727996
rect 378786 727876 378792 727928
rect 378844 727916 378850 727928
rect 593514 727916 593520 727928
rect 378844 727888 593520 727916
rect 378844 727876 378850 727888
rect 593514 727876 593520 727888
rect 593572 727876 593578 727928
rect 367654 727808 367660 727860
rect 367712 727848 367718 727860
rect 585602 727848 585608 727860
rect 367712 727820 585608 727848
rect 367712 727808 367718 727820
rect 585602 727808 585608 727820
rect 585660 727808 585666 727860
rect 499582 726856 499588 726908
rect 499640 726896 499646 726908
rect 594618 726896 594624 726908
rect 499640 726868 594624 726896
rect 499640 726856 499646 726868
rect 594618 726856 594624 726868
rect 594676 726856 594682 726908
rect 491026 726788 491032 726840
rect 491084 726828 491090 726840
rect 596826 726828 596832 726840
rect 491084 726800 596832 726828
rect 491084 726788 491090 726800
rect 596826 726788 596832 726800
rect 596884 726788 596890 726840
rect 382282 726720 382288 726772
rect 382340 726760 382346 726772
rect 569870 726760 569876 726772
rect 382340 726732 569876 726760
rect 382340 726720 382346 726732
rect 569870 726720 569876 726732
rect 569928 726720 569934 726772
rect 584682 726720 584688 726772
rect 584740 726760 584746 726772
rect 595722 726760 595728 726772
rect 584740 726732 595728 726760
rect 584740 726720 584746 726732
rect 595722 726720 595728 726732
rect 595780 726720 595786 726772
rect 568858 725700 568864 725752
rect 568916 725740 568922 725752
rect 583578 725740 583584 725752
rect 568916 725712 583584 725740
rect 568916 725700 568922 725712
rect 583578 725700 583584 725712
rect 583636 725700 583642 725752
rect 246306 725632 246312 725684
rect 246364 725672 246370 725684
rect 578426 725672 578432 725684
rect 246364 725644 578432 725672
rect 246364 725632 246370 725644
rect 578426 725632 578432 725644
rect 578484 725632 578490 725684
rect 246811 725452 246817 725504
rect 246869 725492 246875 725504
rect 649298 725492 649350 725499
rect 246869 725479 246979 725492
rect 246869 725464 649298 725479
rect 246869 725452 246875 725464
rect 246934 725451 649298 725464
rect 649298 725433 649350 725440
rect 448062 724544 448068 724596
rect 448120 724584 448126 724596
rect 464530 724584 464536 724596
rect 448120 724556 464536 724584
rect 448120 724544 448126 724556
rect 464530 724544 464536 724556
rect 464588 724544 464594 724596
rect 583578 724136 583584 724188
rect 583636 724176 583642 724188
rect 587994 724176 588000 724188
rect 583636 724148 588000 724176
rect 583636 724136 583642 724148
rect 587994 724136 588000 724148
rect 588052 724136 588058 724188
rect 585602 723456 585608 723508
rect 585660 723496 585666 723508
rect 585660 723468 588638 723496
rect 585660 723456 585666 723468
rect 588610 723428 588638 723468
rect 594618 723456 594624 723508
rect 594676 723496 594682 723508
rect 607314 723496 607320 723508
rect 594676 723468 607320 723496
rect 594676 723456 594682 723468
rect 607314 723456 607320 723468
rect 607372 723456 607378 723508
rect 599034 723428 599040 723440
rect 588610 723400 599040 723428
rect 599034 723388 599040 723400
rect 599092 723388 599098 723440
rect 593514 722640 593520 722692
rect 593572 722680 593578 722692
rect 594710 722680 594716 722692
rect 593572 722652 594716 722680
rect 593572 722640 593578 722652
rect 594710 722640 594716 722652
rect 594768 722640 594774 722692
rect 468302 722300 468308 722352
rect 468360 722340 468366 722352
rect 468854 722340 468860 722352
rect 468360 722312 468860 722340
rect 468360 722300 468366 722312
rect 468854 722300 468860 722312
rect 468912 722300 468918 722352
rect 589098 722232 589104 722284
rect 589156 722272 589162 722284
rect 594618 722272 594624 722284
rect 589156 722244 594624 722272
rect 589156 722232 589162 722244
rect 594618 722232 594624 722244
rect 594676 722232 594682 722284
rect 600230 722096 600236 722148
rect 600288 722136 600294 722148
rect 602346 722136 602352 722148
rect 600288 722108 602352 722136
rect 600288 722096 600294 722108
rect 602346 722096 602352 722108
rect 602404 722096 602410 722148
rect 596826 721416 596832 721468
rect 596884 721456 596890 721468
rect 603726 721456 603732 721468
rect 596884 721428 603732 721456
rect 596884 721416 596890 721428
rect 603726 721416 603732 721428
rect 603784 721416 603790 721468
rect 600322 721280 600328 721332
rect 600380 721320 600386 721332
rect 604554 721320 604560 721332
rect 600380 721292 604560 721320
rect 600380 721280 600386 721292
rect 604554 721280 604560 721292
rect 604612 721280 604618 721332
rect 652670 721212 652676 721264
rect 652728 721252 652734 721264
rect 653406 721252 653412 721264
rect 652728 721224 653412 721252
rect 652728 721212 652734 721224
rect 653406 721212 653412 721224
rect 653464 721212 653470 721264
rect 595722 720600 595728 720652
rect 595780 720640 595786 720652
rect 596826 720640 596832 720652
rect 595780 720612 596832 720640
rect 595780 720600 595786 720612
rect 596826 720600 596832 720612
rect 596884 720600 596890 720652
rect 610074 720124 610080 720176
rect 610132 720164 610138 720176
rect 616698 720164 616704 720176
rect 610132 720136 616704 720164
rect 610132 720124 610138 720136
rect 616698 720124 616704 720136
rect 616756 720124 616762 720176
rect 607314 720056 607320 720108
rect 607372 720096 607378 720108
rect 613478 720096 613484 720108
rect 607372 720068 613484 720096
rect 607372 720056 607378 720068
rect 613478 720056 613484 720068
rect 613536 720056 613542 720108
rect 359006 719036 359012 719088
rect 359064 719076 359070 719088
rect 359742 719076 359748 719088
rect 359064 719048 359748 719076
rect 359064 719036 359070 719048
rect 359742 719036 359748 719048
rect 359800 719036 359806 719088
rect 363422 719036 363428 719088
rect 363480 719076 363486 719088
rect 575390 719076 575396 719088
rect 363480 719048 575396 719076
rect 363480 719036 363486 719048
rect 575390 719036 575396 719048
rect 575448 719036 575454 719088
rect 597930 719036 597936 719088
rect 597988 719076 597994 719088
rect 605842 719076 605848 719088
rect 597988 719048 605848 719076
rect 597988 719036 597994 719048
rect 605842 719036 605848 719048
rect 605900 719036 605906 719088
rect 485966 718832 485972 718884
rect 486024 718872 486030 718884
rect 486518 718872 486524 718884
rect 486024 718844 486524 718872
rect 486024 718832 486030 718844
rect 486518 718832 486524 718844
rect 486576 718832 486582 718884
rect 605842 717880 605848 717932
rect 605900 717920 605906 717932
rect 613386 717920 613392 717932
rect 605900 717892 613392 717920
rect 605900 717880 605906 717892
rect 613386 717880 613392 717892
rect 613444 717880 613450 717932
rect 603726 716792 603732 716844
rect 603784 716832 603790 716844
rect 608970 716832 608976 716844
rect 603784 716804 608976 716832
rect 603784 716792 603790 716804
rect 608970 716792 608976 716804
rect 609028 716792 609034 716844
rect 464530 715704 464536 715756
rect 464588 715744 464594 715756
rect 468762 715744 468768 715756
rect 464588 715716 468768 715744
rect 464588 715704 464594 715716
rect 468762 715704 468768 715716
rect 468820 715704 468826 715756
rect 208126 714616 208132 714668
rect 208184 714656 208190 714668
rect 209966 714656 209972 714668
rect 208184 714628 209972 714656
rect 208184 714616 208190 714628
rect 209966 714616 209972 714628
rect 210024 714656 210030 714668
rect 351370 714656 351376 714668
rect 210024 714628 351376 714656
rect 210024 714616 210030 714628
rect 351370 714616 351376 714628
rect 351428 714616 351434 714668
rect 596826 714480 596832 714532
rect 596884 714520 596890 714532
rect 597930 714520 597936 714532
rect 596884 714492 597936 714520
rect 596884 714480 596890 714492
rect 597930 714480 597936 714492
rect 597988 714480 597994 714532
rect 600138 713528 600144 713580
rect 600196 713568 600202 713580
rect 604830 713568 604836 713580
rect 600196 713540 604836 713568
rect 600196 713528 600202 713540
rect 604830 713528 604836 713540
rect 604888 713528 604894 713580
rect 613478 713528 613484 713580
rect 613536 713568 613542 713580
rect 614582 713568 614588 713580
rect 613536 713540 614588 713568
rect 613536 713528 613542 713540
rect 614582 713528 614588 713540
rect 614640 713528 614646 713580
rect 599034 713460 599040 713512
rect 599092 713500 599098 713512
rect 606762 713500 606768 713512
rect 599092 713472 606768 713500
rect 599092 713460 599098 713472
rect 606762 713460 606768 713472
rect 606820 713460 606826 713512
rect 602346 712712 602352 712764
rect 602404 712752 602410 712764
rect 604646 712752 604652 712764
rect 602404 712724 604652 712752
rect 602404 712712 602410 712724
rect 604646 712712 604652 712724
rect 604704 712712 604710 712764
rect 594710 712576 594716 712628
rect 594768 712616 594774 712628
rect 600138 712616 600144 712628
rect 594768 712588 600144 712616
rect 594768 712576 594774 712588
rect 600138 712576 600144 712588
rect 600196 712576 600202 712628
rect 208126 711284 208132 711336
rect 208184 711324 208190 711336
rect 365630 711324 365636 711336
rect 208184 711296 365636 711324
rect 208184 711284 208190 711296
rect 365630 711284 365636 711296
rect 365688 711284 365694 711336
rect 468762 711284 468768 711336
rect 468820 711324 468826 711336
rect 478698 711324 478704 711336
rect 468820 711296 478704 711324
rect 468820 711284 468826 711296
rect 478698 711284 478704 711296
rect 478756 711284 478762 711336
rect 587994 711284 588000 711336
rect 588052 711324 588058 711336
rect 604738 711324 604744 711336
rect 588052 711296 604744 711324
rect 588052 711284 588058 711296
rect 604738 711284 604744 711296
rect 604796 711284 604802 711336
rect 594618 710264 594624 710316
rect 594676 710304 594682 710316
rect 598022 710304 598028 710316
rect 594676 710276 598028 710304
rect 594676 710264 594682 710276
rect 598022 710264 598028 710276
rect 598080 710264 598086 710316
rect 600138 708292 600144 708344
rect 600196 708332 600202 708344
rect 602346 708332 602352 708344
rect 600196 708304 602352 708332
rect 600196 708292 600202 708304
rect 602346 708292 602352 708304
rect 602404 708292 602410 708344
rect 608970 708292 608976 708344
rect 609028 708332 609034 708344
rect 611178 708332 611184 708344
rect 609028 708304 611184 708332
rect 609028 708292 609034 708304
rect 611178 708292 611184 708304
rect 611236 708292 611242 708344
rect 320734 707952 320740 708004
rect 320792 707992 320798 708004
rect 595262 707992 595268 708004
rect 320792 707964 595268 707992
rect 320792 707952 320798 707964
rect 595262 707952 595268 707964
rect 595320 707952 595326 708004
rect 604738 707272 604744 707324
rect 604796 707312 604802 707324
rect 605842 707312 605848 707324
rect 604796 707284 605848 707312
rect 604796 707272 604802 707284
rect 605842 707272 605848 707284
rect 605900 707272 605906 707324
rect 606762 707000 606768 707052
rect 606820 707040 606826 707052
rect 608050 707040 608056 707052
rect 606820 707012 608056 707040
rect 606820 707000 606826 707012
rect 608050 707000 608056 707012
rect 608108 707000 608114 707052
rect 604646 706320 604652 706372
rect 604704 706360 604710 706372
rect 607866 706360 607872 706372
rect 604704 706332 607872 706360
rect 604704 706320 604710 706332
rect 607866 706320 607872 706332
rect 607924 706320 607930 706372
rect 351278 705776 351284 705828
rect 351336 705816 351342 705828
rect 512462 705816 512468 705828
rect 351336 705788 512468 705816
rect 351336 705776 351342 705788
rect 512462 705776 512468 705788
rect 512520 705776 512526 705828
rect 344654 704688 344660 704740
rect 344712 704728 344718 704740
rect 541258 704728 541264 704740
rect 344712 704700 541264 704728
rect 344712 704688 344718 704700
rect 541258 704688 541264 704700
rect 541316 704688 541322 704740
rect 257898 703668 257904 703720
rect 257956 703708 257962 703720
rect 354590 703708 354596 703720
rect 257956 703680 354596 703708
rect 257956 703668 257962 703680
rect 354590 703668 354596 703680
rect 354648 703668 354654 703720
rect 354682 703532 354688 703584
rect 354740 703572 354746 703584
rect 513566 703572 513572 703584
rect 354740 703544 513572 703572
rect 354740 703532 354746 703544
rect 513566 703532 513572 703544
rect 513624 703532 513630 703584
rect 675946 702512 675952 702564
rect 676004 702552 676010 702564
rect 676222 702552 676228 702564
rect 676004 702524 676228 702552
rect 676004 702512 676010 702524
rect 676222 702512 676228 702524
rect 676280 702512 676286 702564
rect 598022 702444 598028 702496
rect 598080 702484 598086 702496
rect 605658 702484 605664 702496
rect 598080 702456 605664 702484
rect 598080 702444 598086 702456
rect 605658 702444 605664 702456
rect 605716 702444 605722 702496
rect 646506 701968 646512 702020
rect 646564 702008 646570 702020
rect 676038 702008 676044 702020
rect 646564 701980 676044 702008
rect 646564 701968 646570 701980
rect 676038 701968 676044 701980
rect 676096 701968 676102 702020
rect 323034 701356 323040 701408
rect 323092 701396 323098 701408
rect 383386 701396 383392 701408
rect 323092 701368 383392 701396
rect 323092 701356 323098 701368
rect 383386 701356 383392 701368
rect 383444 701356 383450 701408
rect 675854 701084 675860 701136
rect 675912 701124 675918 701136
rect 676314 701124 676320 701136
rect 675912 701096 676320 701124
rect 675912 701084 675918 701096
rect 676314 701084 676320 701096
rect 676372 701084 676378 701136
rect 605842 701016 605848 701068
rect 605900 701056 605906 701068
rect 607958 701056 607964 701068
rect 605900 701028 607964 701056
rect 605900 701016 605906 701028
rect 607958 701016 607964 701028
rect 608016 701016 608022 701068
rect 604830 700472 604836 700524
rect 604888 700512 604894 700524
rect 610074 700512 610080 700524
rect 604888 700484 610080 700512
rect 604888 700472 604894 700484
rect 610074 700472 610080 700484
rect 610132 700472 610138 700524
rect 597930 700404 597936 700456
rect 597988 700444 597994 700456
rect 600138 700444 600144 700456
rect 597988 700416 600144 700444
rect 597988 700404 597994 700416
rect 600138 700404 600144 700416
rect 600196 700404 600202 700456
rect 605658 700336 605664 700388
rect 605716 700376 605722 700388
rect 611270 700376 611276 700388
rect 605716 700348 611276 700376
rect 605716 700336 605722 700348
rect 611270 700336 611276 700348
rect 611328 700336 611334 700388
rect 248974 700268 248980 700320
rect 249032 700308 249038 700320
rect 386606 700308 386612 700320
rect 249032 700280 386612 700308
rect 249032 700268 249038 700280
rect 386606 700268 386612 700280
rect 386664 700268 386670 700320
rect 614582 699996 614588 700048
rect 614640 700036 614646 700048
rect 615594 700036 615600 700048
rect 614640 700008 615600 700036
rect 614640 699996 614646 700008
rect 615594 699996 615600 700008
rect 615652 699996 615658 700048
rect 613386 699860 613392 699912
rect 613444 699900 613450 699912
rect 614490 699900 614496 699912
rect 613444 699872 614496 699900
rect 613444 699860 613450 699872
rect 614490 699860 614496 699872
rect 614548 699860 614554 699912
rect 321102 699792 321108 699844
rect 321160 699832 321166 699844
rect 358730 699832 358736 699844
rect 321160 699804 358736 699832
rect 321160 699792 321166 699804
rect 358730 699792 358736 699804
rect 358788 699792 358794 699844
rect 604554 699792 604560 699844
rect 604612 699832 604618 699844
rect 605658 699832 605664 699844
rect 604612 699804 605664 699832
rect 604612 699792 604618 699804
rect 605658 699792 605664 699804
rect 605716 699792 605722 699844
rect 288718 699724 288724 699776
rect 288776 699764 288782 699776
rect 384950 699764 384956 699776
rect 288776 699736 384956 699764
rect 288776 699724 288782 699736
rect 384950 699724 384956 699736
rect 385008 699724 385014 699776
rect 255690 699520 255696 699572
rect 255748 699560 255754 699572
rect 308130 699560 308136 699572
rect 255748 699532 308136 699560
rect 255748 699520 255754 699532
rect 308130 699520 308136 699532
rect 308188 699520 308194 699572
rect 287246 699452 287252 699504
rect 287304 699492 287310 699504
rect 299850 699492 299856 699504
rect 287304 699464 299856 699492
rect 287304 699452 287310 699464
rect 299850 699452 299856 699464
rect 299908 699452 299914 699504
rect 302610 699452 302616 699504
rect 302668 699492 302674 699504
rect 329658 699492 329664 699504
rect 302668 699464 329664 699492
rect 302668 699452 302674 699464
rect 329658 699452 329664 699464
rect 329716 699452 329722 699504
rect 250170 699384 250176 699436
rect 250228 699424 250234 699436
rect 301138 699424 301144 699436
rect 250228 699396 301144 699424
rect 250228 699384 250234 699396
rect 301138 699384 301144 699396
rect 301196 699384 301202 699436
rect 303898 699384 303904 699436
rect 303956 699424 303962 699436
rect 321562 699424 321568 699436
rect 303956 699396 321568 699424
rect 303956 699384 303962 699396
rect 321562 699384 321568 699396
rect 321620 699384 321626 699436
rect 210426 699316 210432 699368
rect 210484 699356 210490 699368
rect 309418 699356 309424 699368
rect 210484 699328 309424 699356
rect 210484 699316 210490 699328
rect 309418 699316 309424 699328
rect 309476 699316 309482 699368
rect 317698 699316 317704 699368
rect 317756 699356 317762 699368
rect 324782 699356 324788 699368
rect 317756 699328 324788 699356
rect 317756 699316 317762 699328
rect 324782 699316 324788 699328
rect 324840 699316 324846 699368
rect 288626 699248 288632 699300
rect 288684 699288 288690 699300
rect 330762 699288 330768 699300
rect 288684 699260 330768 699288
rect 288684 699248 288690 699260
rect 330762 699248 330768 699260
rect 330820 699248 330826 699300
rect 289086 699180 289092 699232
rect 289144 699220 289150 699232
rect 361766 699220 361772 699232
rect 289144 699192 361772 699220
rect 289144 699180 289150 699192
rect 361766 699180 361772 699192
rect 361824 699180 361830 699232
rect 249618 699112 249624 699164
rect 249676 699152 249682 699164
rect 292858 699152 292864 699164
rect 249676 699124 292864 699152
rect 249676 699112 249682 699124
rect 292858 699112 292864 699124
rect 292916 699152 292922 699164
rect 321838 699152 321844 699164
rect 292916 699124 321844 699152
rect 292916 699112 292922 699124
rect 321838 699112 321844 699124
rect 321896 699112 321902 699164
rect 249526 699044 249532 699096
rect 249584 699084 249590 699096
rect 295618 699084 295624 699096
rect 249584 699056 295624 699084
rect 249584 699044 249590 699056
rect 295618 699044 295624 699056
rect 295676 699044 295682 699096
rect 297274 699044 297280 699096
rect 297332 699084 297338 699096
rect 322022 699084 322028 699096
rect 297332 699056 322028 699084
rect 297332 699044 297338 699056
rect 322022 699044 322028 699056
rect 322080 699044 322086 699096
rect 294974 698976 294980 699028
rect 295032 699016 295038 699028
rect 301782 699016 301788 699028
rect 295032 698988 301788 699016
rect 295032 698976 295038 698988
rect 301782 698976 301788 698988
rect 301840 698976 301846 699028
rect 302536 698988 302840 699016
rect 249342 698908 249348 698960
rect 249400 698948 249406 698960
rect 302536 698948 302564 698988
rect 249400 698920 302564 698948
rect 302812 698948 302840 698988
rect 305554 698976 305560 699028
rect 305612 699016 305618 699028
rect 328554 699016 328560 699028
rect 305612 698988 328560 699016
rect 305612 698976 305618 698988
rect 328554 698976 328560 698988
rect 328612 698976 328618 699028
rect 306658 698948 306664 698960
rect 302812 698920 306664 698948
rect 249400 698908 249406 698920
rect 306658 698908 306664 698920
rect 306716 698908 306722 698960
rect 316594 698908 316600 698960
rect 316652 698948 316658 698960
rect 596826 698948 596832 698960
rect 316652 698920 596832 698948
rect 316652 698908 316658 698920
rect 596826 698908 596832 698920
rect 596884 698908 596890 698960
rect 250630 698840 250636 698892
rect 250688 698880 250694 698892
rect 301690 698880 301696 698892
rect 250688 698852 301696 698880
rect 250688 698840 250694 698852
rect 301690 698840 301696 698852
rect 301748 698840 301754 698892
rect 301782 698840 301788 698892
rect 301840 698840 301846 698892
rect 306842 698840 306848 698892
rect 306900 698880 306906 698892
rect 313650 698880 313656 698892
rect 306900 698852 313656 698880
rect 306900 698840 306906 698852
rect 313650 698840 313656 698852
rect 313708 698840 313714 698892
rect 314220 698852 318158 698880
rect 301800 698812 301828 698840
rect 314220 698812 314248 698852
rect 301800 698784 314248 698812
rect 318130 698812 318158 698852
rect 320642 698840 320648 698892
rect 320700 698880 320706 698892
rect 361674 698880 361680 698892
rect 320700 698852 361680 698880
rect 320700 698840 320706 698852
rect 361674 698840 361680 698852
rect 361732 698840 361738 698892
rect 474282 698812 474288 698824
rect 318130 698784 474288 698812
rect 474282 698772 474288 698784
rect 474340 698772 474346 698824
rect 251274 698704 251280 698756
rect 251332 698744 251338 698756
rect 314818 698744 314824 698754
rect 251332 698716 314824 698744
rect 251332 698704 251338 698716
rect 314818 698702 314824 698716
rect 314876 698702 314882 698754
rect 321194 698704 321200 698756
rect 321252 698744 321258 698756
rect 576954 698744 576960 698756
rect 321252 698716 576960 698744
rect 321252 698704 321258 698716
rect 576954 698704 576960 698716
rect 577012 698704 577018 698756
rect 676314 698744 676320 698756
rect 670306 698716 676320 698744
rect 654234 698636 654240 698688
rect 654292 698676 654298 698688
rect 670306 698676 670334 698716
rect 676314 698704 676320 698716
rect 676372 698704 676378 698756
rect 654292 698648 670334 698676
rect 654292 698636 654298 698648
rect 323678 698092 323684 698144
rect 323736 698132 323742 698144
rect 390010 698132 390016 698144
rect 323736 698104 390016 698132
rect 323736 698092 323742 698104
rect 390010 698092 390016 698104
rect 390068 698092 390074 698144
rect 321562 698024 321568 698076
rect 321620 698064 321626 698076
rect 508138 698064 508144 698076
rect 321620 698036 508144 698064
rect 321620 698024 321626 698036
rect 508138 698024 508144 698036
rect 508196 698024 508202 698076
rect 675946 697948 675952 698000
rect 676004 697988 676010 698000
rect 676320 697990 676326 698002
rect 676038 697988 676326 697990
rect 676004 697962 676326 697988
rect 676004 697960 676076 697962
rect 676004 697948 676010 697960
rect 676320 697950 676326 697962
rect 676378 697950 676384 698002
rect 675670 697480 675676 697532
rect 675728 697520 675734 697532
rect 676038 697520 676044 697532
rect 675728 697492 676044 697520
rect 675728 697480 675734 697492
rect 676038 697480 676044 697492
rect 676096 697480 676102 697532
rect 478698 696936 478704 696988
rect 478756 696976 478762 696988
rect 489738 696976 489744 696988
rect 478756 696948 489744 696976
rect 478756 696936 478762 696948
rect 489738 696936 489744 696948
rect 489796 696936 489802 696988
rect 664814 696936 664820 696988
rect 664872 696976 664878 696988
rect 667482 696976 667488 696988
rect 664872 696948 667488 696976
rect 664872 696936 664878 696948
rect 667482 696936 667488 696948
rect 667540 696936 667546 696988
rect 675578 696528 675584 696580
rect 675636 696568 675642 696580
rect 675854 696568 675860 696580
rect 675636 696540 675860 696568
rect 675636 696528 675642 696540
rect 675854 696528 675860 696540
rect 675912 696568 675918 696580
rect 676314 696568 676320 696580
rect 675912 696540 676320 696568
rect 675912 696528 675918 696540
rect 676314 696528 676320 696540
rect 676372 696528 676378 696580
rect 654878 696460 654884 696512
rect 654936 696500 654942 696512
rect 676038 696500 676044 696512
rect 654936 696472 676044 696500
rect 654936 696460 654942 696472
rect 676038 696460 676044 696472
rect 676096 696460 676102 696512
rect 675762 696052 675768 696104
rect 675820 696092 675826 696104
rect 676038 696092 676044 696104
rect 675820 696064 676044 696092
rect 675820 696052 675826 696064
rect 676038 696052 676044 696064
rect 676096 696052 676102 696104
rect 320550 695780 320556 695832
rect 320608 695820 320614 695832
rect 321194 695820 321200 695832
rect 320608 695792 321200 695820
rect 320608 695780 320614 695792
rect 321194 695780 321200 695792
rect 321252 695780 321258 695832
rect 557082 695372 557088 695424
rect 557140 695412 557146 695424
rect 675854 695412 675860 695424
rect 557140 695384 675860 695412
rect 557140 695372 557146 695384
rect 675854 695372 675860 695384
rect 675912 695412 675918 695424
rect 676038 695412 676044 695424
rect 675912 695384 676044 695412
rect 675912 695372 675918 695384
rect 676038 695372 676044 695384
rect 676096 695372 676102 695424
rect 384950 695304 384956 695356
rect 385008 695344 385014 695356
rect 387158 695344 387164 695356
rect 385008 695316 387164 695344
rect 385008 695304 385014 695316
rect 387158 695304 387164 695316
rect 387216 695344 387222 695356
rect 619642 695344 619648 695356
rect 387216 695316 619648 695344
rect 387216 695304 387222 695316
rect 619642 695304 619648 695316
rect 619700 695304 619706 695356
rect 320642 695100 320648 695152
rect 320700 695140 320706 695152
rect 322574 695140 322580 695152
rect 320700 695112 322580 695140
rect 320700 695100 320706 695112
rect 322574 695100 322580 695112
rect 322632 695100 322638 695152
rect 321930 694760 321936 694812
rect 321988 694800 321994 694812
rect 370782 694800 370788 694812
rect 321988 694772 370788 694800
rect 321988 694760 321994 694772
rect 370782 694760 370788 694772
rect 370840 694760 370846 694812
rect 361858 694692 361864 694744
rect 361916 694732 361922 694744
rect 376670 694732 376676 694744
rect 361916 694704 376676 694732
rect 361916 694692 361922 694704
rect 376670 694692 376676 694704
rect 376728 694692 376734 694744
rect 358730 694624 358736 694676
rect 358788 694664 358794 694676
rect 372806 694664 372812 694676
rect 358788 694636 372812 694664
rect 358788 694624 358794 694636
rect 372806 694624 372812 694636
rect 372864 694624 372870 694676
rect 381270 694624 381276 694676
rect 381328 694664 381334 694676
rect 460574 694664 460580 694676
rect 381328 694636 460580 694664
rect 381328 694624 381334 694636
rect 460574 694624 460580 694636
rect 460632 694624 460638 694676
rect 321838 694556 321844 694608
rect 321896 694596 321902 694608
rect 388814 694596 388820 694608
rect 321896 694568 388820 694596
rect 321896 694556 321902 694568
rect 388814 694556 388820 694568
rect 388872 694556 388878 694608
rect 321010 694488 321016 694540
rect 321068 694528 321074 694540
rect 375198 694528 375204 694540
rect 321068 694500 375204 694528
rect 321068 694488 321074 694500
rect 375198 694488 375204 694500
rect 375256 694528 375262 694540
rect 625070 694528 625076 694540
rect 375256 694500 625076 694528
rect 375256 694488 375262 694500
rect 625070 694488 625076 694500
rect 625128 694488 625134 694540
rect 675670 694488 675676 694540
rect 675728 694528 675734 694540
rect 676130 694528 676136 694540
rect 675728 694500 676136 694528
rect 675728 694488 675734 694500
rect 676130 694488 676136 694500
rect 676188 694488 676194 694540
rect 624426 694216 624432 694268
rect 624484 694256 624490 694268
rect 676038 694256 676044 694268
rect 624484 694228 676044 694256
rect 624484 694216 624490 694228
rect 676038 694216 676044 694228
rect 676096 694216 676102 694268
rect 675854 694012 675860 694064
rect 675912 694052 675918 694064
rect 676130 694052 676136 694064
rect 675912 694024 676136 694052
rect 675912 694012 675918 694024
rect 676130 694012 676136 694024
rect 676188 694012 676194 694064
rect 208126 693944 208132 693996
rect 208184 693984 208190 693996
rect 208310 693984 208316 693996
rect 208184 693956 208316 693984
rect 208184 693944 208190 693956
rect 208310 693944 208316 693956
rect 208368 693944 208374 693996
rect 324782 693128 324788 693180
rect 324840 693168 324846 693180
rect 356982 693168 356988 693180
rect 324840 693140 356988 693168
rect 324840 693128 324846 693140
rect 356982 693128 356988 693140
rect 357040 693128 357046 693180
rect 450730 693128 450736 693180
rect 450788 693168 450794 693180
rect 676314 693168 676320 693180
rect 450788 693140 676320 693168
rect 450788 693128 450794 693140
rect 676314 693128 676320 693140
rect 676372 693128 676378 693180
rect 226248 692698 226776 692716
rect 208126 692516 208132 692568
rect 208184 692556 208190 692568
rect 208954 692556 208960 692568
rect 208184 692528 208960 692556
rect 208184 692516 208190 692528
rect 208954 692516 208960 692528
rect 209012 692556 209018 692568
rect 226248 692556 226265 692698
rect 209012 692528 226265 692556
rect 209012 692516 209018 692528
rect 226248 692383 226265 692528
rect 226757 692556 226776 692698
rect 287706 692556 287712 692568
rect 226757 692528 287712 692556
rect 226757 692383 226776 692528
rect 287706 692516 287712 692528
rect 287764 692516 287770 692568
rect 226248 692366 226776 692383
rect 608050 692040 608056 692092
rect 608108 692080 608114 692092
rect 611454 692080 611460 692092
rect 608108 692052 611460 692080
rect 608108 692040 608114 692052
rect 611454 692040 611460 692052
rect 611512 692040 611518 692092
rect 320642 691428 320648 691480
rect 320700 691468 320706 691480
rect 321102 691468 321108 691480
rect 320700 691440 321108 691468
rect 320700 691428 320706 691440
rect 321102 691428 321108 691440
rect 321160 691428 321166 691480
rect 676222 691162 676228 691214
rect 676280 691202 676286 691214
rect 676280 691174 676437 691202
rect 676280 691162 676286 691174
rect 611178 690612 611184 690664
rect 611236 690652 611242 690664
rect 612282 690652 612288 690664
rect 611236 690624 612288 690652
rect 611236 690612 611242 690624
rect 612282 690612 612288 690624
rect 612340 690612 612346 690664
rect 675854 690272 675860 690324
rect 675912 690312 675918 690324
rect 676314 690312 676320 690324
rect 675912 690284 676320 690312
rect 675912 690272 675918 690284
rect 676314 690272 676320 690284
rect 676372 690272 676378 690324
rect 506298 689796 506304 689848
rect 506356 689836 506362 689848
rect 675854 689836 675860 689848
rect 506356 689808 675860 689836
rect 506356 689796 506362 689808
rect 675854 689796 675860 689808
rect 675912 689796 675918 689848
rect 576954 689184 576960 689236
rect 577012 689224 577018 689236
rect 590202 689224 590208 689236
rect 577012 689196 590208 689224
rect 577012 689184 577018 689196
rect 590202 689184 590208 689196
rect 590260 689184 590266 689236
rect 676038 688096 676044 688148
rect 676096 688136 676102 688148
rect 676314 688136 676320 688148
rect 676096 688108 676320 688136
rect 676096 688096 676102 688108
rect 676314 688096 676320 688108
rect 676372 688096 676378 688148
rect 251734 687620 251740 687672
rect 251792 687660 251798 687672
rect 279886 687660 279892 687672
rect 251792 687632 279892 687660
rect 251792 687620 251798 687632
rect 279886 687620 279892 687632
rect 279944 687620 279950 687672
rect 667482 687620 667488 687672
rect 667540 687660 667546 687672
rect 675946 687660 675952 687672
rect 667540 687632 675952 687660
rect 667540 687620 667546 687632
rect 675946 687620 675952 687632
rect 676004 687620 676010 687672
rect 675670 687076 675676 687128
rect 675728 687116 675734 687128
rect 676314 687116 676320 687128
rect 675728 687088 676320 687116
rect 675728 687076 675734 687088
rect 676314 687076 676320 687088
rect 676372 687076 676378 687128
rect 489738 687008 489744 687060
rect 489796 687048 489802 687060
rect 496362 687048 496368 687060
rect 489796 687020 496368 687048
rect 489796 687008 489802 687020
rect 496362 687008 496368 687020
rect 496420 687008 496426 687060
rect 675762 687008 675768 687060
rect 675820 687048 675826 687060
rect 676222 687048 676228 687060
rect 675820 687020 676228 687048
rect 675820 687008 675826 687020
rect 676222 687008 676228 687020
rect 676280 687008 676286 687060
rect 602346 684764 602352 684816
rect 602404 684804 602410 684816
rect 611178 684804 611184 684816
rect 602404 684776 611184 684804
rect 602404 684764 602410 684776
rect 611178 684764 611184 684776
rect 611236 684764 611242 684816
rect 614490 684560 614496 684612
rect 614548 684600 614554 684612
rect 615686 684600 615692 684612
rect 614548 684572 615692 684600
rect 614548 684560 614554 684572
rect 615686 684560 615692 684572
rect 615744 684560 615750 684612
rect 596826 684492 596832 684544
rect 596884 684532 596890 684544
rect 603542 684532 603548 684544
rect 596884 684504 603548 684532
rect 596884 684492 596890 684504
rect 603542 684492 603548 684504
rect 603600 684492 603606 684544
rect 322022 684288 322028 684340
rect 322080 684328 322086 684340
rect 360662 684328 360668 684340
rect 322080 684300 360668 684328
rect 322080 684288 322086 684300
rect 360662 684288 360668 684300
rect 360720 684288 360726 684340
rect 616698 684084 616704 684136
rect 616756 684124 616762 684136
rect 617894 684124 617900 684136
rect 616756 684096 617900 684124
rect 616756 684084 616762 684096
rect 617894 684084 617900 684096
rect 617952 684084 617958 684136
rect 600138 683064 600144 683116
rect 600196 683104 600202 683116
rect 603450 683104 603456 683116
rect 600196 683076 603456 683104
rect 600196 683064 600202 683076
rect 603450 683064 603456 683076
rect 603508 683064 603514 683116
rect 330762 682112 330768 682164
rect 330820 682152 330826 682164
rect 359834 682152 359840 682164
rect 330820 682124 359840 682152
rect 330820 682112 330826 682124
rect 359834 682112 359840 682124
rect 359892 682112 359898 682164
rect 496362 682112 496368 682164
rect 496420 682152 496426 682164
rect 506390 682152 506396 682164
rect 496420 682124 506396 682152
rect 496420 682112 496426 682124
rect 506390 682112 506396 682124
rect 506448 682112 506454 682164
rect 590202 681500 590208 681552
rect 590260 681540 590266 681552
rect 600138 681540 600144 681552
rect 590260 681512 600144 681540
rect 590260 681500 590266 681512
rect 600138 681500 600144 681512
rect 600196 681500 600202 681552
rect 607958 681432 607964 681484
rect 608016 681472 608022 681484
rect 612558 681472 612564 681484
rect 608016 681444 612564 681472
rect 608016 681432 608022 681444
rect 612558 681432 612564 681444
rect 612616 681432 612622 681484
rect 611270 681092 611276 681144
rect 611328 681132 611334 681144
rect 612466 681132 612472 681144
rect 611328 681104 612472 681132
rect 611328 681092 611334 681104
rect 612466 681092 612472 681104
rect 612524 681092 612530 681144
rect 611454 681024 611460 681076
rect 611512 681064 611518 681076
rect 614582 681064 614588 681076
rect 611512 681036 614588 681064
rect 611512 681024 611518 681036
rect 614582 681024 614588 681036
rect 614640 681024 614646 681076
rect 610074 680956 610080 681008
rect 610132 680996 610138 681008
rect 613386 680996 613392 681008
rect 610132 680968 613392 680996
rect 610132 680956 610138 680968
rect 613386 680956 613392 680968
rect 613444 680956 613450 681008
rect 650922 680956 650928 681008
rect 650980 680996 650986 681008
rect 654234 680996 654240 681008
rect 650980 680968 654240 680996
rect 650980 680956 650986 680968
rect 654234 680956 654240 680968
rect 654292 680956 654298 681008
rect 328554 678780 328560 678832
rect 328612 678820 328618 678832
rect 362594 678820 362600 678832
rect 328612 678792 362600 678820
rect 328612 678780 328618 678792
rect 362594 678780 362600 678792
rect 362652 678780 362658 678832
rect 612558 677760 612564 677812
rect 612616 677800 612622 677812
rect 614490 677800 614496 677812
rect 612616 677772 614496 677800
rect 612616 677760 612622 677772
rect 614490 677760 614496 677772
rect 614548 677760 614554 677812
rect 208126 677556 208132 677608
rect 208184 677596 208190 677608
rect 209966 677596 209972 677608
rect 208184 677568 209972 677596
rect 208184 677556 208190 677568
rect 209966 677556 209972 677568
rect 210024 677556 210030 677608
rect 390194 676604 390200 676656
rect 390252 676644 390258 676656
rect 390654 676644 390660 676656
rect 390252 676616 390660 676644
rect 390252 676604 390258 676616
rect 390654 676604 390660 676616
rect 390712 676604 390718 676656
rect 607866 676604 607872 676656
rect 607924 676644 607930 676656
rect 608970 676644 608976 676656
rect 607924 676616 608976 676644
rect 607924 676604 607930 676616
rect 608970 676604 608976 676616
rect 609028 676604 609034 676656
rect 605658 676468 605664 676520
rect 605716 676508 605722 676520
rect 606854 676508 606860 676520
rect 605716 676480 606860 676508
rect 605716 676468 605722 676480
rect 606854 676468 606860 676480
rect 606912 676468 606918 676520
rect 390194 676264 390200 676316
rect 390252 676304 390258 676316
rect 390378 676304 390384 676316
rect 390252 676276 390384 676304
rect 390252 676264 390258 676276
rect 390378 676264 390384 676276
rect 390436 676264 390442 676316
rect 614582 676264 614588 676316
rect 614640 676304 614646 676316
rect 616698 676304 616704 676316
rect 614640 676276 616704 676304
rect 614640 676264 614646 676276
rect 616698 676264 616704 676276
rect 616756 676264 616762 676316
rect 612466 676128 612472 676180
rect 612524 676168 612530 676180
rect 614582 676168 614588 676180
rect 612524 676140 614588 676168
rect 612524 676128 612530 676140
rect 614582 676128 614588 676140
rect 614640 676128 614646 676180
rect 643194 675924 643200 675976
rect 643252 675964 643258 675976
rect 650922 675964 650928 675976
rect 643252 675936 650928 675964
rect 643252 675924 643258 675936
rect 650922 675924 650928 675936
rect 650980 675924 650986 675976
rect 603542 674836 603548 674888
rect 603600 674876 603606 674888
rect 610810 674876 610816 674888
rect 603600 674848 610816 674876
rect 603600 674836 603606 674848
rect 610810 674836 610816 674848
rect 610868 674836 610874 674888
rect 248146 674360 248152 674412
rect 248204 674400 248210 674412
rect 287982 674400 287988 674412
rect 248204 674372 287988 674400
rect 248204 674360 248210 674372
rect 287982 674360 287988 674372
rect 288040 674360 288046 674412
rect 603450 673340 603456 673392
rect 603508 673380 603514 673392
rect 606762 673380 606768 673392
rect 603508 673352 606768 673380
rect 603508 673340 603514 673352
rect 606762 673340 606768 673352
rect 606820 673340 606826 673392
rect 329658 673272 329664 673324
rect 329716 673312 329722 673324
rect 360754 673312 360760 673324
rect 329716 673284 360760 673312
rect 329716 673272 329722 673284
rect 360754 673272 360760 673284
rect 360812 673272 360818 673324
rect 417518 671504 417524 671556
rect 417576 671544 417582 671556
rect 536750 671544 536756 671556
rect 417576 671516 536756 671544
rect 417576 671504 417582 671516
rect 536750 671504 536756 671516
rect 536808 671504 536814 671556
rect 600138 671504 600144 671556
rect 600196 671544 600202 671556
rect 612374 671544 612380 671556
rect 600196 671516 612380 671544
rect 600196 671504 600202 671516
rect 612374 671504 612380 671516
rect 612432 671504 612438 671556
rect 251642 671028 251648 671080
rect 251700 671068 251706 671080
rect 251700 671040 283934 671068
rect 251700 671028 251706 671040
rect 283906 671000 283934 671040
rect 286418 671000 286424 671012
rect 283906 670972 286424 671000
rect 286418 670960 286424 670972
rect 286476 670960 286482 671012
rect 341066 670416 341072 670468
rect 341124 670456 341130 670468
rect 352382 670456 352388 670468
rect 341124 670428 352388 670456
rect 341124 670416 341130 670428
rect 352382 670416 352388 670428
rect 352440 670416 352446 670468
rect 208126 669804 208132 669856
rect 208184 669844 208190 669856
rect 209046 669844 209052 669856
rect 208184 669816 209052 669844
rect 208184 669804 208190 669816
rect 209046 669804 209052 669816
rect 209104 669804 209110 669856
rect 610810 669328 610816 669380
rect 610868 669368 610874 669380
rect 617802 669368 617808 669380
rect 610868 669340 617808 669368
rect 610868 669328 610874 669340
rect 617802 669328 617808 669340
rect 617860 669328 617866 669380
rect 613386 668716 613392 668768
rect 613444 668756 613450 668768
rect 616974 668756 616980 668768
rect 613444 668728 616980 668756
rect 613444 668716 613450 668728
rect 616974 668716 616980 668728
rect 617032 668716 617038 668768
rect 489278 668240 489284 668292
rect 489336 668280 489342 668292
rect 516878 668280 516884 668292
rect 489336 668252 516884 668280
rect 489336 668240 489342 668252
rect 516878 668240 516884 668252
rect 516936 668240 516942 668292
rect 340928 667890 342850 667912
rect 340928 667818 341506 667890
rect 342830 667818 342850 667890
rect 252838 667764 252844 667816
rect 252896 667804 252902 667816
rect 286602 667804 286608 667816
rect 252896 667776 286608 667804
rect 252896 667764 252902 667776
rect 286602 667764 286608 667776
rect 286660 667804 286666 667816
rect 286878 667804 286884 667816
rect 286660 667776 286884 667804
rect 286660 667764 286666 667776
rect 286878 667764 286884 667776
rect 286936 667764 286942 667816
rect 340928 667794 342850 667818
rect 220034 667728 222160 667758
rect 209322 667560 209328 667612
rect 209380 667600 209386 667612
rect 210150 667600 210156 667612
rect 209380 667572 210156 667600
rect 209380 667560 209386 667572
rect 210150 667560 210156 667572
rect 210208 667560 210214 667612
rect 220034 667552 220076 667728
rect 222120 667677 222160 667728
rect 222120 667581 268866 667677
rect 615594 667628 615600 667680
rect 615652 667668 615658 667680
rect 618906 667668 618912 667680
rect 615652 667640 618912 667668
rect 615652 667628 615658 667640
rect 618906 667628 618912 667640
rect 618964 667628 618970 667680
rect 222120 667552 222160 667581
rect 335546 667560 335552 667612
rect 335604 667600 335610 667612
rect 342265 667603 342323 667609
rect 342265 667600 342277 667603
rect 335604 667572 342277 667600
rect 335604 667560 335610 667572
rect 342265 667569 342277 667572
rect 342311 667569 342323 667603
rect 342265 667563 342323 667569
rect 220034 667516 222160 667552
rect 342538 667532 342544 667544
rect 337404 667504 342544 667532
rect 240850 667368 256334 667396
rect 208126 667288 208132 667340
rect 208184 667328 208190 667340
rect 210058 667328 210064 667340
rect 208184 667300 210064 667328
rect 208184 667288 208190 667300
rect 210058 667288 210064 667300
rect 210116 667288 210122 667340
rect 228185 667331 228243 667337
rect 228185 667297 228197 667331
rect 228231 667328 228243 667331
rect 240850 667328 240878 667368
rect 228231 667300 240878 667328
rect 248425 667331 248483 667337
rect 228231 667297 228243 667300
rect 228185 667291 228243 667297
rect 248425 667297 248437 667331
rect 248471 667328 248483 667331
rect 256306 667328 256334 667368
rect 286878 667356 286884 667408
rect 286936 667396 286942 667408
rect 337294 667396 337300 667408
rect 286936 667368 337300 667396
rect 286936 667356 286942 667368
rect 337294 667356 337300 667368
rect 337352 667356 337358 667408
rect 268757 667331 268815 667337
rect 248471 667300 248606 667328
rect 256306 667300 264062 667328
rect 248471 667297 248483 667300
rect 248425 667291 248483 667297
rect 248578 667192 248606 667300
rect 264034 667260 264062 667300
rect 268757 667297 268769 667331
rect 268803 667328 268815 667331
rect 270226 667328 270232 667340
rect 268803 667300 270232 667328
rect 268803 667297 268815 667300
rect 268757 667291 268815 667297
rect 270226 667288 270232 667300
rect 270284 667288 270290 667340
rect 290742 667328 290748 667340
rect 271762 667300 290748 667328
rect 267390 667260 268230 667280
rect 271762 667260 271790 667300
rect 290742 667288 290748 667300
rect 290800 667288 290806 667340
rect 315490 667288 315496 667340
rect 315548 667328 315554 667340
rect 316042 667328 316048 667340
rect 315548 667300 316048 667328
rect 315548 667288 315554 667300
rect 316042 667288 316048 667300
rect 316100 667328 316106 667340
rect 337404 667328 337432 667504
rect 342538 667492 342544 667504
rect 342596 667492 342602 667544
rect 341066 667430 341072 667476
rect 340992 667424 341072 667430
rect 341124 667424 341130 667476
rect 338950 667356 338956 667408
rect 339008 667396 339014 667408
rect 340992 667402 341081 667424
rect 340992 667396 341020 667402
rect 339008 667368 341020 667396
rect 341069 667399 341081 667402
rect 341115 667399 341127 667424
rect 341069 667393 341127 667399
rect 342464 667368 372254 667396
rect 339008 667356 339014 667368
rect 342464 667328 342492 667368
rect 316100 667300 337432 667328
rect 337496 667300 342492 667328
rect 316100 667288 316106 667300
rect 303162 667260 303168 667272
rect 264034 667252 271790 667260
rect 264034 667232 267430 667252
rect 268196 667232 271790 667252
rect 279490 667232 303168 667260
rect 267834 667212 267840 667224
rect 267556 667192 267840 667212
rect 248578 667184 267840 667192
rect 248578 667164 267588 667184
rect 267834 667172 267840 667184
rect 267892 667172 267898 667224
rect 270226 667152 270232 667204
rect 270284 667192 270290 667204
rect 279490 667192 279518 667232
rect 303162 667220 303168 667232
rect 303220 667220 303226 667272
rect 337294 667220 337300 667272
rect 337352 667260 337358 667272
rect 337496 667260 337524 667300
rect 342538 667288 342544 667340
rect 342596 667328 342602 667340
rect 362318 667328 362324 667340
rect 342596 667300 362324 667328
rect 342596 667288 342602 667300
rect 362318 667288 362324 667300
rect 362376 667288 362382 667340
rect 372226 667328 372254 667368
rect 382926 667328 382932 667340
rect 372226 667300 382932 667328
rect 382926 667288 382932 667300
rect 382984 667288 382990 667340
rect 337352 667232 337524 667260
rect 337352 667220 337358 667232
rect 360478 667220 360484 667272
rect 360536 667260 360542 667272
rect 362410 667260 362416 667272
rect 360536 667232 362416 667260
rect 360536 667220 360542 667232
rect 362410 667220 362416 667232
rect 362468 667220 362474 667272
rect 270284 667164 279518 667192
rect 340914 667170 342572 667192
rect 270284 667152 270290 667164
rect 227016 667037 269080 667133
rect 308222 667084 308228 667136
rect 308280 667124 308286 667136
rect 321930 667124 321936 667136
rect 308280 667096 321936 667124
rect 308280 667084 308286 667096
rect 321930 667084 321936 667096
rect 321988 667084 321994 667136
rect 340914 667088 340998 667170
rect 342546 667088 342572 667170
rect 361122 667152 361128 667204
rect 361180 667192 361186 667204
rect 361858 667192 361864 667204
rect 361180 667164 361864 667192
rect 361180 667152 361186 667164
rect 361858 667152 361864 667164
rect 361916 667152 361922 667204
rect 362686 667152 362692 667204
rect 362744 667192 362750 667204
rect 363882 667192 363888 667204
rect 362744 667164 363888 667192
rect 362744 667152 362750 667164
rect 363882 667152 363888 667164
rect 363940 667152 363946 667204
rect 390102 667152 390108 667204
rect 390160 667192 390166 667204
rect 569226 667192 569232 667204
rect 390160 667164 569232 667192
rect 390160 667152 390166 667164
rect 569226 667152 569232 667164
rect 569284 667152 569290 667204
rect 635466 667152 635472 667204
rect 635524 667192 635530 667204
rect 643194 667192 643200 667204
rect 635524 667164 643200 667192
rect 635524 667152 635530 667164
rect 643194 667152 643200 667164
rect 643252 667152 643258 667204
rect 340914 667070 342572 667088
rect 342906 667084 342912 667136
rect 342964 667124 342970 667136
rect 342964 667096 345758 667124
rect 342964 667084 342970 667096
rect 236436 667020 243140 667037
rect 236436 665954 236536 667020
rect 242984 665954 243140 667020
rect 310154 667016 310160 667068
rect 310212 667056 310218 667068
rect 345730 667056 345758 667096
rect 361766 667084 361772 667136
rect 361824 667124 361830 667136
rect 381086 667124 381092 667136
rect 361824 667096 381092 667124
rect 361824 667084 361830 667096
rect 381086 667084 381092 667096
rect 381144 667084 381150 667136
rect 361214 667056 361220 667068
rect 310212 667028 336236 667056
rect 345730 667028 361220 667056
rect 310212 667016 310218 667028
rect 318158 666948 318164 667000
rect 318216 666988 318222 667000
rect 336208 666988 336236 667028
rect 361214 667016 361220 667028
rect 361272 667016 361278 667068
rect 342722 666988 342728 667000
rect 318216 666960 335776 666988
rect 336208 666960 342728 666988
rect 318216 666948 318222 666960
rect 297550 666880 297556 666932
rect 297608 666920 297614 666932
rect 335638 666920 335644 666932
rect 297608 666892 335644 666920
rect 297608 666880 297614 666892
rect 335638 666880 335644 666892
rect 335696 666880 335702 666932
rect 335748 666920 335776 666960
rect 342722 666948 342728 666960
rect 342780 666948 342786 667000
rect 342906 666948 342912 667000
rect 342964 666988 342970 667000
rect 375198 666988 375204 667000
rect 342964 666960 375204 666988
rect 342964 666948 342970 666960
rect 375198 666948 375204 666960
rect 375256 666948 375262 667000
rect 342814 666920 342820 666932
rect 335748 666892 342820 666920
rect 342814 666880 342820 666892
rect 342872 666880 342878 666932
rect 344102 666880 344108 666932
rect 344160 666920 344166 666932
rect 360478 666920 360484 666932
rect 344160 666892 360484 666920
rect 344160 666880 344166 666892
rect 360478 666880 360484 666892
rect 360536 666880 360542 666932
rect 361674 666880 361680 666932
rect 361732 666920 361738 666932
rect 368850 666920 368856 666932
rect 361732 666892 368856 666920
rect 361732 666880 361738 666892
rect 368850 666880 368856 666892
rect 368908 666920 368914 666932
rect 369126 666920 369132 666932
rect 368908 666892 369132 666920
rect 368908 666880 368914 666892
rect 369126 666880 369132 666892
rect 369184 666880 369190 666932
rect 290650 666812 290656 666864
rect 290708 666852 290714 666864
rect 390470 666852 390476 666864
rect 290708 666824 390476 666852
rect 290708 666812 290714 666824
rect 390470 666812 390476 666824
rect 390528 666812 390534 666864
rect 251550 666744 251556 666796
rect 251608 666784 251614 666796
rect 289362 666784 289368 666796
rect 251608 666756 289368 666784
rect 251608 666744 251614 666756
rect 289362 666744 289368 666756
rect 289420 666744 289426 666796
rect 298746 666744 298752 666796
rect 298804 666784 298810 666796
rect 373174 666784 373180 666796
rect 298804 666756 373180 666784
rect 298804 666744 298810 666756
rect 373174 666744 373180 666756
rect 373232 666744 373238 666796
rect 377130 666744 377136 666796
rect 377188 666784 377194 666796
rect 379246 666784 379252 666796
rect 377188 666756 379252 666784
rect 377188 666744 377194 666756
rect 379246 666744 379252 666756
rect 379304 666784 379310 666796
rect 576494 666784 576500 666796
rect 379304 666756 576500 666784
rect 379304 666744 379310 666756
rect 576494 666744 576500 666756
rect 576552 666744 576558 666796
rect 250538 666676 250544 666728
rect 250596 666716 250602 666728
rect 296170 666716 296176 666728
rect 250596 666688 296176 666716
rect 250596 666676 250602 666688
rect 296170 666676 296176 666688
rect 296228 666716 296234 666728
rect 377222 666716 377228 666728
rect 296228 666688 377228 666716
rect 296228 666676 296234 666688
rect 377222 666676 377228 666688
rect 377280 666676 377286 666728
rect 389366 666676 389372 666728
rect 389424 666716 389430 666728
rect 612926 666716 612932 666728
rect 389424 666688 612932 666716
rect 389424 666676 389430 666688
rect 612926 666676 612932 666688
rect 612984 666676 612990 666728
rect 252746 666608 252752 666660
rect 252804 666648 252810 666660
rect 290650 666648 290656 666660
rect 252804 666620 290656 666648
rect 252804 666608 252810 666620
rect 290650 666608 290656 666620
rect 290708 666608 290714 666660
rect 321010 666608 321016 666660
rect 321068 666648 321074 666660
rect 365078 666648 365084 666660
rect 321068 666620 365084 666648
rect 321068 666608 321074 666620
rect 365078 666608 365084 666620
rect 365136 666608 365142 666660
rect 385318 666608 385324 666660
rect 385376 666648 385382 666660
rect 615778 666648 615784 666660
rect 385376 666620 615784 666648
rect 385376 666608 385382 666620
rect 615778 666608 615784 666620
rect 615836 666608 615842 666660
rect 316870 666540 316876 666592
rect 316928 666580 316934 666592
rect 637214 666580 637220 666592
rect 316928 666552 637220 666580
rect 316928 666540 316934 666552
rect 637214 666540 637220 666552
rect 637272 666540 637278 666592
rect 314110 666472 314116 666524
rect 314168 666512 314174 666524
rect 598574 666512 598580 666524
rect 314168 666484 598580 666512
rect 314168 666472 314174 666484
rect 598574 666472 598580 666484
rect 598632 666472 598638 666524
rect 294790 666404 294796 666456
rect 294848 666444 294854 666456
rect 370506 666444 370512 666456
rect 294848 666416 370512 666444
rect 294848 666404 294854 666416
rect 370506 666404 370512 666416
rect 370564 666444 370570 666456
rect 371150 666444 371156 666456
rect 370564 666416 371156 666444
rect 370564 666404 370570 666416
rect 371150 666404 371156 666416
rect 371208 666404 371214 666456
rect 288258 666336 288264 666388
rect 288316 666376 288322 666388
rect 335546 666376 335552 666388
rect 288316 666348 335552 666376
rect 288316 666336 288322 666348
rect 335546 666336 335552 666348
rect 335604 666336 335610 666388
rect 335638 666336 335644 666388
rect 335696 666376 335702 666388
rect 344102 666376 344108 666388
rect 335696 666348 344108 666376
rect 335696 666336 335702 666348
rect 344102 666336 344108 666348
rect 344160 666336 344166 666388
rect 611178 666336 611184 666388
rect 611236 666376 611242 666388
rect 613386 666376 613392 666388
rect 611236 666348 613392 666376
rect 611236 666336 611242 666348
rect 613386 666336 613392 666348
rect 613444 666336 613450 666388
rect 290834 666268 290840 666320
rect 290892 666308 290898 666320
rect 298746 666308 298752 666320
rect 290892 666280 298752 666308
rect 290892 666268 290898 666280
rect 298746 666268 298752 666280
rect 298804 666268 298810 666320
rect 321286 666308 321292 666320
rect 310402 666280 321292 666308
rect 288534 666200 288540 666252
rect 288592 666240 288598 666252
rect 306474 666240 306480 666252
rect 288592 666212 306480 666240
rect 288592 666200 288598 666212
rect 306474 666200 306480 666212
rect 306532 666200 306538 666252
rect 252010 666132 252016 666184
rect 252068 666172 252074 666184
rect 310402 666172 310430 666280
rect 321286 666268 321292 666280
rect 321344 666308 321350 666320
rect 363238 666308 363244 666320
rect 321344 666280 363244 666308
rect 321344 666268 321350 666280
rect 363238 666268 363244 666280
rect 363296 666268 363302 666320
rect 375198 666200 375204 666252
rect 375256 666240 375262 666252
rect 605658 666240 605664 666252
rect 375256 666212 605664 666240
rect 375256 666200 375262 666212
rect 605658 666200 605664 666212
rect 605716 666200 605722 666252
rect 252068 666144 310430 666172
rect 252068 666132 252074 666144
rect 362502 666132 362508 666184
rect 362560 666172 362566 666184
rect 615594 666172 615600 666184
rect 362560 666144 615600 666172
rect 362560 666132 362566 666144
rect 615594 666132 615600 666144
rect 615652 666132 615658 666184
rect 288442 666064 288448 666116
rect 288500 666104 288506 666116
rect 594618 666104 594624 666116
rect 288500 666076 594624 666104
rect 288500 666064 288506 666076
rect 594618 666064 594624 666076
rect 594676 666064 594682 666116
rect 606854 666064 606860 666116
rect 606912 666104 606918 666116
rect 613478 666104 613484 666116
rect 606912 666076 613484 666104
rect 606912 666064 606918 666076
rect 613478 666064 613484 666076
rect 613536 666064 613542 666116
rect 288166 665996 288172 666048
rect 288224 666036 288230 666048
rect 598574 666036 598580 666048
rect 288224 666008 598580 666036
rect 288224 665996 288230 666008
rect 598574 665996 598580 666008
rect 598632 665996 598638 666048
rect 236436 665890 243140 665954
rect 290742 665860 290748 665912
rect 290800 665900 290806 665912
rect 321194 665900 321200 665912
rect 290800 665872 321200 665900
rect 290800 665860 290806 665872
rect 321194 665860 321200 665872
rect 321252 665860 321258 665912
rect 267834 665792 267840 665844
rect 267892 665832 267898 665844
rect 320918 665832 320924 665844
rect 267892 665804 320924 665832
rect 267892 665792 267898 665804
rect 320918 665792 320924 665804
rect 320976 665792 320982 665844
rect 251458 665520 251464 665572
rect 251516 665560 251522 665572
rect 290834 665560 290840 665572
rect 251516 665532 290840 665560
rect 251516 665520 251522 665532
rect 290834 665520 290840 665532
rect 290892 665520 290898 665572
rect 287982 665452 287988 665504
rect 288040 665492 288046 665504
rect 390286 665492 390292 665504
rect 288040 665464 390292 665492
rect 288040 665452 288046 665464
rect 390286 665452 390292 665464
rect 390344 665452 390350 665504
rect 320734 665384 320740 665436
rect 320792 665424 320798 665436
rect 389366 665424 389372 665436
rect 320792 665396 389372 665424
rect 320792 665384 320798 665396
rect 389366 665384 389372 665396
rect 389424 665384 389430 665436
rect 297826 665316 297832 665368
rect 297884 665356 297890 665368
rect 298838 665356 298844 665368
rect 297884 665328 298844 665356
rect 297884 665316 297890 665328
rect 298838 665316 298844 665328
rect 298896 665316 298902 665368
rect 304910 665316 304916 665368
rect 304968 665356 304974 665368
rect 305830 665356 305836 665368
rect 304968 665328 305836 665356
rect 304968 665316 304974 665328
rect 305830 665316 305836 665328
rect 305888 665316 305894 665368
rect 320826 665356 320832 665368
rect 310402 665328 320832 665356
rect 209046 665248 209052 665300
rect 209104 665288 209110 665300
rect 310402 665288 310430 665328
rect 320826 665316 320832 665328
rect 320884 665356 320890 665368
rect 377130 665356 377136 665368
rect 320884 665328 377136 665356
rect 320884 665316 320890 665328
rect 377130 665316 377136 665328
rect 377188 665316 377194 665368
rect 209104 665260 310430 665288
rect 209104 665248 209110 665260
rect 248514 665180 248520 665232
rect 248572 665220 248578 665232
rect 362870 665220 362876 665232
rect 248572 665192 362876 665220
rect 248572 665180 248578 665192
rect 362870 665180 362876 665192
rect 362928 665180 362934 665232
rect 378878 665180 378884 665232
rect 378936 665220 378942 665232
rect 506298 665220 506304 665232
rect 378936 665192 506304 665220
rect 378936 665180 378942 665192
rect 506298 665180 506304 665192
rect 506356 665180 506362 665232
rect 210150 665112 210156 665164
rect 210208 665152 210214 665164
rect 338950 665152 338956 665164
rect 210208 665124 338956 665152
rect 210208 665112 210214 665124
rect 338950 665112 338956 665124
rect 339008 665112 339014 665164
rect 362594 665112 362600 665164
rect 362652 665152 362658 665164
rect 532334 665152 532340 665164
rect 362652 665124 532340 665152
rect 362652 665112 362658 665124
rect 532334 665112 532340 665124
rect 532392 665112 532398 665164
rect 288074 665044 288080 665096
rect 288132 665084 288138 665096
rect 301598 665084 301604 665096
rect 288132 665056 301604 665084
rect 288132 665044 288138 665056
rect 301598 665044 301604 665056
rect 301656 665044 301662 665096
rect 304358 665044 304364 665096
rect 304416 665084 304422 665096
rect 610258 665084 610264 665096
rect 304416 665056 610264 665084
rect 304416 665044 304422 665056
rect 610258 665044 610264 665056
rect 610316 665044 610322 665096
rect 292030 664976 292036 665028
rect 292088 665016 292094 665028
rect 604646 665016 604652 665028
rect 292088 664988 604652 665016
rect 292088 664976 292094 664988
rect 604646 664976 604652 664988
rect 604704 664976 604710 665028
rect 289086 664908 289092 664960
rect 289144 664948 289150 664960
rect 615962 664948 615968 664960
rect 289144 664920 615968 664948
rect 289144 664908 289150 664920
rect 615962 664908 615968 664920
rect 616020 664908 616026 664960
rect 287890 664840 287896 664892
rect 287948 664880 287954 664892
rect 321470 664880 321476 664892
rect 287948 664852 321476 664880
rect 287948 664840 287954 664852
rect 321470 664840 321476 664852
rect 321528 664840 321534 664892
rect 319722 664772 319728 664824
rect 319780 664812 319786 664824
rect 367102 664812 367108 664824
rect 319780 664784 367108 664812
rect 319780 664772 319786 664784
rect 367102 664772 367108 664784
rect 367160 664772 367166 664824
rect 617894 664772 617900 664824
rect 617952 664812 617958 664824
rect 620010 664812 620016 664824
rect 617952 664784 620016 664812
rect 617952 664772 617958 664784
rect 620010 664772 620016 664784
rect 620068 664772 620074 664824
rect 608970 664500 608976 664552
rect 609028 664540 609034 664552
rect 612190 664540 612196 664552
rect 609028 664512 612196 664540
rect 609028 664500 609034 664512
rect 612190 664500 612196 664512
rect 612248 664500 612254 664552
rect 569226 663956 569232 664008
rect 569284 663996 569290 664008
rect 574746 663996 574752 664008
rect 569284 663968 574752 663996
rect 569284 663956 569290 663968
rect 574746 663956 574752 663968
rect 574804 663956 574810 664008
rect 675670 663956 675676 664008
rect 675728 663996 675734 664008
rect 676038 663996 676044 664008
rect 675728 663968 676044 663996
rect 675728 663956 675734 663968
rect 676038 663956 676044 663968
rect 676096 663956 676102 664008
rect 306474 663888 306480 663940
rect 306532 663928 306538 663940
rect 604554 663928 604560 663940
rect 306532 663900 604560 663928
rect 306532 663888 306538 663900
rect 604554 663888 604560 663900
rect 604612 663888 604618 663940
rect 300310 663820 300316 663872
rect 300368 663860 300374 663872
rect 610074 663860 610080 663872
rect 300368 663832 610080 663860
rect 300368 663820 300374 663832
rect 610074 663820 610080 663832
rect 610132 663820 610138 663872
rect 615594 663820 615600 663872
rect 615652 663860 615658 663872
rect 621298 663860 621304 663872
rect 615652 663832 621304 663860
rect 615652 663820 615658 663832
rect 621298 663820 621304 663832
rect 621356 663820 621362 663872
rect 676038 663820 676044 663872
rect 676096 663860 676102 663872
rect 676682 663860 676688 663872
rect 676096 663832 676688 663860
rect 676096 663820 676102 663832
rect 676682 663820 676688 663832
rect 676740 663820 676746 663872
rect 675854 663616 675860 663668
rect 675912 663656 675918 663668
rect 676222 663656 676228 663668
rect 675912 663628 676228 663656
rect 675912 663616 675918 663628
rect 676222 663616 676228 663628
rect 676280 663616 676286 663668
rect 676590 663036 676596 663048
rect 676357 663008 676596 663036
rect 675762 662936 675768 662988
rect 675820 662976 675826 662988
rect 676357 662976 676385 663008
rect 676590 662996 676596 663008
rect 676648 662996 676654 663048
rect 675820 662948 676385 662976
rect 675820 662936 675826 662948
rect 614490 662868 614496 662920
rect 614548 662908 614554 662920
rect 619090 662908 619096 662920
rect 614548 662880 619096 662908
rect 614548 662868 614554 662880
rect 619090 662868 619096 662880
rect 619148 662868 619154 662920
rect 252654 662732 252660 662784
rect 252712 662772 252718 662784
rect 293318 662772 293324 662784
rect 252712 662744 293324 662772
rect 252712 662732 252718 662744
rect 293318 662732 293324 662744
rect 293376 662732 293382 662784
rect 362410 662732 362416 662784
rect 362468 662772 362474 662784
rect 584222 662772 584228 662784
rect 362468 662744 584228 662772
rect 362468 662732 362474 662744
rect 584222 662732 584228 662744
rect 584280 662732 584286 662784
rect 604646 662732 604652 662784
rect 604704 662772 604710 662784
rect 614490 662772 614496 662784
rect 604704 662744 614496 662772
rect 604704 662732 604710 662744
rect 614490 662732 614496 662744
rect 614548 662732 614554 662784
rect 675670 662256 675676 662308
rect 675728 662296 675734 662308
rect 676130 662296 676136 662308
rect 675728 662268 676136 662296
rect 675728 662256 675734 662268
rect 676130 662256 676136 662268
rect 676188 662256 676194 662308
rect 671346 661916 671352 661968
rect 671404 661956 671410 661968
rect 676314 661956 676320 661968
rect 671404 661928 676320 661956
rect 671404 661916 671410 661928
rect 676314 661916 676320 661928
rect 676372 661916 676378 661968
rect 615686 661848 615692 661900
rect 615744 661888 615750 661900
rect 616790 661888 616796 661900
rect 615744 661860 616796 661888
rect 615744 661848 615750 661860
rect 616790 661848 616796 661860
rect 616848 661848 616854 661900
rect 604554 661712 604560 661764
rect 604612 661752 604618 661764
rect 610166 661752 610172 661764
rect 604612 661724 610172 661752
rect 604612 661712 604618 661724
rect 610166 661712 610172 661724
rect 610224 661712 610230 661764
rect 612098 661304 612104 661356
rect 612156 661344 612162 661356
rect 619366 661344 619372 661356
rect 612156 661316 619372 661344
rect 612156 661304 612162 661316
rect 619366 661304 619372 661316
rect 619424 661304 619430 661356
rect 251090 661100 251096 661152
rect 251148 661140 251154 661152
rect 671346 661140 671352 661152
rect 251148 661112 671352 661140
rect 251148 661100 251154 661112
rect 671346 661100 671352 661112
rect 671404 661100 671410 661152
rect 359006 660488 359012 660540
rect 359064 660528 359070 660540
rect 541166 660528 541172 660540
rect 359064 660500 541172 660528
rect 359064 660488 359070 660500
rect 541166 660488 541172 660500
rect 541224 660488 541230 660540
rect 675762 660284 675768 660336
rect 675820 660324 675826 660336
rect 676314 660324 676320 660336
rect 675820 660296 676320 660324
rect 675820 660284 675826 660296
rect 676314 660284 676320 660296
rect 676372 660284 676378 660336
rect 606762 660080 606768 660132
rect 606820 660120 606826 660132
rect 609154 660120 609160 660132
rect 606820 660092 609160 660120
rect 606820 660080 606826 660092
rect 609154 660080 609160 660092
rect 609212 660080 609218 660132
rect 613478 659468 613484 659520
rect 613536 659508 613542 659520
rect 618262 659508 618268 659520
rect 613536 659480 618268 659508
rect 613536 659468 613542 659480
rect 618262 659468 618268 659480
rect 618320 659468 618326 659520
rect 402062 659400 402068 659452
rect 402120 659440 402126 659452
rect 485966 659440 485972 659452
rect 402120 659412 485972 659440
rect 402120 659400 402126 659412
rect 485966 659400 485972 659412
rect 486024 659400 486030 659452
rect 614582 659400 614588 659452
rect 614640 659440 614646 659452
rect 615686 659440 615692 659452
rect 614640 659412 615692 659440
rect 614640 659400 614646 659412
rect 615686 659400 615692 659412
rect 615744 659400 615750 659452
rect 616974 659060 616980 659112
rect 617032 659100 617038 659112
rect 621482 659100 621488 659112
rect 617032 659072 621488 659100
rect 617032 659060 617038 659072
rect 621482 659060 621488 659072
rect 621540 659060 621546 659112
rect 610074 658924 610080 658976
rect 610132 658964 610138 658976
rect 612282 658964 612288 658976
rect 610132 658936 612288 658964
rect 610132 658924 610138 658936
rect 612282 658924 612288 658936
rect 612340 658924 612346 658976
rect 615778 658448 615784 658500
rect 615836 658488 615842 658500
rect 620102 658488 620108 658500
rect 615836 658460 620108 658488
rect 615836 658448 615842 658460
rect 620102 658448 620108 658460
rect 620160 658448 620166 658500
rect 615962 658380 615968 658432
rect 616020 658420 616026 658432
rect 621022 658420 621028 658432
rect 616020 658392 621028 658420
rect 616020 658380 616026 658392
rect 621022 658380 621028 658392
rect 621080 658380 621086 658432
rect 307118 658312 307124 658364
rect 307176 658352 307182 658364
rect 437482 658352 437488 658364
rect 307176 658324 437488 658352
rect 307176 658312 307182 658324
rect 437482 658312 437488 658324
rect 437540 658312 437546 658364
rect 468302 658312 468308 658364
rect 468360 658352 468366 658364
rect 522490 658352 522496 658364
rect 468360 658324 522496 658352
rect 468360 658312 468366 658324
rect 522490 658312 522496 658324
rect 522548 658312 522554 658364
rect 574746 658312 574752 658364
rect 574804 658352 574810 658364
rect 584682 658352 584688 658364
rect 574804 658324 584688 658352
rect 574804 658312 574810 658324
rect 584682 658312 584688 658324
rect 584740 658312 584746 658364
rect 675670 658108 675676 658160
rect 675728 658148 675734 658160
rect 676038 658148 676044 658160
rect 675728 658120 676044 658148
rect 675728 658108 675734 658120
rect 676038 658108 676044 658120
rect 676096 658108 676102 658160
rect 637674 657768 637680 657820
rect 637732 657808 637738 657820
rect 676222 657808 676228 657820
rect 637732 657780 676228 657808
rect 637732 657768 637738 657780
rect 676222 657768 676228 657780
rect 676280 657768 676286 657820
rect 675578 657360 675584 657412
rect 675636 657400 675642 657412
rect 676222 657400 676228 657412
rect 675636 657372 676228 657400
rect 675636 657360 675642 657372
rect 676222 657360 676228 657372
rect 676280 657360 676286 657412
rect 506390 657224 506396 657276
rect 506448 657264 506454 657276
rect 514026 657264 514032 657276
rect 506448 657236 514032 657264
rect 506448 657224 506454 657236
rect 514026 657224 514032 657236
rect 514084 657224 514090 657276
rect 610258 657224 610264 657276
rect 610316 657264 610322 657276
rect 618998 657264 619004 657276
rect 610316 657236 619004 657264
rect 610316 657224 610322 657236
rect 618998 657224 619004 657236
rect 619056 657224 619062 657276
rect 282922 657156 282928 657208
rect 282980 657196 282986 657208
rect 548894 657196 548900 657208
rect 282980 657168 548900 657196
rect 282980 657156 282986 657168
rect 548894 657156 548900 657168
rect 548952 657156 548958 657208
rect 594618 657156 594624 657208
rect 594676 657196 594682 657208
rect 612190 657196 612196 657208
rect 594676 657168 612196 657196
rect 594676 657156 594682 657168
rect 612190 657156 612196 657168
rect 612248 657156 612254 657208
rect 675578 656680 675584 656732
rect 675636 656720 675642 656732
rect 676314 656720 676320 656732
rect 675636 656692 676320 656720
rect 675636 656680 675642 656692
rect 676314 656680 676320 656692
rect 676372 656680 676378 656732
rect 605658 656204 605664 656256
rect 605716 656244 605722 656256
rect 614398 656244 614404 656256
rect 605716 656216 614404 656244
rect 605716 656204 605722 656216
rect 614398 656204 614404 656216
rect 614456 656204 614462 656256
rect 675854 656204 675860 656256
rect 675912 656244 675918 656256
rect 676314 656244 676320 656256
rect 675912 656216 676320 656244
rect 675912 656204 675918 656216
rect 676314 656204 676320 656216
rect 676372 656204 676378 656256
rect 248422 656136 248428 656188
rect 248480 656176 248486 656188
rect 522582 656176 522588 656188
rect 248480 656148 522588 656176
rect 248480 656136 248486 656148
rect 522582 656136 522588 656148
rect 522640 656136 522646 656188
rect 584682 656136 584688 656188
rect 584740 656176 584746 656188
rect 595722 656176 595728 656188
rect 584740 656148 595728 656176
rect 584740 656136 584746 656148
rect 595722 656136 595728 656148
rect 595780 656136 595786 656188
rect 247318 656068 247324 656120
rect 247376 656108 247382 656120
rect 312638 656108 312644 656120
rect 247376 656080 312644 656108
rect 247376 656068 247382 656080
rect 312638 656068 312644 656080
rect 312696 656068 312702 656120
rect 315950 656068 315956 656120
rect 316008 656108 316014 656120
rect 624426 656108 624432 656120
rect 316008 656080 624432 656108
rect 316008 656068 316014 656080
rect 624426 656068 624432 656080
rect 624484 656068 624490 656120
rect 675762 656000 675768 656052
rect 675820 656040 675826 656052
rect 676130 656040 676136 656052
rect 675820 656012 676136 656040
rect 675820 656000 675826 656012
rect 676130 656000 676136 656012
rect 676188 656000 676194 656052
rect 675670 655592 675676 655644
rect 675728 655632 675734 655644
rect 676314 655632 676320 655644
rect 675728 655604 676320 655632
rect 675728 655592 675734 655604
rect 676314 655592 676320 655604
rect 676372 655592 676378 655644
rect 610166 655048 610172 655100
rect 610224 655088 610230 655100
rect 615502 655088 615508 655100
rect 610224 655060 615508 655088
rect 610224 655048 610230 655060
rect 615502 655048 615508 655060
rect 615560 655048 615566 655100
rect 620102 654912 620108 654964
rect 620160 654952 620166 654964
rect 622126 654952 622132 654964
rect 620160 654924 622132 654952
rect 620160 654912 620166 654924
rect 622126 654912 622132 654924
rect 622184 654912 622190 654964
rect 621482 654708 621488 654760
rect 621540 654748 621546 654760
rect 623138 654748 623144 654760
rect 621540 654720 623144 654748
rect 621540 654708 621546 654720
rect 623138 654708 623144 654720
rect 623196 654708 623202 654760
rect 213462 654504 213468 654556
rect 213520 654544 213526 654556
rect 619274 654544 619280 654556
rect 213520 654516 619280 654544
rect 213520 654504 213526 654516
rect 619274 654504 619280 654516
rect 619332 654504 619338 654556
rect 675486 654232 675492 654284
rect 675544 654272 675550 654284
rect 675946 654272 675952 654284
rect 675544 654244 675952 654272
rect 675544 654232 675550 654244
rect 675946 654232 675952 654244
rect 676004 654232 676010 654284
rect 675762 654164 675768 654216
rect 675820 654204 675826 654216
rect 676038 654204 676044 654216
rect 675820 654176 676044 654204
rect 675820 654164 675826 654176
rect 676038 654164 676044 654176
rect 676096 654164 676102 654216
rect 258542 653960 258548 654012
rect 258600 654000 258606 654012
rect 413102 654000 413108 654012
rect 258600 653972 413108 654000
rect 258600 653960 258606 653972
rect 413102 653960 413108 653972
rect 413160 653960 413166 654012
rect 501422 653960 501428 654012
rect 501480 654000 501486 654012
rect 546686 654000 546692 654012
rect 501480 653972 546692 654000
rect 501480 653960 501486 653972
rect 546686 653960 546692 653972
rect 546744 653960 546750 654012
rect 618262 653960 618268 654012
rect 618320 654000 618326 654012
rect 619458 654000 619464 654012
rect 618320 653972 619464 654000
rect 618320 653960 618326 653972
rect 619458 653960 619464 653972
rect 619516 653960 619522 654012
rect 250262 653892 250268 653944
rect 250320 653932 250326 653944
rect 519178 653932 519184 653944
rect 250320 653904 519184 653932
rect 250320 653892 250326 653904
rect 519178 653892 519184 653904
rect 519236 653892 519242 653944
rect 553310 653892 553316 653944
rect 553368 653932 553374 653944
rect 617894 653932 617900 653944
rect 553368 653904 617900 653932
rect 553368 653892 553374 653904
rect 617894 653892 617900 653904
rect 617952 653892 617958 653944
rect 620010 653620 620016 653672
rect 620068 653660 620074 653672
rect 622586 653660 622592 653672
rect 620068 653632 622592 653660
rect 620068 653620 620074 653632
rect 622586 653620 622592 653632
rect 622644 653620 622650 653672
rect 250998 652940 251004 652992
rect 251056 652980 251062 652992
rect 440702 652980 440708 652992
rect 251056 652952 440708 652980
rect 251056 652940 251062 652952
rect 440702 652940 440708 652952
rect 440760 652940 440766 652992
rect 250078 652872 250084 652924
rect 250136 652912 250142 652924
rect 459470 652912 459476 652924
rect 250136 652884 459476 652912
rect 250136 652872 250142 652884
rect 459470 652872 459476 652884
rect 459528 652872 459534 652924
rect 517982 652872 517988 652924
rect 518040 652912 518046 652924
rect 529206 652912 529212 652924
rect 518040 652884 529212 652912
rect 518040 652872 518046 652884
rect 529206 652872 529212 652884
rect 529264 652872 529270 652924
rect 609154 652872 609160 652924
rect 609212 652912 609218 652924
rect 615594 652912 615600 652924
rect 609212 652884 615600 652912
rect 609212 652872 609218 652884
rect 615594 652872 615600 652884
rect 615652 652872 615658 652924
rect 368850 652804 368856 652856
rect 368908 652844 368914 652856
rect 622954 652844 622960 652856
rect 368908 652816 622960 652844
rect 368908 652804 368914 652816
rect 622954 652804 622960 652816
rect 623012 652804 623018 652856
rect 361122 652736 361128 652788
rect 361180 652776 361186 652788
rect 621666 652776 621672 652788
rect 361180 652748 621672 652776
rect 361180 652736 361186 652748
rect 621666 652736 621672 652748
rect 621724 652736 621730 652788
rect 676222 652436 676228 652448
rect 673618 652408 676228 652436
rect 616698 652328 616704 652380
rect 616756 652368 616762 652380
rect 619182 652368 619188 652380
rect 616756 652340 619188 652368
rect 616756 652328 616762 652340
rect 619182 652328 619188 652340
rect 619240 652328 619246 652380
rect 673618 652368 673646 652408
rect 676222 652396 676228 652408
rect 676280 652396 676286 652448
rect 670306 652340 673646 652368
rect 208126 652260 208132 652312
rect 208184 652300 208190 652312
rect 209966 652300 209972 652312
rect 208184 652272 209972 652300
rect 208184 652260 208190 652272
rect 209966 652260 209972 652272
rect 210024 652260 210030 652312
rect 633258 652260 633264 652312
rect 633316 652300 633322 652312
rect 670306 652300 670334 652340
rect 633316 652272 670334 652300
rect 633316 652260 633322 652272
rect 208954 652056 208960 652108
rect 209012 652096 209018 652108
rect 209138 652096 209144 652108
rect 209012 652068 209144 652096
rect 209012 652056 209018 652068
rect 209138 652056 209144 652068
rect 209196 652056 209202 652108
rect 619090 651920 619096 651972
rect 619148 651960 619154 651972
rect 621114 651960 621120 651972
rect 619148 651932 621120 651960
rect 619148 651920 619154 651932
rect 621114 651920 621120 651932
rect 621172 651920 621178 651972
rect 250354 651784 250360 651836
rect 250412 651824 250418 651836
rect 419910 651824 419916 651836
rect 250412 651796 419916 651824
rect 250412 651784 250418 651796
rect 419910 651784 419916 651796
rect 419968 651784 419974 651836
rect 615686 651784 615692 651836
rect 615744 651824 615750 651836
rect 620838 651824 620844 651836
rect 615744 651796 620844 651824
rect 615744 651784 615750 651796
rect 620838 651784 620844 651796
rect 620896 651784 620902 651836
rect 251826 651716 251832 651768
rect 251884 651756 251890 651768
rect 431870 651756 431876 651768
rect 251884 651728 431876 651756
rect 251884 651716 251890 651728
rect 431870 651716 431876 651728
rect 431928 651716 431934 651768
rect 595722 651716 595728 651768
rect 595780 651756 595786 651768
rect 607866 651756 607872 651768
rect 595780 651728 607872 651756
rect 595780 651716 595786 651728
rect 607866 651716 607872 651728
rect 607924 651716 607930 651768
rect 249250 651648 249256 651700
rect 249308 651688 249314 651700
rect 463978 651688 463984 651700
rect 249308 651660 463984 651688
rect 249308 651648 249314 651660
rect 463978 651648 463984 651660
rect 464036 651648 464042 651700
rect 561222 651648 561228 651700
rect 561280 651688 561286 651700
rect 652670 651688 652676 651700
rect 561280 651660 652676 651688
rect 561280 651648 561286 651660
rect 652670 651648 652676 651660
rect 652728 651648 652734 651700
rect 668586 651648 668592 651700
rect 668644 651688 668650 651700
rect 676038 651688 676044 651700
rect 668644 651660 676044 651688
rect 668644 651648 668650 651660
rect 676038 651648 676044 651660
rect 676096 651648 676102 651700
rect 675578 651580 675584 651632
rect 675636 651620 675642 651632
rect 675854 651620 675860 651632
rect 675636 651592 675860 651620
rect 675636 651580 675642 651592
rect 675854 651580 675860 651592
rect 675912 651580 675918 651632
rect 675762 651376 675768 651428
rect 675820 651416 675826 651428
rect 676222 651416 676228 651428
rect 675820 651388 676228 651416
rect 675820 651376 675826 651388
rect 676222 651376 676228 651388
rect 676280 651376 676286 651428
rect 615594 651036 615600 651088
rect 615652 651076 615658 651088
rect 621390 651076 621396 651088
rect 615652 651048 621396 651076
rect 615652 651036 615658 651048
rect 621390 651036 621396 651048
rect 621448 651036 621454 651088
rect 618998 650832 619004 650884
rect 619056 650872 619062 650884
rect 622218 650872 622224 650884
rect 619056 650844 622224 650872
rect 619056 650832 619062 650844
rect 622218 650832 622224 650844
rect 622276 650832 622282 650884
rect 495902 650764 495908 650816
rect 495960 650804 495966 650816
rect 615594 650804 615600 650816
rect 495960 650776 615600 650804
rect 495960 650764 495966 650776
rect 615594 650764 615600 650776
rect 615652 650764 615658 650816
rect 619366 650764 619372 650816
rect 619424 650804 619430 650816
rect 622402 650804 622408 650816
rect 619424 650776 622408 650804
rect 619424 650764 619430 650776
rect 622402 650764 622408 650776
rect 622460 650764 622466 650816
rect 390010 650696 390016 650748
rect 390068 650736 390074 650748
rect 621850 650736 621856 650748
rect 390068 650708 621856 650736
rect 390068 650696 390074 650708
rect 621850 650696 621856 650708
rect 621908 650696 621914 650748
rect 389918 650628 389924 650680
rect 389976 650668 389982 650680
rect 613294 650668 613300 650680
rect 389976 650640 613300 650668
rect 389976 650628 389982 650640
rect 613294 650628 613300 650640
rect 613352 650628 613358 650680
rect 613386 650628 613392 650680
rect 613444 650668 613450 650680
rect 620930 650668 620936 650680
rect 613444 650640 620936 650668
rect 613444 650628 613450 650640
rect 620930 650628 620936 650640
rect 620988 650628 620994 650680
rect 370506 650560 370512 650612
rect 370564 650600 370570 650612
rect 619734 650600 619740 650612
rect 370564 650572 619740 650600
rect 370564 650560 370570 650572
rect 619734 650560 619740 650572
rect 619792 650560 619798 650612
rect 615594 650492 615600 650544
rect 615652 650532 615658 650544
rect 621942 650532 621948 650544
rect 615652 650504 621948 650532
rect 615652 650492 615658 650504
rect 621942 650492 621948 650504
rect 622000 650492 622006 650544
rect 613294 650424 613300 650476
rect 613352 650464 613358 650476
rect 622862 650464 622868 650476
rect 613352 650436 622868 650464
rect 613352 650424 613358 650436
rect 622862 650424 622868 650436
rect 622920 650424 622926 650476
rect 612098 650356 612104 650408
rect 612156 650396 612162 650408
rect 618998 650396 619004 650408
rect 612156 650368 619004 650396
rect 612156 650356 612162 650368
rect 618998 650356 619004 650368
rect 619056 650356 619062 650408
rect 676130 650362 676136 650414
rect 676188 650402 676194 650414
rect 676188 650374 676437 650402
rect 676188 650362 676194 650374
rect 614490 650288 614496 650340
rect 614548 650328 614554 650340
rect 622494 650328 622500 650340
rect 614548 650300 622500 650328
rect 614548 650288 614554 650300
rect 622494 650288 622500 650300
rect 622552 650288 622558 650340
rect 217050 650084 217056 650136
rect 217108 650124 217114 650136
rect 551654 650124 551660 650136
rect 217108 650096 551660 650124
rect 217108 650084 217114 650096
rect 551654 650084 551660 650096
rect 551712 650084 551718 650136
rect 607866 649540 607872 649592
rect 607924 649580 607930 649592
rect 619090 649580 619096 649592
rect 607924 649552 619096 649580
rect 607924 649540 607930 649552
rect 619090 649540 619096 649552
rect 619148 649540 619154 649592
rect 514026 649472 514032 649524
rect 514084 649512 514090 649524
rect 514084 649484 611822 649512
rect 514084 649472 514090 649484
rect 611794 649444 611822 649484
rect 617802 649472 617808 649524
rect 617860 649512 617866 649524
rect 621206 649512 621212 649524
rect 617860 649484 621212 649512
rect 617860 649472 617866 649484
rect 621206 649472 621212 649484
rect 621264 649472 621270 649524
rect 623046 649444 623052 649456
rect 611794 649416 623052 649444
rect 623046 649404 623052 649416
rect 623104 649404 623110 649456
rect 569226 649064 569232 649116
rect 569284 649104 569290 649116
rect 676222 649104 676228 649116
rect 569284 649076 676228 649104
rect 569284 649064 569290 649076
rect 676222 649064 676228 649076
rect 676280 649064 676286 649116
rect 252286 648996 252292 649048
rect 252344 649036 252350 649048
rect 675854 649036 675860 649048
rect 252344 649008 675860 649036
rect 252344 648996 252350 649008
rect 675854 648996 675860 649008
rect 675912 648996 675918 649048
rect 675486 648928 675492 648980
rect 675544 648968 675550 648980
rect 675946 648968 675952 648980
rect 675544 648940 675952 648968
rect 675544 648928 675550 648940
rect 675946 648928 675952 648940
rect 676004 648928 676010 648980
rect 615502 648724 615508 648776
rect 615560 648764 615566 648776
rect 619918 648764 619924 648776
rect 615560 648736 619924 648764
rect 615560 648724 615566 648736
rect 619918 648724 619924 648736
rect 619976 648724 619982 648776
rect 248054 648656 248060 648708
rect 248112 648696 248118 648708
rect 304910 648696 304916 648708
rect 248112 648668 304916 648696
rect 248112 648656 248118 648668
rect 304910 648656 304916 648668
rect 304968 648656 304974 648708
rect 249434 648588 249440 648640
rect 249492 648628 249498 648640
rect 316042 648628 316048 648640
rect 249492 648600 316048 648628
rect 249492 648588 249498 648600
rect 316042 648588 316048 648600
rect 316100 648588 316106 648640
rect 252562 648520 252568 648572
rect 252620 648560 252626 648572
rect 319722 648560 319728 648572
rect 252620 648532 319728 648560
rect 252620 648520 252626 648532
rect 319722 648520 319728 648532
rect 319780 648520 319786 648572
rect 248238 648452 248244 648504
rect 248296 648492 248302 648504
rect 321102 648492 321108 648504
rect 248296 648464 321108 648492
rect 248296 648452 248302 648464
rect 321102 648452 321108 648464
rect 321160 648452 321166 648504
rect 470142 648452 470148 648504
rect 470200 648492 470206 648504
rect 569226 648492 569232 648504
rect 470200 648464 569232 648492
rect 470200 648452 470206 648464
rect 569226 648452 569232 648464
rect 569284 648452 569290 648504
rect 248330 648384 248336 648436
rect 248388 648424 248394 648436
rect 324782 648424 324788 648436
rect 248388 648396 324788 648424
rect 248388 648384 248394 648396
rect 324782 648384 324788 648396
rect 324840 648384 324846 648436
rect 494798 648384 494804 648436
rect 494856 648424 494862 648436
rect 494856 648396 611822 648424
rect 494856 648384 494862 648396
rect 611794 648356 611822 648396
rect 618906 648384 618912 648436
rect 618964 648424 618970 648436
rect 620654 648424 620660 648436
rect 618964 648396 620660 648424
rect 618964 648384 618970 648396
rect 620654 648384 620660 648396
rect 620712 648384 620718 648436
rect 628842 648384 628848 648436
rect 628900 648424 628906 648436
rect 635466 648424 635472 648436
rect 628900 648396 635472 648424
rect 628900 648384 628906 648396
rect 635466 648384 635472 648396
rect 635524 648384 635530 648436
rect 622034 648356 622040 648368
rect 611794 648328 622040 648356
rect 622034 648316 622040 648328
rect 622092 648316 622098 648368
rect 374278 647976 374284 648028
rect 374336 648016 374342 648028
rect 624426 648016 624432 648028
rect 374336 647988 624432 648016
rect 374336 647976 374342 647988
rect 624426 647976 624432 647988
rect 624484 647976 624490 648028
rect 233610 647908 233616 647960
rect 233668 647948 233674 647960
rect 623230 647948 623236 647960
rect 233668 647920 623236 647948
rect 233668 647908 233674 647920
rect 623230 647908 623236 647920
rect 623288 647908 623294 647960
rect 252470 647840 252476 647892
rect 252528 647880 252534 647892
rect 671070 647880 671076 647892
rect 252528 647852 671076 647880
rect 252528 647840 252534 647852
rect 671070 647840 671076 647852
rect 671128 647840 671134 647892
rect 223674 647568 223680 647620
rect 223732 647608 223738 647620
rect 622310 647608 622316 647620
rect 223732 647580 622316 647608
rect 223732 647568 223738 647580
rect 622310 647568 622316 647580
rect 622368 647568 622374 647620
rect 252102 647432 252108 647484
rect 252160 647472 252166 647484
rect 320642 647472 320648 647484
rect 252160 647444 320648 647472
rect 252160 647432 252166 647444
rect 320642 647432 320648 647444
rect 320700 647432 320706 647484
rect 381086 647432 381092 647484
rect 381144 647472 381150 647484
rect 388630 647472 388636 647484
rect 381144 647444 388636 647472
rect 381144 647432 381150 647444
rect 388630 647432 388636 647444
rect 388688 647432 388694 647484
rect 405374 647432 405380 647484
rect 405432 647472 405438 647484
rect 426902 647472 426908 647484
rect 405432 647444 426908 647472
rect 405432 647432 405438 647444
rect 426902 647432 426908 647444
rect 426960 647432 426966 647484
rect 479710 647432 479716 647484
rect 479768 647472 479774 647484
rect 625530 647472 625536 647484
rect 479768 647444 625536 647472
rect 479768 647432 479774 647444
rect 625530 647432 625536 647444
rect 625588 647432 625594 647484
rect 252194 647364 252200 647416
rect 252252 647404 252258 647416
rect 321010 647404 321016 647416
rect 252252 647376 321016 647404
rect 252252 647364 252258 647376
rect 321010 647364 321016 647376
rect 321068 647364 321074 647416
rect 363882 647364 363888 647416
rect 363940 647404 363946 647416
rect 412550 647404 412556 647416
rect 363940 647376 412556 647404
rect 363940 647364 363946 647376
rect 412550 647364 412556 647376
rect 412608 647364 412614 647416
rect 494062 647364 494068 647416
rect 494120 647404 494126 647416
rect 645402 647404 645408 647416
rect 494120 647376 645408 647404
rect 494120 647364 494126 647376
rect 645402 647364 645408 647376
rect 645460 647364 645466 647416
rect 219258 647296 219264 647348
rect 219316 647336 219322 647348
rect 288810 647336 288816 647348
rect 219316 647308 288816 647336
rect 219316 647296 219322 647308
rect 288810 647296 288816 647308
rect 288868 647296 288874 647348
rect 365262 647296 365268 647348
rect 365320 647336 365326 647348
rect 383846 647336 383852 647348
rect 365320 647308 383852 647336
rect 365320 647296 365326 647308
rect 383846 647296 383852 647308
rect 383904 647296 383910 647348
rect 390378 647296 390384 647348
rect 390436 647336 390442 647348
rect 619826 647336 619832 647348
rect 390436 647308 619832 647336
rect 390436 647296 390442 647308
rect 619826 647296 619832 647308
rect 619884 647296 619890 647348
rect 251366 647228 251372 647280
rect 251424 647268 251430 647280
rect 544478 647268 544484 647280
rect 251424 647240 544484 647268
rect 251424 647228 251430 647240
rect 544478 647228 544484 647240
rect 544536 647228 544542 647280
rect 594710 647228 594716 647280
rect 594768 647268 594774 647280
rect 642090 647268 642096 647280
rect 594768 647240 642096 647268
rect 594768 647228 594774 647240
rect 642090 647228 642096 647240
rect 642148 647228 642154 647280
rect 320550 647160 320556 647212
rect 320608 647200 320614 647212
rect 503630 647200 503636 647212
rect 320608 647172 503636 647200
rect 320608 647160 320614 647172
rect 503630 647160 503636 647172
rect 503688 647160 503694 647212
rect 556438 647160 556444 647212
rect 556496 647200 556502 647212
rect 620746 647200 620752 647212
rect 556496 647172 620752 647200
rect 556496 647160 556502 647172
rect 620746 647160 620752 647172
rect 620804 647160 620810 647212
rect 288810 647092 288816 647144
rect 288868 647132 288874 647144
rect 407766 647132 407772 647144
rect 288868 647104 407772 647132
rect 288868 647092 288874 647104
rect 407766 647092 407772 647104
rect 407824 647092 407830 647144
rect 455790 647092 455796 647144
rect 455848 647132 455854 647144
rect 640986 647132 640992 647144
rect 455848 647104 640992 647132
rect 455848 647092 455854 647104
rect 640986 647092 640992 647104
rect 641044 647092 641050 647144
rect 297550 647024 297556 647076
rect 297608 647064 297614 647076
rect 308222 647064 308228 647076
rect 297608 647036 308228 647064
rect 297608 647024 297614 647036
rect 308222 647024 308228 647036
rect 308280 647024 308286 647076
rect 320458 647024 320464 647076
rect 320516 647064 320522 647076
rect 393414 647064 393420 647076
rect 320516 647036 393420 647064
rect 320516 647024 320522 647036
rect 393414 647024 393420 647036
rect 393472 647024 393478 647076
rect 398198 647024 398204 647076
rect 398256 647064 398262 647076
rect 671898 647064 671904 647076
rect 398256 647036 671904 647064
rect 398256 647024 398262 647036
rect 671898 647024 671904 647036
rect 671956 647024 671962 647076
rect 241338 646956 241344 647008
rect 241396 646996 241402 647008
rect 619366 646996 619372 647008
rect 241396 646968 619372 646996
rect 241396 646956 241402 646968
rect 619366 646956 619372 646968
rect 619424 646956 619430 647008
rect 675670 646956 675676 647008
rect 675728 646996 675734 647008
rect 676314 646996 676320 647008
rect 675728 646968 676320 646996
rect 675728 646956 675734 646968
rect 676314 646956 676320 646968
rect 676372 646956 676378 647008
rect 292766 646888 292772 646940
rect 292824 646928 292830 646940
rect 323034 646928 323040 646940
rect 292824 646900 323040 646928
rect 292824 646888 292830 646900
rect 323034 646888 323040 646900
rect 323092 646888 323098 646940
rect 326254 646888 326260 646940
rect 326312 646928 326318 646940
rect 635466 646928 635472 646940
rect 326312 646900 635472 646928
rect 326312 646888 326318 646900
rect 635466 646888 635472 646900
rect 635524 646888 635530 646940
rect 252378 646820 252384 646872
rect 252436 646860 252442 646872
rect 255690 646860 255696 646872
rect 252436 646832 255696 646860
rect 252436 646820 252442 646832
rect 255690 646820 255696 646832
rect 255748 646820 255754 646872
rect 609062 646820 609068 646872
rect 609120 646860 609126 646872
rect 631050 646860 631056 646872
rect 609120 646832 631056 646860
rect 609120 646820 609126 646832
rect 631050 646820 631056 646832
rect 631108 646820 631114 646872
rect 208402 646752 208408 646804
rect 208460 646792 208466 646804
rect 268662 646792 268668 646804
rect 208460 646764 268668 646792
rect 208460 646752 208466 646764
rect 268662 646752 268668 646764
rect 268720 646752 268726 646804
rect 273630 646752 273636 646804
rect 273688 646792 273694 646804
rect 297826 646792 297832 646804
rect 273688 646764 297832 646792
rect 273688 646752 273694 646764
rect 297826 646752 297832 646764
rect 297884 646752 297890 646804
rect 311902 646752 311908 646804
rect 311960 646792 311966 646804
rect 638778 646792 638784 646804
rect 311960 646764 638784 646792
rect 311960 646752 311966 646764
rect 638778 646752 638784 646764
rect 638836 646752 638842 646804
rect 676222 646752 676228 646804
rect 676280 646752 676286 646804
rect 676240 646532 676268 646752
rect 676222 646480 676228 646532
rect 676280 646480 676286 646532
rect 671070 646140 671076 646192
rect 671128 646180 671134 646192
rect 676130 646180 676136 646192
rect 671128 646152 676136 646180
rect 671128 646140 671134 646152
rect 676130 646140 676136 646152
rect 676188 646140 676194 646192
rect 666746 645936 666752 645988
rect 666804 645976 666810 645988
rect 676590 645976 676596 645988
rect 666804 645948 676596 645976
rect 666804 645936 666810 645948
rect 676590 645936 676596 645948
rect 676648 645936 676654 645988
rect 208310 644984 208316 645036
rect 208368 645024 208374 645036
rect 210058 645024 210064 645036
rect 208368 644996 210064 645024
rect 208368 644984 208374 644996
rect 210058 644984 210064 644996
rect 210116 644984 210122 645036
rect 675762 644780 675768 644832
rect 675820 644820 675826 644832
rect 676498 644820 676504 644832
rect 675820 644792 676504 644820
rect 675820 644780 675826 644792
rect 676498 644780 676504 644792
rect 676556 644780 676562 644832
rect 209414 643964 209420 644016
rect 209472 644004 209478 644016
rect 233610 644004 233616 644016
rect 209472 643976 233616 644004
rect 209472 643964 209478 643976
rect 233610 643964 233616 643976
rect 233668 643964 233674 644016
rect 675578 643896 675584 643948
rect 675636 643936 675642 643948
rect 676406 643936 676412 643948
rect 675636 643908 676412 643936
rect 675636 643896 675642 643908
rect 676406 643896 676412 643908
rect 676464 643896 676470 643948
rect 208034 640700 208040 640752
rect 208092 640740 208098 640752
rect 208678 640740 208684 640752
rect 208092 640712 208684 640740
rect 208092 640700 208098 640712
rect 208678 640700 208684 640712
rect 208736 640700 208742 640752
rect 208586 640632 208592 640684
rect 208644 640672 208650 640684
rect 209966 640672 209972 640684
rect 208644 640644 209972 640672
rect 208644 640632 208650 640644
rect 209966 640632 209972 640644
rect 210024 640632 210030 640684
rect 208218 640292 208224 640344
rect 208276 640332 208282 640344
rect 208862 640332 208868 640344
rect 208276 640304 208868 640332
rect 208276 640292 208282 640304
rect 208862 640292 208868 640304
rect 208920 640292 208926 640344
rect 208218 639884 208224 639936
rect 208276 639924 208282 639936
rect 208770 639924 208776 639936
rect 208276 639896 208776 639924
rect 208276 639884 208282 639896
rect 208770 639884 208776 639896
rect 208828 639884 208834 639936
rect 208034 638932 208040 638984
rect 208092 638972 208098 638984
rect 208954 638972 208960 638984
rect 208092 638944 208960 638972
rect 208092 638932 208098 638944
rect 208954 638932 208960 638944
rect 209012 638932 209018 638984
rect 209322 638388 209328 638440
rect 209380 638428 209386 638440
rect 223674 638428 223680 638440
rect 209380 638400 223680 638428
rect 209380 638388 209386 638400
rect 223674 638388 223680 638400
rect 223732 638388 223738 638440
rect 661962 637844 661968 637896
rect 662020 637884 662026 637896
rect 668586 637884 668592 637896
rect 662020 637856 668592 637884
rect 662020 637844 662026 637856
rect 668586 637844 668592 637856
rect 668644 637844 668650 637896
rect 208678 636756 208684 636808
rect 208736 636796 208742 636808
rect 208862 636796 208868 636808
rect 208736 636768 208868 636796
rect 208736 636756 208742 636768
rect 208862 636756 208868 636768
rect 208920 636756 208926 636808
rect 208770 636688 208776 636740
rect 208828 636728 208834 636740
rect 209138 636728 209144 636740
rect 208828 636700 209144 636728
rect 208828 636688 208834 636700
rect 209138 636688 209144 636700
rect 209196 636688 209202 636740
rect 208402 636620 208408 636672
rect 208460 636660 208466 636672
rect 208460 636632 208816 636660
rect 208460 636620 208466 636632
rect 208788 636604 208816 636632
rect 208310 636552 208316 636604
rect 208368 636592 208374 636604
rect 208678 636592 208684 636604
rect 208368 636564 208684 636592
rect 208368 636552 208374 636564
rect 208678 636552 208684 636564
rect 208736 636552 208742 636604
rect 208770 636552 208776 636604
rect 208828 636552 208834 636604
rect 208034 636484 208040 636536
rect 208092 636524 208098 636536
rect 208494 636524 208500 636536
rect 208092 636496 208500 636524
rect 208092 636484 208098 636496
rect 208494 636484 208500 636496
rect 208552 636484 208558 636536
rect 208954 635640 208960 635652
rect 208052 635626 208960 635640
rect 207962 635612 208960 635626
rect 207962 635598 208080 635612
rect 208954 635600 208960 635612
rect 209012 635600 209018 635652
rect 623322 635124 623328 635176
rect 623380 635164 623386 635176
rect 628842 635164 628848 635176
rect 623380 635136 628848 635164
rect 623380 635124 623386 635136
rect 628842 635124 628848 635136
rect 628900 635124 628906 635176
rect 208006 633070 208012 633122
rect 208064 633112 208070 633122
rect 208224 633112 208230 633120
rect 208064 633074 208230 633112
rect 208064 633070 208070 633074
rect 208224 633068 208230 633074
rect 208282 633068 208288 633120
rect 230298 632880 230304 632932
rect 230356 632920 230362 632932
rect 241338 632920 241344 632932
rect 230356 632892 241344 632920
rect 230356 632880 230362 632892
rect 241338 632880 241344 632892
rect 241396 632880 241402 632932
rect 621482 632404 621488 632456
rect 621540 632444 621546 632456
rect 641906 632444 641912 632456
rect 621540 632416 641912 632444
rect 621540 632404 621546 632416
rect 641906 632404 641912 632416
rect 641964 632404 641970 632456
rect 208218 632200 208224 632252
rect 208276 632200 208282 632252
rect 208236 632104 208264 632200
rect 208310 632132 208316 632184
rect 208368 632172 208374 632184
rect 208586 632172 208592 632184
rect 208368 632144 208592 632172
rect 208368 632132 208374 632144
rect 208586 632132 208592 632144
rect 208644 632132 208650 632184
rect 208494 632104 208500 632116
rect 208236 632076 208500 632104
rect 208494 632064 208500 632076
rect 208552 632064 208558 632116
rect 208034 631996 208040 632048
rect 208092 632036 208098 632048
rect 208586 632036 208592 632048
rect 208092 632008 208592 632036
rect 208092 631996 208098 632008
rect 208586 631996 208592 632008
rect 208644 631996 208650 632048
rect 208402 631928 208408 631980
rect 208460 631968 208466 631980
rect 208770 631968 208776 631980
rect 208460 631940 208776 631968
rect 208460 631928 208466 631940
rect 208770 631928 208776 631940
rect 208828 631928 208834 631980
rect 208770 631792 208776 631844
rect 208828 631832 208834 631844
rect 208954 631832 208960 631844
rect 208828 631804 208960 631832
rect 208828 631792 208834 631804
rect 208954 631792 208960 631804
rect 209012 631792 209018 631844
rect 675854 631724 675860 631776
rect 675912 631764 675918 631776
rect 676314 631764 676320 631776
rect 675912 631736 676320 631764
rect 675912 631724 675918 631736
rect 676314 631724 676320 631736
rect 676372 631724 676378 631776
rect 676314 631588 676320 631640
rect 676372 631628 676378 631640
rect 676682 631628 676688 631640
rect 676372 631600 676688 631628
rect 676372 631588 676378 631600
rect 676682 631588 676688 631600
rect 676740 631588 676746 631640
rect 676498 631452 676504 631504
rect 676556 631492 676562 631504
rect 676682 631492 676688 631504
rect 676556 631464 676688 631492
rect 676556 631452 676562 631464
rect 676682 631452 676688 631464
rect 676740 631452 676746 631504
rect 208126 631044 208132 631096
rect 208184 631084 208190 631096
rect 208954 631084 208960 631096
rect 208184 631056 208960 631084
rect 208184 631044 208190 631056
rect 208954 631044 208960 631056
rect 209012 631044 209018 631096
rect 208034 630772 208040 630824
rect 208092 630812 208098 630824
rect 208678 630812 208684 630824
rect 208092 630784 208684 630812
rect 208092 630772 208098 630784
rect 208678 630772 208684 630784
rect 208736 630772 208742 630824
rect 641906 630704 641912 630756
rect 641964 630744 641970 630756
rect 652026 630744 652032 630756
rect 641964 630716 652032 630744
rect 641964 630704 641970 630716
rect 652026 630704 652032 630716
rect 652084 630704 652090 630756
rect 208034 630024 208040 630076
rect 208092 630064 208098 630076
rect 208310 630064 208316 630076
rect 208092 630036 208316 630064
rect 208092 630024 208098 630036
rect 208310 630024 208316 630036
rect 208368 630064 208374 630076
rect 209138 630064 209144 630076
rect 208368 630036 209144 630064
rect 208368 630024 208374 630036
rect 209138 630024 209144 630036
rect 209196 630024 209202 630076
rect 208034 629276 208040 629328
rect 208092 629316 208098 629328
rect 208092 629288 208172 629316
rect 208092 629276 208098 629288
rect 208144 629124 208172 629288
rect 208126 629072 208132 629124
rect 208184 629112 208190 629124
rect 208770 629112 208776 629124
rect 208184 629084 208776 629112
rect 208184 629072 208190 629084
rect 208770 629072 208776 629084
rect 208828 629072 208834 629124
rect 208034 628800 208040 628852
rect 208092 628840 208098 628852
rect 208586 628840 208592 628852
rect 208092 628812 208592 628840
rect 208092 628800 208098 628812
rect 208586 628800 208592 628812
rect 208644 628800 208650 628852
rect 675762 628732 675768 628784
rect 675820 628772 675826 628784
rect 676314 628772 676320 628784
rect 675820 628744 676320 628772
rect 675820 628732 675826 628744
rect 676314 628732 676320 628744
rect 676372 628732 676378 628784
rect 675670 628664 675676 628716
rect 675728 628704 675734 628716
rect 676222 628704 676228 628716
rect 675728 628676 676228 628704
rect 675728 628664 675734 628676
rect 676222 628664 676228 628676
rect 676280 628664 676286 628716
rect 208402 628528 208408 628580
rect 208460 628568 208466 628580
rect 208678 628568 208684 628580
rect 208460 628540 208684 628568
rect 208460 628528 208466 628540
rect 208678 628528 208684 628540
rect 208736 628528 208742 628580
rect 676222 628528 676228 628580
rect 676280 628568 676286 628580
rect 676682 628568 676688 628580
rect 676280 628540 676688 628568
rect 676280 628528 676286 628540
rect 676682 628528 676688 628540
rect 676740 628528 676746 628580
rect 645494 626284 645500 626336
rect 645552 626324 645558 626336
rect 661962 626324 661968 626336
rect 645552 626296 661968 626324
rect 645552 626284 645558 626296
rect 661962 626284 661968 626296
rect 662020 626284 662026 626336
rect 228090 626012 228096 626064
rect 228148 626052 228154 626064
rect 230298 626052 230304 626064
rect 228148 626024 230304 626052
rect 228148 626012 228154 626024
rect 230298 626012 230304 626024
rect 230356 626012 230362 626064
rect 208126 625740 208132 625792
rect 208184 625740 208190 625792
rect 208144 625656 208172 625740
rect 208126 625604 208132 625656
rect 208184 625604 208190 625656
rect 619090 624516 619096 624568
rect 619148 624516 619154 624568
rect 208402 624108 208408 624160
rect 208460 624108 208466 624160
rect 208034 623904 208040 623956
rect 208092 623904 208098 623956
rect 208218 623904 208224 623956
rect 208276 623944 208282 623956
rect 208420 623944 208448 624108
rect 208276 623916 208448 623944
rect 208276 623904 208282 623916
rect 208052 623876 208080 623904
rect 208402 623876 208408 623888
rect 208052 623848 208408 623876
rect 208402 623836 208408 623848
rect 208460 623836 208466 623888
rect 208310 623768 208316 623820
rect 208368 623808 208374 623820
rect 208678 623808 208684 623820
rect 208368 623780 208684 623808
rect 208368 623768 208374 623780
rect 208678 623768 208684 623780
rect 208736 623768 208742 623820
rect 208034 623632 208040 623684
rect 208092 623672 208098 623684
rect 208862 623672 208868 623684
rect 208092 623644 208868 623672
rect 208092 623632 208098 623644
rect 208862 623632 208868 623644
rect 208920 623632 208926 623684
rect 619108 621236 619136 624516
rect 675578 622340 675584 622392
rect 675636 622380 675642 622392
rect 676498 622380 676504 622392
rect 675636 622352 676504 622380
rect 675636 622340 675642 622352
rect 676498 622340 676504 622352
rect 676556 622340 676562 622392
rect 675302 621320 675308 621372
rect 675360 621360 675366 621372
rect 675854 621360 675860 621372
rect 675360 621332 675860 621360
rect 675360 621320 675366 621332
rect 675854 621320 675860 621332
rect 675912 621320 675918 621372
rect 619090 621184 619096 621236
rect 619148 621184 619154 621236
rect 675854 621184 675860 621236
rect 675912 621224 675918 621236
rect 676222 621224 676228 621236
rect 675912 621196 676228 621224
rect 675912 621184 675918 621196
rect 676222 621184 676228 621196
rect 676280 621184 676286 621236
rect 675670 620980 675676 621032
rect 675728 621020 675734 621032
rect 676314 621020 676320 621032
rect 675728 620992 676320 621020
rect 675728 620980 675734 620992
rect 676314 620980 676320 620992
rect 676372 620980 676378 621032
rect 675854 619484 675860 619536
rect 675912 619524 675918 619536
rect 676314 619524 676320 619536
rect 675912 619496 676320 619524
rect 675912 619484 675918 619496
rect 676314 619484 676320 619496
rect 676372 619484 676378 619536
rect 619090 619212 619096 619264
rect 619148 619252 619154 619264
rect 620010 619252 620016 619264
rect 619148 619224 620016 619252
rect 619148 619212 619154 619224
rect 620010 619212 620016 619224
rect 620068 619212 620074 619264
rect 619090 617376 619096 617428
rect 619148 617416 619154 617428
rect 620010 617416 620016 617428
rect 619148 617388 620016 617416
rect 619148 617376 619154 617388
rect 620010 617376 620016 617388
rect 620068 617376 620074 617428
rect 620010 617172 620016 617224
rect 620068 617212 620074 617224
rect 620654 617212 620660 617224
rect 620068 617184 620660 617212
rect 620068 617172 620074 617184
rect 620654 617172 620660 617184
rect 620712 617172 620718 617224
rect 643194 616968 643200 617020
rect 643252 617008 643258 617020
rect 676314 617008 676320 617020
rect 643252 616980 676320 617008
rect 643252 616968 643258 616980
rect 676314 616968 676320 616980
rect 676372 616968 676378 617020
rect 676222 616424 676228 616476
rect 676280 616424 676286 616476
rect 676240 616260 676268 616424
rect 676314 616260 676320 616272
rect 676240 616232 676320 616260
rect 676314 616220 676320 616232
rect 676372 616220 676378 616272
rect 675578 616084 675584 616136
rect 675636 616084 675642 616136
rect 675486 615880 675492 615932
rect 675544 615920 675550 615932
rect 675596 615920 675624 616084
rect 675544 615892 675624 615920
rect 675544 615880 675550 615892
rect 625530 615812 625536 615864
rect 625588 615852 625594 615864
rect 675762 615852 675768 615864
rect 625588 615824 675768 615852
rect 625588 615812 625594 615824
rect 675762 615812 675768 615824
rect 675820 615852 675826 615864
rect 676222 615852 676228 615864
rect 675820 615824 676228 615852
rect 675820 615812 675826 615824
rect 676222 615812 676228 615824
rect 676280 615812 676286 615864
rect 676314 615812 676320 615864
rect 676372 615812 676378 615864
rect 675394 615744 675400 615796
rect 675452 615784 675458 615796
rect 676332 615784 676360 615812
rect 675452 615756 676360 615784
rect 675452 615744 675458 615756
rect 675486 615676 675492 615728
rect 675544 615716 675550 615728
rect 676222 615716 676228 615728
rect 675544 615688 676228 615716
rect 675544 615676 675550 615688
rect 676222 615676 676228 615688
rect 676280 615676 676286 615728
rect 652026 615608 652032 615660
rect 652084 615648 652090 615660
rect 654234 615648 654240 615660
rect 652084 615620 654240 615648
rect 652084 615608 652090 615620
rect 654234 615608 654240 615620
rect 654292 615608 654298 615660
rect 675854 614928 675860 614980
rect 675912 614968 675918 614980
rect 676222 614968 676228 614980
rect 675912 614940 676228 614968
rect 675912 614928 675918 614940
rect 676222 614928 676228 614940
rect 676280 614928 676286 614980
rect 675302 614248 675308 614300
rect 675360 614288 675366 614300
rect 676314 614288 676320 614300
rect 675360 614260 676320 614288
rect 675360 614248 675366 614260
rect 676314 614248 676320 614260
rect 676372 614248 676378 614300
rect 213738 614112 213744 614164
rect 213796 614152 213802 614164
rect 228090 614152 228096 614164
rect 213796 614124 228096 614152
rect 213796 614112 213802 614124
rect 228090 614112 228096 614124
rect 228148 614112 228154 614164
rect 675394 613500 675400 613552
rect 675452 613540 675458 613552
rect 675670 613540 675676 613552
rect 675452 613512 675676 613540
rect 675452 613500 675458 613512
rect 675670 613500 675676 613512
rect 675728 613540 675734 613552
rect 676222 613540 676228 613552
rect 675728 613512 676228 613540
rect 675728 613500 675734 613512
rect 676222 613500 676228 613512
rect 676280 613500 676286 613552
rect 619458 613200 619464 613212
rect 619016 613172 619464 613200
rect 619016 612928 619044 613172
rect 619458 613160 619464 613172
rect 619516 613160 619522 613212
rect 675578 613092 675584 613144
rect 675636 613132 675642 613144
rect 676314 613132 676320 613144
rect 675636 613104 676320 613132
rect 675636 613092 675642 613104
rect 676314 613092 676320 613104
rect 676372 613092 676378 613144
rect 619090 613024 619096 613076
rect 619148 613064 619154 613076
rect 619458 613064 619464 613076
rect 619148 613036 619464 613064
rect 619148 613024 619154 613036
rect 619458 613024 619464 613036
rect 619516 613024 619522 613076
rect 619090 612928 619096 612940
rect 619016 612900 619096 612928
rect 619090 612888 619096 612900
rect 619148 612888 619154 612940
rect 675670 612208 675676 612260
rect 675728 612248 675734 612260
rect 676222 612248 676228 612260
rect 675728 612220 676228 612248
rect 675728 612208 675734 612220
rect 676222 612208 676228 612220
rect 676280 612208 676286 612260
rect 675854 611936 675860 611988
rect 675912 611976 675918 611988
rect 676314 611976 676320 611988
rect 675912 611948 676320 611976
rect 675912 611936 675918 611948
rect 676314 611936 676320 611948
rect 676372 611936 676378 611988
rect 207942 611800 207948 611852
rect 208000 611840 208006 611852
rect 208678 611840 208684 611852
rect 208000 611812 208684 611840
rect 208000 611800 208006 611812
rect 208678 611800 208684 611812
rect 208736 611800 208742 611852
rect 208494 611732 208500 611784
rect 208552 611772 208558 611784
rect 217050 611772 217056 611784
rect 208552 611744 217056 611772
rect 208552 611732 208558 611744
rect 217050 611732 217056 611744
rect 217108 611732 217114 611784
rect 208402 611638 208408 611690
rect 208460 611638 208466 611690
rect 208420 611244 208448 611638
rect 624426 611460 624432 611512
rect 624484 611500 624490 611512
rect 676222 611500 676228 611512
rect 624484 611472 676228 611500
rect 624484 611460 624490 611472
rect 676222 611460 676228 611472
rect 676280 611460 676286 611512
rect 675486 611324 675492 611376
rect 675544 611364 675550 611376
rect 676222 611364 676228 611376
rect 675544 611336 676228 611364
rect 675544 611324 675550 611336
rect 676222 611324 676228 611336
rect 676280 611324 676286 611376
rect 208494 611244 208500 611256
rect 208043 611177 208049 611229
rect 208101 611217 208107 611229
rect 208382 611217 208500 611244
rect 208101 611216 208500 611217
rect 208101 611189 208410 611216
rect 208494 611204 208500 611216
rect 208552 611204 208558 611256
rect 208101 611177 208107 611189
rect 209506 610848 209512 610900
rect 209564 610888 209570 610900
rect 213738 610888 213744 610900
rect 209564 610860 213744 610888
rect 209564 610848 209570 610860
rect 213738 610848 213744 610860
rect 213796 610848 213802 610900
rect 619090 610576 619096 610628
rect 619148 610616 619154 610628
rect 619458 610616 619464 610628
rect 619148 610588 619464 610616
rect 619148 610576 619154 610588
rect 619458 610576 619464 610588
rect 619516 610576 619522 610628
rect 675302 609556 675308 609608
rect 675360 609596 675366 609608
rect 675360 609568 676437 609596
rect 675360 609556 675366 609568
rect 208034 609148 208040 609200
rect 208092 609188 208098 609200
rect 209782 609188 209788 609200
rect 208092 609160 209788 609188
rect 208092 609148 208098 609160
rect 209782 609148 209788 609160
rect 209840 609148 209846 609200
rect 675854 609080 675860 609132
rect 675912 609120 675918 609132
rect 676314 609120 676320 609132
rect 675912 609092 676320 609120
rect 675912 609080 675918 609092
rect 676314 609080 676320 609092
rect 676372 609080 676378 609132
rect 675486 609012 675492 609064
rect 675544 609052 675550 609064
rect 675946 609052 675952 609064
rect 675544 609024 675952 609052
rect 675544 609012 675550 609024
rect 675946 609012 675952 609024
rect 676004 609012 676010 609064
rect 675762 608944 675768 608996
rect 675820 608984 675826 608996
rect 676314 608984 676320 608996
rect 675820 608956 676320 608984
rect 675820 608944 675826 608956
rect 676314 608944 676320 608956
rect 676372 608944 676378 608996
rect 208126 608536 208132 608588
rect 208184 608576 208190 608588
rect 208770 608576 208776 608588
rect 208184 608548 208776 608576
rect 208184 608536 208190 608548
rect 208770 608536 208776 608548
rect 208828 608536 208834 608588
rect 208218 608236 208224 608248
rect 207962 608208 208224 608236
rect 208218 608196 208224 608208
rect 208276 608236 208282 608248
rect 208494 608236 208500 608248
rect 208276 608208 208500 608236
rect 208276 608196 208282 608208
rect 208494 608196 208500 608208
rect 208552 608196 208558 608248
rect 675762 608128 675768 608180
rect 675820 608168 675826 608180
rect 676222 608168 676228 608180
rect 675820 608140 676228 608168
rect 675820 608128 675826 608140
rect 676222 608128 676228 608140
rect 676280 608128 676286 608180
rect 675302 606564 675308 606616
rect 675360 606604 675366 606616
rect 676314 606604 676320 606616
rect 675360 606576 676320 606604
rect 675360 606564 675366 606576
rect 676314 606564 676320 606576
rect 676372 606564 676378 606616
rect 675394 606156 675400 606208
rect 675452 606196 675458 606208
rect 676314 606196 676320 606208
rect 675452 606168 676320 606196
rect 675452 606156 675458 606168
rect 676314 606156 676320 606168
rect 676372 606156 676378 606208
rect 233610 605884 233616 605936
rect 233668 605924 233674 605936
rect 252378 605924 252384 605936
rect 233668 605896 252384 605924
rect 233668 605884 233674 605896
rect 252378 605884 252384 605896
rect 252436 605884 252442 605936
rect 625530 605884 625536 605936
rect 625588 605924 625594 605936
rect 669690 605924 669696 605936
rect 625588 605896 669696 605924
rect 625588 605884 625594 605896
rect 669690 605884 669696 605896
rect 669748 605884 669754 605936
rect 675578 605816 675584 605868
rect 675636 605856 675642 605868
rect 676314 605856 676320 605868
rect 675636 605828 676320 605856
rect 675636 605816 675642 605828
rect 676314 605816 676320 605828
rect 676372 605816 676378 605868
rect 643286 605340 643292 605392
rect 643344 605380 643350 605392
rect 645494 605380 645500 605392
rect 643344 605352 645500 605380
rect 643344 605340 643350 605352
rect 645494 605340 645500 605352
rect 645552 605340 645558 605392
rect 675854 605340 675860 605392
rect 675912 605380 675918 605392
rect 676498 605380 676504 605392
rect 675912 605352 676504 605380
rect 675912 605340 675918 605352
rect 676498 605340 676504 605352
rect 676556 605340 676562 605392
rect 675670 605272 675676 605324
rect 675728 605312 675734 605324
rect 676590 605312 676596 605324
rect 675728 605284 676596 605312
rect 675728 605272 675734 605284
rect 676590 605272 676596 605284
rect 676648 605272 676654 605324
rect 675302 605204 675308 605256
rect 675360 605244 675366 605256
rect 675854 605244 675860 605256
rect 675360 605216 675860 605244
rect 675360 605204 675366 605216
rect 675854 605204 675860 605216
rect 675912 605204 675918 605256
rect 675486 605136 675492 605188
rect 675544 605176 675550 605188
rect 675946 605176 675952 605188
rect 675544 605148 675952 605176
rect 675544 605136 675550 605148
rect 675946 605136 675952 605148
rect 676004 605136 676010 605188
rect 675762 605068 675768 605120
rect 675820 605108 675826 605120
rect 676222 605108 676228 605120
rect 675820 605080 676228 605108
rect 675820 605068 675826 605080
rect 676222 605068 676228 605080
rect 676280 605068 676286 605120
rect 208402 605000 208408 605052
rect 208460 605000 208466 605052
rect 208420 604780 208448 605000
rect 208402 604728 208408 604780
rect 208460 604728 208466 604780
rect 208034 603232 208040 603284
rect 208092 603272 208098 603284
rect 208586 603272 208592 603284
rect 208092 603244 208592 603272
rect 208092 603232 208098 603244
rect 208586 603232 208592 603244
rect 208644 603232 208650 603284
rect 654234 602008 654240 602060
rect 654292 602048 654298 602060
rect 659754 602048 659760 602060
rect 654292 602020 659760 602048
rect 654292 602008 654298 602020
rect 659754 602008 659760 602020
rect 659812 602008 659818 602060
rect 208034 601396 208040 601448
rect 208092 601436 208098 601448
rect 208310 601436 208316 601448
rect 208092 601408 208316 601436
rect 208092 601396 208098 601408
rect 208310 601396 208316 601408
rect 208368 601436 208374 601448
rect 209322 601436 209328 601448
rect 208368 601408 209328 601436
rect 208368 601396 208374 601408
rect 209322 601396 209328 601408
rect 209380 601396 209386 601448
rect 639882 601396 639888 601448
rect 639940 601436 639946 601448
rect 643286 601436 643292 601448
rect 639940 601408 643292 601436
rect 639940 601396 639946 601408
rect 643286 601396 643292 601408
rect 643344 601396 643350 601448
rect 211530 599288 211536 599340
rect 211588 599328 211594 599340
rect 244650 599328 244656 599340
rect 211588 599300 244656 599328
rect 211588 599288 211594 599300
rect 244650 599288 244656 599300
rect 244708 599288 244714 599340
rect 208126 598948 208132 599000
rect 208184 598988 208190 599000
rect 208770 598988 208776 599000
rect 208184 598960 208776 598988
rect 208184 598948 208190 598960
rect 208770 598948 208776 598960
rect 208828 598948 208834 599000
rect 208034 598812 208040 598864
rect 208092 598852 208098 598864
rect 208770 598852 208776 598864
rect 208092 598824 208776 598852
rect 208092 598812 208098 598824
rect 208770 598812 208776 598824
rect 208828 598812 208834 598864
rect 208034 597792 208040 597844
rect 208092 597832 208098 597844
rect 208494 597832 208500 597844
rect 208092 597804 208500 597832
rect 208092 597792 208098 597804
rect 208494 597792 208500 597804
rect 208552 597832 208558 597844
rect 208678 597832 208684 597844
rect 208552 597804 208684 597832
rect 208552 597792 208558 597804
rect 208678 597792 208684 597804
rect 208736 597792 208742 597844
rect 208034 596772 208040 596824
rect 208092 596812 208098 596824
rect 208770 596812 208776 596824
rect 208092 596784 208776 596812
rect 208092 596772 208098 596784
rect 208770 596772 208776 596784
rect 208828 596772 208834 596824
rect 208218 595072 208224 595124
rect 208276 595112 208282 595124
rect 208586 595112 208592 595124
rect 208276 595084 208592 595112
rect 208276 595072 208282 595084
rect 208586 595072 208592 595084
rect 208644 595072 208650 595124
rect 209782 590448 209788 590500
rect 209840 590488 209846 590500
rect 219350 590488 219356 590500
rect 209840 590460 219356 590488
rect 209840 590448 209846 590460
rect 219350 590448 219356 590460
rect 219408 590448 219414 590500
rect 659754 587660 659760 587712
rect 659812 587700 659818 587712
rect 667482 587700 667488 587712
rect 659812 587672 667488 587700
rect 659812 587660 659818 587672
rect 667482 587660 667488 587672
rect 667540 587660 667546 587712
rect 637766 587184 637772 587236
rect 637824 587224 637830 587236
rect 639882 587224 639888 587236
rect 637824 587196 639888 587224
rect 637824 587184 637830 587196
rect 639882 587184 639888 587196
rect 639940 587184 639946 587236
rect 208402 585484 208408 585536
rect 208460 585524 208466 585536
rect 249066 585524 249072 585536
rect 208460 585496 249072 585524
rect 208460 585484 208466 585496
rect 249066 585484 249072 585496
rect 249124 585484 249130 585536
rect 208126 585416 208132 585468
rect 208184 585456 208190 585468
rect 252378 585456 252384 585468
rect 208184 585428 252384 585456
rect 208184 585416 208190 585428
rect 252378 585416 252384 585428
rect 252436 585416 252442 585468
rect 208034 583852 208040 583904
rect 208092 583892 208098 583904
rect 208770 583892 208776 583904
rect 208092 583864 208776 583892
rect 208092 583852 208098 583864
rect 208770 583852 208776 583864
rect 208828 583852 208834 583904
rect 209690 583852 209696 583904
rect 209748 583892 209754 583904
rect 249158 583892 249164 583904
rect 209748 583864 249164 583892
rect 209748 583852 209754 583864
rect 249158 583852 249164 583864
rect 249216 583852 249222 583904
rect 676314 582220 676320 582272
rect 676372 582220 676378 582272
rect 676332 582124 676360 582220
rect 675780 582096 676360 582124
rect 675780 582068 675808 582096
rect 675762 582016 675768 582068
rect 675820 582016 675826 582068
rect 635558 581880 635564 581932
rect 635616 581920 635622 581932
rect 637766 581920 637772 581932
rect 635616 581892 637772 581920
rect 635616 581880 635622 581892
rect 637766 581880 637772 581892
rect 637824 581880 637830 581932
rect 208034 581744 208040 581796
rect 208092 581784 208098 581796
rect 208494 581784 208500 581796
rect 208092 581756 208500 581784
rect 208092 581744 208098 581756
rect 208494 581744 208500 581756
rect 208552 581744 208558 581796
rect 675578 581404 675584 581456
rect 675636 581444 675642 581456
rect 676498 581444 676504 581456
rect 675636 581416 676504 581444
rect 675636 581404 675642 581416
rect 676498 581404 676504 581416
rect 676556 581404 676562 581456
rect 624426 581336 624432 581388
rect 624484 581376 624490 581388
rect 673370 581376 673376 581388
rect 624484 581348 673376 581376
rect 624484 581336 624490 581348
rect 673370 581336 673376 581348
rect 673428 581336 673434 581388
rect 208862 580832 208868 580844
rect 207962 580804 208868 580832
rect 208862 580792 208868 580804
rect 208920 580792 208926 580844
rect 676314 580628 676320 580640
rect 673618 580600 676320 580628
rect 673370 580520 673376 580572
rect 673428 580560 673434 580572
rect 673618 580560 673646 580600
rect 676314 580588 676320 580600
rect 676372 580588 676378 580640
rect 673428 580532 673646 580560
rect 673428 580520 673434 580532
rect 676314 580180 676320 580232
rect 676372 580180 676378 580232
rect 676332 580096 676360 580180
rect 675394 580044 675400 580096
rect 675452 580084 675458 580096
rect 675854 580084 675860 580096
rect 675452 580056 675860 580084
rect 675452 580044 675458 580056
rect 675854 580044 675860 580056
rect 675912 580084 675918 580096
rect 676314 580084 676320 580096
rect 675912 580056 676320 580084
rect 675912 580044 675918 580056
rect 676314 580044 676320 580056
rect 676372 580044 676378 580096
rect 208310 578820 208316 578872
rect 208368 578860 208374 578872
rect 208586 578860 208592 578872
rect 208368 578832 208592 578860
rect 208368 578820 208374 578832
rect 208586 578820 208592 578832
rect 208644 578820 208650 578872
rect 675670 578820 675676 578872
rect 675728 578860 675734 578872
rect 676222 578860 676228 578872
rect 675728 578832 676228 578860
rect 675728 578820 675734 578832
rect 676222 578820 676228 578832
rect 676280 578820 676286 578872
rect 675578 578684 675584 578736
rect 675636 578724 675642 578736
rect 676222 578724 676228 578736
rect 675636 578696 676228 578724
rect 675636 578684 675642 578696
rect 676222 578684 676228 578696
rect 676280 578684 676286 578736
rect 208034 578344 208040 578396
rect 208092 578384 208098 578396
rect 208678 578384 208684 578396
rect 208092 578356 208684 578384
rect 208092 578344 208098 578356
rect 208678 578344 208684 578356
rect 208736 578344 208742 578396
rect 675394 578208 675400 578260
rect 675452 578248 675458 578260
rect 676222 578248 676228 578260
rect 675452 578220 676228 578248
rect 675452 578208 675458 578220
rect 676222 578208 676228 578220
rect 676280 578208 676286 578260
rect 675486 578140 675492 578192
rect 675544 578180 675550 578192
rect 675946 578180 675952 578192
rect 675544 578152 675952 578180
rect 675544 578140 675550 578152
rect 675946 578140 675952 578152
rect 676004 578140 676010 578192
rect 676130 578072 676136 578124
rect 676188 578072 676194 578124
rect 676148 577988 676176 578072
rect 676130 577936 676136 577988
rect 676188 577936 676194 577988
rect 208218 577460 208224 577512
rect 208276 577460 208282 577512
rect 208236 577172 208264 577460
rect 208218 577120 208224 577172
rect 208276 577120 208282 577172
rect 219350 576848 219356 576900
rect 219408 576888 219414 576900
rect 221558 576888 221564 576900
rect 219408 576860 221564 576888
rect 219408 576848 219414 576860
rect 221558 576848 221564 576860
rect 221616 576848 221622 576900
rect 676314 576100 676320 576152
rect 676372 576100 676378 576152
rect 676130 576032 676136 576084
rect 676188 576032 676194 576084
rect 676148 575948 676176 576032
rect 676130 575896 676136 575948
rect 676188 575896 676194 575948
rect 675670 575760 675676 575812
rect 675728 575800 675734 575812
rect 675946 575800 675952 575812
rect 675728 575772 675952 575800
rect 675728 575760 675734 575772
rect 675946 575760 675952 575772
rect 676004 575760 676010 575812
rect 675854 575692 675860 575744
rect 675912 575732 675918 575744
rect 676222 575732 676228 575744
rect 675912 575704 676228 575732
rect 675912 575692 675918 575704
rect 676222 575692 676228 575704
rect 676280 575692 676286 575744
rect 675486 575556 675492 575608
rect 675544 575596 675550 575608
rect 676222 575596 676228 575608
rect 675544 575568 676228 575596
rect 675544 575556 675550 575568
rect 676222 575556 676228 575568
rect 676280 575556 676286 575608
rect 676222 575420 676228 575472
rect 676280 575460 676286 575472
rect 676332 575460 676360 576100
rect 676280 575432 676360 575460
rect 676280 575420 676286 575432
rect 208034 575216 208040 575268
rect 208092 575256 208098 575268
rect 208494 575256 208500 575268
rect 208092 575228 208500 575256
rect 208092 575216 208098 575228
rect 208494 575216 208500 575228
rect 208552 575216 208558 575268
rect 208310 575148 208316 575200
rect 208368 575188 208374 575200
rect 208770 575188 208776 575200
rect 208368 575160 208776 575188
rect 208368 575148 208374 575160
rect 208770 575148 208776 575160
rect 208828 575148 208834 575200
rect 675854 575080 675860 575132
rect 675912 575120 675918 575132
rect 676314 575120 676320 575132
rect 675912 575092 676320 575120
rect 675912 575080 675918 575092
rect 676314 575080 676320 575092
rect 676372 575080 676378 575132
rect 208034 574944 208040 574996
rect 208092 574984 208098 574996
rect 208770 574984 208776 574996
rect 208092 574956 208776 574984
rect 208092 574944 208098 574956
rect 208770 574944 208776 574956
rect 208828 574944 208834 574996
rect 675302 574944 675308 574996
rect 675360 574984 675366 574996
rect 675670 574984 675676 574996
rect 675360 574956 675676 574984
rect 675360 574944 675366 574956
rect 675670 574944 675676 574956
rect 675728 574944 675734 574996
rect 676038 574944 676044 574996
rect 676096 574944 676102 574996
rect 676130 574944 676136 574996
rect 676188 574944 676194 574996
rect 208678 574876 208684 574928
rect 208736 574916 208742 574928
rect 208862 574916 208868 574928
rect 208736 574888 208868 574916
rect 208736 574876 208742 574888
rect 208862 574876 208868 574888
rect 208920 574876 208926 574928
rect 675762 574876 675768 574928
rect 675820 574876 675826 574928
rect 675670 574808 675676 574860
rect 675728 574848 675734 574860
rect 675780 574848 675808 574876
rect 676056 574860 676084 574944
rect 676148 574860 676176 574944
rect 675728 574820 675808 574848
rect 675728 574808 675734 574820
rect 676038 574808 676044 574860
rect 676096 574808 676102 574860
rect 676130 574808 676136 574860
rect 676188 574808 676194 574860
rect 208218 574740 208224 574792
rect 208276 574780 208282 574792
rect 208678 574780 208684 574792
rect 208276 574752 208684 574780
rect 208276 574740 208282 574752
rect 208678 574740 208684 574752
rect 208736 574740 208742 574792
rect 675946 574740 675952 574792
rect 676004 574780 676010 574792
rect 676314 574780 676320 574792
rect 676004 574752 676320 574780
rect 676004 574740 676010 574752
rect 676314 574740 676320 574752
rect 676372 574740 676378 574792
rect 208310 574536 208316 574588
rect 208368 574576 208374 574588
rect 208494 574576 208500 574588
rect 208368 574548 208500 574576
rect 208368 574536 208374 574548
rect 208494 574536 208500 574548
rect 208552 574536 208558 574588
rect 675302 574128 675308 574180
rect 675360 574168 675366 574180
rect 676314 574168 676320 574180
rect 675360 574140 676320 574168
rect 675360 574128 675366 574140
rect 676314 574128 676320 574140
rect 676372 574128 676378 574180
rect 208034 573584 208040 573636
rect 208092 573624 208098 573636
rect 208862 573624 208868 573636
rect 208092 573596 208868 573624
rect 208092 573584 208098 573596
rect 208862 573584 208868 573596
rect 208920 573584 208926 573636
rect 675486 573584 675492 573636
rect 675544 573624 675550 573636
rect 676314 573624 676320 573636
rect 675544 573596 676320 573624
rect 675544 573584 675550 573596
rect 676314 573584 676320 573596
rect 676372 573584 676378 573636
rect 674106 572292 674112 572344
rect 674164 572332 674170 572344
rect 676222 572332 676228 572344
rect 674164 572304 676228 572332
rect 674164 572292 674170 572304
rect 676222 572292 676228 572304
rect 676280 572292 676286 572344
rect 208218 571748 208224 571800
rect 208276 571788 208282 571800
rect 208494 571788 208500 571800
rect 208276 571760 208500 571788
rect 208276 571748 208282 571760
rect 208494 571748 208500 571760
rect 208552 571748 208558 571800
rect 208126 571612 208132 571664
rect 208184 571652 208190 571664
rect 208494 571652 208500 571664
rect 208184 571624 208500 571652
rect 208184 571612 208190 571624
rect 208494 571612 208500 571624
rect 208552 571612 208558 571664
rect 675854 571476 675860 571528
rect 675912 571516 675918 571528
rect 676222 571516 676228 571528
rect 675912 571488 676228 571516
rect 675912 571476 675918 571488
rect 676222 571476 676228 571488
rect 676280 571476 676286 571528
rect 675578 571136 675584 571188
rect 675636 571176 675642 571188
rect 676314 571176 676320 571188
rect 675636 571148 676320 571176
rect 675636 571136 675642 571148
rect 676314 571136 676320 571148
rect 676372 571136 676378 571188
rect 675578 571000 675584 571052
rect 675636 571040 675642 571052
rect 675946 571040 675952 571052
rect 675636 571012 675952 571040
rect 675636 571000 675642 571012
rect 675946 571000 675952 571012
rect 676004 571000 676010 571052
rect 208218 570728 208224 570780
rect 208276 570768 208282 570780
rect 208678 570768 208684 570780
rect 208276 570740 208684 570768
rect 208276 570728 208282 570740
rect 208678 570728 208684 570740
rect 208736 570728 208742 570780
rect 667482 570592 667488 570644
rect 667540 570632 667546 570644
rect 676222 570632 676228 570644
rect 667540 570604 676228 570632
rect 667540 570592 667546 570604
rect 676222 570592 676228 570604
rect 676280 570592 676286 570644
rect 208034 569164 208040 569216
rect 208092 569204 208098 569216
rect 208678 569204 208684 569216
rect 208092 569176 208684 569204
rect 208092 569164 208098 569176
rect 208678 569164 208684 569176
rect 208736 569204 208742 569216
rect 208862 569204 208868 569216
rect 208736 569176 208868 569204
rect 208736 569164 208742 569176
rect 208862 569164 208868 569176
rect 208920 569164 208926 569216
rect 208126 569096 208132 569148
rect 208184 569136 208190 569148
rect 208586 569136 208592 569148
rect 208184 569108 208592 569136
rect 208184 569096 208190 569108
rect 208586 569096 208592 569108
rect 208644 569096 208650 569148
rect 208034 568756 208040 568808
rect 208092 568796 208098 568808
rect 208770 568796 208776 568808
rect 208092 568768 208776 568796
rect 208092 568756 208098 568768
rect 208770 568756 208776 568768
rect 208828 568756 208834 568808
rect 675394 568756 675400 568808
rect 675452 568796 675458 568808
rect 675946 568796 675952 568808
rect 675452 568768 675952 568796
rect 675452 568756 675458 568768
rect 675946 568756 675952 568768
rect 676004 568796 676010 568808
rect 676004 568768 676437 568796
rect 676004 568756 676010 568768
rect 619274 568416 619280 568468
rect 619332 568456 619338 568468
rect 629762 568456 629768 568468
rect 619332 568428 629768 568456
rect 619332 568416 619338 568428
rect 629762 568416 629768 568428
rect 629820 568416 629826 568468
rect 623414 568348 623420 568400
rect 623472 568388 623478 568400
rect 635558 568388 635564 568400
rect 623472 568360 635564 568388
rect 623472 568348 623478 568360
rect 635558 568348 635564 568360
rect 635616 568348 635622 568400
rect 675394 567804 675400 567856
rect 675452 567844 675458 567856
rect 675670 567844 675676 567856
rect 675452 567816 675676 567844
rect 675452 567804 675458 567816
rect 675670 567804 675676 567816
rect 675728 567804 675734 567856
rect 208126 567736 208132 567788
rect 208184 567776 208190 567788
rect 221466 567776 221472 567788
rect 208184 567748 221472 567776
rect 208184 567736 208190 567748
rect 221466 567736 221472 567748
rect 221524 567736 221530 567788
rect 675670 567668 675676 567720
rect 675728 567708 675734 567720
rect 675946 567708 675952 567720
rect 675728 567680 675952 567708
rect 675728 567668 675734 567680
rect 675946 567668 675952 567680
rect 676004 567668 676010 567720
rect 208126 566648 208132 566700
rect 208184 566688 208190 566700
rect 209046 566688 209052 566700
rect 208184 566660 209052 566688
rect 208184 566648 208190 566660
rect 209046 566648 209052 566660
rect 209104 566648 209110 566700
rect 629762 566648 629768 566700
rect 629820 566688 629826 566700
rect 645494 566688 645500 566700
rect 629820 566660 645500 566688
rect 629820 566648 629826 566660
rect 645494 566648 645500 566660
rect 645552 566648 645558 566700
rect 675670 565696 675676 565748
rect 675728 565736 675734 565748
rect 676222 565736 676228 565748
rect 675728 565708 676228 565736
rect 675728 565696 675734 565708
rect 676222 565696 676228 565708
rect 676280 565696 676286 565748
rect 221558 565560 221564 565612
rect 221616 565600 221622 565612
rect 225882 565600 225888 565612
rect 221616 565572 225888 565600
rect 221616 565560 221622 565572
rect 225882 565560 225888 565572
rect 225940 565560 225946 565612
rect 675486 565356 675492 565408
rect 675544 565396 675550 565408
rect 676314 565396 676320 565408
rect 675544 565368 676320 565396
rect 675544 565356 675550 565368
rect 676314 565356 676320 565368
rect 676372 565356 676378 565408
rect 675394 565016 675400 565068
rect 675452 565056 675458 565068
rect 676314 565056 676320 565068
rect 675452 565028 676320 565056
rect 675452 565016 675458 565028
rect 676314 565016 676320 565028
rect 676372 565016 676378 565068
rect 675762 564540 675768 564592
rect 675820 564580 675826 564592
rect 676590 564580 676596 564592
rect 675820 564552 676596 564580
rect 675820 564540 675826 564552
rect 676590 564540 676596 564552
rect 676648 564540 676654 564592
rect 675302 563792 675308 563844
rect 675360 563832 675366 563844
rect 676682 563832 676688 563844
rect 675360 563804 676688 563832
rect 675360 563792 675366 563804
rect 676682 563792 676688 563804
rect 676740 563792 676746 563844
rect 675578 563384 675584 563436
rect 675636 563424 675642 563436
rect 676222 563424 676228 563436
rect 675636 563396 676228 563424
rect 675636 563384 675642 563396
rect 676222 563384 676228 563396
rect 676280 563384 676286 563436
rect 645494 561888 645500 561940
rect 645552 561928 645558 561940
rect 649818 561928 649824 561940
rect 645552 561900 649824 561928
rect 645552 561888 645558 561900
rect 649818 561888 649824 561900
rect 649876 561888 649882 561940
rect 676498 558964 676504 559016
rect 676556 559004 676562 559016
rect 676682 559004 676688 559016
rect 676556 558976 676688 559004
rect 676556 558964 676562 558976
rect 676682 558964 676688 558976
rect 676740 558964 676746 559016
rect 664170 558896 664176 558948
rect 664228 558936 664234 558948
rect 670794 558936 670800 558948
rect 664228 558908 670800 558936
rect 664228 558896 664234 558908
rect 670794 558896 670800 558908
rect 670852 558896 670858 558948
rect 676406 558828 676412 558880
rect 676464 558868 676470 558880
rect 676682 558868 676688 558880
rect 676464 558840 676688 558868
rect 676464 558828 676470 558840
rect 676682 558828 676688 558840
rect 676740 558828 676746 558880
rect 208494 557808 208500 557860
rect 208552 557848 208558 557860
rect 251182 557848 251188 557860
rect 208552 557820 251188 557848
rect 208552 557808 208558 557820
rect 251182 557808 251188 557820
rect 251240 557808 251246 557860
rect 208126 557672 208132 557724
rect 208184 557712 208190 557724
rect 208494 557712 208500 557724
rect 208184 557684 208500 557712
rect 208184 557672 208190 557684
rect 208494 557672 208500 557684
rect 208552 557672 208558 557724
rect 208034 556924 208040 556976
rect 208092 556964 208098 556976
rect 208954 556964 208960 556976
rect 208092 556936 208960 556964
rect 208092 556924 208098 556936
rect 208954 556924 208960 556936
rect 209012 556924 209018 556976
rect 208052 556772 208080 556924
rect 225882 556856 225888 556908
rect 225940 556896 225946 556908
rect 234714 556896 234720 556908
rect 225940 556868 234720 556896
rect 225940 556856 225946 556868
rect 234714 556856 234720 556868
rect 234772 556856 234778 556908
rect 208034 556720 208040 556772
rect 208092 556720 208098 556772
rect 208034 556516 208040 556568
rect 208092 556556 208098 556568
rect 208678 556556 208684 556568
rect 208092 556528 208684 556556
rect 208092 556516 208098 556528
rect 208678 556516 208684 556528
rect 208736 556516 208742 556568
rect 208402 556244 208408 556296
rect 208460 556284 208466 556296
rect 244650 556284 244656 556296
rect 208460 556256 244656 556284
rect 208460 556244 208466 556256
rect 244650 556244 244656 556256
rect 244708 556244 244714 556296
rect 619090 554680 619096 554732
rect 619148 554720 619154 554732
rect 619274 554720 619280 554732
rect 619148 554692 619280 554720
rect 619148 554680 619154 554692
rect 619274 554680 619280 554692
rect 619332 554680 619338 554732
rect 208310 554408 208316 554460
rect 208368 554448 208374 554460
rect 208770 554448 208776 554460
rect 208368 554420 208776 554448
rect 208368 554408 208374 554420
rect 208770 554408 208776 554420
rect 208828 554408 208834 554460
rect 208218 554340 208224 554392
rect 208276 554380 208282 554392
rect 208862 554380 208868 554392
rect 208276 554352 208868 554380
rect 208276 554340 208282 554352
rect 208862 554340 208868 554352
rect 208920 554340 208926 554392
rect 208218 553428 208224 553440
rect 207962 553400 208224 553428
rect 208218 553388 208224 553400
rect 208276 553428 208282 553440
rect 208678 553428 208684 553440
rect 208276 553400 208684 553428
rect 208276 553388 208282 553400
rect 208678 553388 208684 553400
rect 208736 553388 208742 553440
rect 208126 552300 208132 552352
rect 208184 552340 208190 552352
rect 208678 552340 208684 552352
rect 208184 552312 208684 552340
rect 208184 552300 208190 552312
rect 208678 552300 208684 552312
rect 208736 552300 208742 552352
rect 208034 550866 208040 550918
rect 208092 550906 208098 550918
rect 208494 550906 208500 550918
rect 208092 550878 208500 550906
rect 208092 550866 208098 550878
rect 208494 550866 208500 550878
rect 208552 550866 208558 550918
rect 208034 549920 208040 549972
rect 208092 549960 208098 549972
rect 208218 549960 208224 549972
rect 208092 549932 208224 549960
rect 208092 549920 208098 549932
rect 208218 549920 208224 549932
rect 208276 549920 208282 549972
rect 208034 549444 208040 549496
rect 208092 549484 208098 549496
rect 208678 549484 208684 549496
rect 208092 549456 208684 549484
rect 208092 549444 208098 549456
rect 208678 549444 208684 549456
rect 208736 549444 208742 549496
rect 234714 548968 234720 549020
rect 234772 549008 234778 549020
rect 243546 549008 243552 549020
rect 234772 548980 243552 549008
rect 234772 548968 234778 548980
rect 243546 548968 243552 548980
rect 243604 548968 243610 549020
rect 208034 548016 208040 548068
rect 208092 548056 208098 548068
rect 208402 548056 208408 548068
rect 208092 548028 208408 548056
rect 208092 548016 208098 548028
rect 208402 548016 208408 548028
rect 208460 548056 208466 548068
rect 208770 548056 208776 548068
rect 208460 548028 208776 548056
rect 208460 548016 208466 548028
rect 208770 548016 208776 548028
rect 208828 548016 208834 548068
rect 208034 547676 208040 547728
rect 208092 547716 208098 547728
rect 208862 547716 208868 547728
rect 208092 547688 208868 547716
rect 208092 547676 208098 547688
rect 208862 547676 208868 547688
rect 208920 547676 208926 547728
rect 620010 547404 620016 547456
rect 620068 547444 620074 547456
rect 641078 547444 641084 547456
rect 620068 547416 641084 547444
rect 620068 547404 620074 547416
rect 641078 547404 641084 547416
rect 641136 547404 641142 547456
rect 208034 546588 208040 546640
rect 208092 546628 208098 546640
rect 208218 546628 208224 546640
rect 208092 546600 208224 546628
rect 208092 546588 208098 546600
rect 208218 546588 208224 546600
rect 208276 546628 208282 546640
rect 209414 546628 209420 546640
rect 208276 546600 209420 546628
rect 208276 546588 208282 546600
rect 209414 546588 209420 546600
rect 209472 546588 209478 546640
rect 208218 546384 208224 546436
rect 208276 546424 208282 546436
rect 208862 546424 208868 546436
rect 208276 546396 208868 546424
rect 208276 546384 208282 546396
rect 208862 546384 208868 546396
rect 208920 546384 208926 546436
rect 208034 546180 208040 546232
rect 208092 546220 208098 546232
rect 208770 546220 208776 546232
rect 208092 546192 208776 546220
rect 208092 546180 208098 546192
rect 208770 546180 208776 546192
rect 208828 546180 208834 546232
rect 649818 545704 649824 545756
rect 649876 545744 649882 545756
rect 651290 545744 651296 545756
rect 649876 545716 651296 545744
rect 649876 545704 649882 545716
rect 651290 545704 651296 545716
rect 651348 545704 651354 545756
rect 619090 545228 619096 545280
rect 619148 545268 619154 545280
rect 619366 545268 619372 545280
rect 619148 545240 619372 545268
rect 619148 545228 619154 545240
rect 619366 545228 619372 545240
rect 619424 545228 619430 545280
rect 208034 544072 208040 544124
rect 208092 544112 208098 544124
rect 208954 544112 208960 544124
rect 208092 544084 208960 544112
rect 208092 544072 208098 544084
rect 208954 544072 208960 544084
rect 209012 544072 209018 544124
rect 208402 543936 208408 543988
rect 208460 543976 208466 543988
rect 208586 543976 208592 543988
rect 208460 543948 208592 543976
rect 208460 543936 208466 543948
rect 208586 543936 208592 543948
rect 208644 543936 208650 543988
rect 208034 543868 208040 543920
rect 208092 543908 208098 543920
rect 208678 543908 208684 543920
rect 208092 543880 208684 543908
rect 208092 543868 208098 543880
rect 208678 543868 208684 543880
rect 208736 543868 208742 543920
rect 675854 543664 675860 543716
rect 675912 543704 675918 543716
rect 676222 543704 676228 543716
rect 675912 543676 676228 543704
rect 675912 543664 675918 543676
rect 676222 543664 676228 543676
rect 676280 543664 676286 543716
rect 675762 543596 675768 543648
rect 675820 543636 675826 543648
rect 676314 543636 676320 543648
rect 675820 543608 676320 543636
rect 675820 543596 675826 543608
rect 676314 543596 676320 543608
rect 676372 543596 676378 543648
rect 619090 543528 619096 543580
rect 619148 543568 619154 543580
rect 619274 543568 619280 543580
rect 619148 543540 619280 543568
rect 619148 543528 619154 543540
rect 619274 543528 619280 543540
rect 619332 543528 619338 543580
rect 651290 543120 651296 543172
rect 651348 543160 651354 543172
rect 661962 543160 661968 543172
rect 651348 543132 661968 543160
rect 651348 543120 651354 543132
rect 661962 543120 661968 543132
rect 662020 543120 662026 543172
rect 208034 541964 208040 542016
rect 208092 542004 208098 542016
rect 208770 542004 208776 542016
rect 208092 541976 208776 542004
rect 208092 541964 208098 541976
rect 208770 541964 208776 541976
rect 208828 541964 208834 542016
rect 641078 541896 641084 541948
rect 641136 541936 641142 541948
rect 644298 541936 644304 541948
rect 641136 541908 644304 541936
rect 641136 541896 641142 541908
rect 644298 541896 644304 541908
rect 644356 541896 644362 541948
rect 208310 541664 208316 541676
rect 208236 541636 208316 541664
rect 208236 541608 208264 541636
rect 208310 541624 208316 541636
rect 208368 541624 208374 541676
rect 208218 541556 208224 541608
rect 208276 541556 208282 541608
rect 675394 540536 675400 540588
rect 675452 540576 675458 540588
rect 676682 540576 676688 540588
rect 675452 540548 676688 540576
rect 675452 540536 675458 540548
rect 676682 540536 676688 540548
rect 676740 540536 676746 540588
rect 675578 540468 675584 540520
rect 675636 540508 675642 540520
rect 676498 540508 676504 540520
rect 675636 540480 676504 540508
rect 675636 540468 675642 540480
rect 676498 540468 676504 540480
rect 676556 540468 676562 540520
rect 675670 540400 675676 540452
rect 675728 540440 675734 540452
rect 676590 540440 676596 540452
rect 675728 540412 676596 540440
rect 675728 540400 675734 540412
rect 676590 540400 676596 540412
rect 676648 540400 676654 540452
rect 208034 540196 208040 540248
rect 208092 540236 208098 540248
rect 208678 540236 208684 540248
rect 208092 540208 208684 540236
rect 208092 540196 208098 540208
rect 208678 540196 208684 540208
rect 208736 540196 208742 540248
rect 208494 540128 208500 540180
rect 208552 540168 208558 540180
rect 214842 540168 214848 540180
rect 208552 540140 214848 540168
rect 208552 540128 208558 540140
rect 214842 540128 214848 540140
rect 214900 540128 214906 540180
rect 671898 539788 671904 539840
rect 671956 539828 671962 539840
rect 671956 539800 676360 539828
rect 671956 539788 671962 539800
rect 676332 539704 676360 539800
rect 676130 539652 676136 539704
rect 676188 539652 676194 539704
rect 676314 539652 676320 539704
rect 676372 539652 676378 539704
rect 676148 539500 676176 539652
rect 676130 539448 676136 539500
rect 676188 539448 676194 539500
rect 675486 539176 675492 539228
rect 675544 539216 675550 539228
rect 676222 539216 676228 539228
rect 675544 539188 676228 539216
rect 675544 539176 675550 539188
rect 676222 539176 676228 539188
rect 676280 539176 676286 539228
rect 644298 538700 644304 538752
rect 644356 538740 644362 538752
rect 648714 538740 648720 538752
rect 644356 538712 648720 538740
rect 644356 538700 644362 538712
rect 648714 538700 648720 538712
rect 648772 538700 648778 538752
rect 675578 537680 675584 537732
rect 675636 537720 675642 537732
rect 676314 537720 676320 537732
rect 675636 537692 676320 537720
rect 675636 537680 675642 537692
rect 676314 537680 676320 537692
rect 676372 537680 676378 537732
rect 676222 537000 676228 537052
rect 676280 537040 676286 537052
rect 676314 537040 676320 537052
rect 676280 537012 676320 537040
rect 676280 537000 676286 537012
rect 676314 537000 676320 537012
rect 676372 537000 676378 537052
rect 675670 536796 675676 536848
rect 675728 536836 675734 536848
rect 676314 536836 676320 536848
rect 675728 536808 676320 536836
rect 675728 536796 675734 536808
rect 676314 536796 676320 536808
rect 676372 536796 676378 536848
rect 675670 535980 675676 536032
rect 675728 536020 675734 536032
rect 676130 536020 676136 536032
rect 675728 535992 676136 536020
rect 675728 535980 675734 535992
rect 676130 535980 676136 535992
rect 676188 535980 676194 536032
rect 620010 535232 620016 535284
rect 620068 535272 620074 535284
rect 676130 535272 676136 535284
rect 620068 535244 676136 535272
rect 620068 535232 620074 535244
rect 676130 535232 676136 535244
rect 676188 535232 676194 535284
rect 675394 535164 675400 535216
rect 675452 535204 675458 535216
rect 675854 535204 675860 535216
rect 675452 535176 675860 535204
rect 675452 535164 675458 535176
rect 675854 535164 675860 535176
rect 675912 535164 675918 535216
rect 676038 535028 676044 535080
rect 676096 535028 676102 535080
rect 676056 534944 676084 535028
rect 676038 534892 676044 534944
rect 676096 534892 676102 534944
rect 675670 534552 675676 534604
rect 675728 534592 675734 534604
rect 676222 534592 676228 534604
rect 675728 534564 676228 534592
rect 675728 534552 675734 534564
rect 676222 534552 676228 534564
rect 676280 534552 676286 534604
rect 676038 534212 676044 534264
rect 676096 534212 676102 534264
rect 676056 534128 676084 534212
rect 676038 534076 676044 534128
rect 676096 534076 676102 534128
rect 675394 533872 675400 533924
rect 675452 533912 675458 533924
rect 675946 533912 675952 533924
rect 675452 533884 675952 533912
rect 675452 533872 675458 533884
rect 675946 533872 675952 533884
rect 676004 533912 676010 533924
rect 676314 533912 676320 533924
rect 676004 533884 676320 533912
rect 676004 533872 676010 533884
rect 676314 533872 676320 533884
rect 676372 533872 676378 533924
rect 675578 533192 675584 533244
rect 675636 533232 675642 533244
rect 676130 533232 676136 533244
rect 675636 533204 676136 533232
rect 675636 533192 675642 533204
rect 676130 533192 676136 533204
rect 676188 533192 676194 533244
rect 675486 532580 675492 532632
rect 675544 532620 675550 532632
rect 676314 532620 676320 532632
rect 675544 532592 676320 532620
rect 675544 532580 675550 532592
rect 676314 532580 676320 532592
rect 676372 532580 676378 532632
rect 620102 532512 620108 532564
rect 620160 532552 620166 532564
rect 622494 532552 622500 532564
rect 620160 532524 622500 532552
rect 620160 532512 620166 532524
rect 622494 532512 622500 532524
rect 622552 532512 622558 532564
rect 675762 532376 675768 532428
rect 675820 532416 675826 532428
rect 676130 532416 676136 532428
rect 675820 532388 676136 532416
rect 675820 532376 675826 532388
rect 676130 532376 676136 532388
rect 676188 532376 676194 532428
rect 631050 530812 631056 530864
rect 631108 530852 631114 530864
rect 676130 530852 676136 530864
rect 631108 530824 676136 530852
rect 631108 530812 631114 530824
rect 676130 530812 676136 530824
rect 676188 530812 676194 530864
rect 675670 530200 675676 530252
rect 675728 530240 675734 530252
rect 676314 530240 676320 530252
rect 675728 530212 676320 530240
rect 675728 530200 675734 530212
rect 676314 530200 676320 530212
rect 676372 530200 676378 530252
rect 635466 529724 635472 529776
rect 635524 529764 635530 529776
rect 676130 529764 676136 529776
rect 635524 529736 676136 529764
rect 635524 529724 635530 529736
rect 676130 529724 676136 529736
rect 676188 529724 676194 529776
rect 675946 529588 675952 529640
rect 676004 529628 676010 529640
rect 676130 529628 676136 529640
rect 676004 529600 676136 529628
rect 676004 529588 676010 529600
rect 676130 529588 676136 529600
rect 676188 529588 676194 529640
rect 208034 529180 208040 529232
rect 208092 529220 208098 529232
rect 208586 529220 208592 529232
rect 208092 529192 208592 529220
rect 208092 529180 208098 529192
rect 208586 529180 208592 529192
rect 208644 529180 208650 529232
rect 208126 529112 208132 529164
rect 208184 529112 208190 529164
rect 208218 529112 208224 529164
rect 208276 529112 208282 529164
rect 208144 528960 208172 529112
rect 208236 528960 208264 529112
rect 208126 528908 208132 528960
rect 208184 528908 208190 528960
rect 208218 528908 208224 528960
rect 208276 528908 208282 528960
rect 675670 527752 675676 527804
rect 675728 527792 675734 527804
rect 676222 527792 676228 527804
rect 675728 527764 676228 527792
rect 675728 527752 675734 527764
rect 676222 527752 676228 527764
rect 676280 527792 676286 527804
rect 676280 527764 676437 527792
rect 676280 527752 676286 527764
rect 208034 527004 208040 527056
rect 208092 527044 208098 527056
rect 208092 527016 208172 527044
rect 208092 527004 208098 527016
rect 208144 526908 208172 527016
rect 208218 527004 208224 527056
rect 208276 527044 208282 527056
rect 208586 527044 208592 527056
rect 208276 527016 208592 527044
rect 208276 527004 208282 527016
rect 208586 527004 208592 527016
rect 208644 527004 208650 527056
rect 208218 526908 208224 526920
rect 208144 526880 208224 526908
rect 208218 526868 208224 526880
rect 208276 526868 208282 526920
rect 208218 526024 208224 526036
rect 207962 525996 208224 526024
rect 208218 525984 208224 525996
rect 208276 525984 208282 526036
rect 659754 525100 659760 525152
rect 659812 525140 659818 525152
rect 664170 525140 664176 525152
rect 659812 525112 664176 525140
rect 659812 525100 659818 525112
rect 664170 525100 664176 525112
rect 664228 525100 664234 525152
rect 675578 524624 675584 524676
rect 675636 524664 675642 524676
rect 676314 524664 676320 524676
rect 675636 524636 676320 524664
rect 675636 524624 675642 524636
rect 676314 524624 676320 524636
rect 676372 524624 676378 524676
rect 675854 523944 675860 523996
rect 675912 523984 675918 523996
rect 676222 523984 676228 523996
rect 675912 523956 676228 523984
rect 675912 523944 675918 523956
rect 676222 523944 676228 523956
rect 676280 523944 676286 523996
rect 208017 523507 208023 523519
rect 208014 523479 208023 523507
rect 208017 523467 208023 523479
rect 208075 523508 208081 523519
rect 208303 523508 208309 523513
rect 208075 523471 208309 523508
rect 208075 523467 208081 523471
rect 208303 523461 208309 523471
rect 208361 523461 208367 523513
rect 208034 522816 208040 522868
rect 208092 522856 208098 522868
rect 208678 522856 208684 522868
rect 208092 522828 208684 522856
rect 208092 522816 208098 522828
rect 208678 522816 208684 522828
rect 208736 522816 208742 522868
rect 208037 522458 208089 522464
rect 209182 522453 209188 522463
rect 208089 522414 209188 522453
rect 209182 522411 209188 522414
rect 209240 522411 209246 522463
rect 208037 522399 208089 522406
rect 208402 522312 208408 522364
rect 208460 522352 208466 522364
rect 209506 522352 209512 522364
rect 208460 522324 209512 522352
rect 208460 522312 208466 522324
rect 209506 522312 209512 522324
rect 209564 522312 209570 522364
rect 648714 521360 648720 521412
rect 648772 521400 648778 521412
rect 658650 521400 658656 521412
rect 648772 521372 658656 521400
rect 648772 521360 648778 521372
rect 658650 521360 658656 521372
rect 658708 521360 658714 521412
rect 208218 521292 208224 521344
rect 208276 521332 208282 521344
rect 208586 521332 208592 521344
rect 208276 521304 208592 521332
rect 208276 521292 208282 521304
rect 208586 521292 208592 521304
rect 208644 521292 208650 521344
rect 208494 520816 208500 520868
rect 208552 520856 208558 520868
rect 208770 520856 208776 520868
rect 208552 520828 208776 520856
rect 208552 520816 208558 520828
rect 208770 520816 208776 520828
rect 208828 520816 208834 520868
rect 208218 520748 208224 520800
rect 208276 520788 208282 520800
rect 208586 520788 208592 520800
rect 208276 520760 208592 520788
rect 208276 520748 208282 520760
rect 208586 520748 208592 520760
rect 208644 520748 208650 520800
rect 208126 520680 208132 520732
rect 208184 520720 208190 520732
rect 208494 520720 208500 520732
rect 208184 520692 208500 520720
rect 208184 520680 208190 520692
rect 208494 520680 208500 520692
rect 208552 520680 208558 520732
rect 676314 520612 676320 520664
rect 676372 520652 676378 520664
rect 676372 520624 676452 520652
rect 676372 520612 676378 520624
rect 676424 520460 676452 520624
rect 676406 520408 676412 520460
rect 676464 520408 676470 520460
rect 675762 520272 675768 520324
rect 675820 520312 675826 520324
rect 676130 520312 676136 520324
rect 675820 520284 676136 520312
rect 675820 520272 675826 520284
rect 676130 520272 676136 520284
rect 676188 520272 676194 520324
rect 208034 519660 208040 519712
rect 208092 519700 208098 519712
rect 208586 519700 208592 519712
rect 208092 519672 208592 519700
rect 208092 519660 208098 519672
rect 208586 519660 208592 519672
rect 208644 519660 208650 519712
rect 208034 519524 208040 519576
rect 208092 519564 208098 519576
rect 208310 519564 208316 519576
rect 208092 519536 208316 519564
rect 208092 519524 208098 519536
rect 208310 519524 208316 519536
rect 208368 519564 208374 519576
rect 208770 519564 208776 519576
rect 208368 519536 208776 519564
rect 208368 519524 208374 519536
rect 208770 519524 208776 519536
rect 208828 519524 208834 519576
rect 208126 518164 208132 518216
rect 208184 518204 208190 518216
rect 208184 518176 208356 518204
rect 208184 518164 208190 518176
rect 208328 518012 208356 518176
rect 208310 517960 208316 518012
rect 208368 517960 208374 518012
rect 208218 517892 208224 517944
rect 208276 517932 208282 517944
rect 208586 517932 208592 517944
rect 208276 517904 208592 517932
rect 208276 517892 208282 517904
rect 208586 517892 208592 517904
rect 208644 517892 208650 517944
rect 668586 517008 668592 517060
rect 668644 517048 668650 517060
rect 674198 517048 674204 517060
rect 668644 517020 674204 517048
rect 668644 517008 668650 517020
rect 674198 517008 674204 517020
rect 674256 517008 674262 517060
rect 208034 516804 208040 516856
rect 208092 516844 208098 516856
rect 208770 516844 208776 516856
rect 208092 516816 208776 516844
rect 208092 516804 208098 516816
rect 208770 516804 208776 516816
rect 208828 516804 208834 516856
rect 208126 516124 208132 516176
rect 208184 516124 208190 516176
rect 208144 516040 208172 516124
rect 208126 515988 208132 516040
rect 208184 515988 208190 516040
rect 208126 514628 208132 514680
rect 208184 514668 208190 514680
rect 208494 514668 208500 514680
rect 208184 514640 208500 514668
rect 208184 514628 208190 514640
rect 208494 514628 208500 514640
rect 208552 514628 208558 514680
rect 208034 514356 208040 514408
rect 208092 514396 208098 514408
rect 208494 514396 208500 514408
rect 208092 514368 208500 514396
rect 208092 514356 208098 514368
rect 208494 514356 208500 514368
rect 208552 514356 208558 514408
rect 214842 514288 214848 514340
rect 214900 514328 214906 514340
rect 250814 514328 250820 514340
rect 214900 514300 250820 514328
rect 214900 514288 214906 514300
rect 250814 514288 250820 514300
rect 250872 514288 250878 514340
rect 244854 514222 244906 514228
rect 208030 514169 208036 514221
rect 208088 514210 208094 514221
rect 208088 514181 244854 514210
rect 208088 514169 208094 514181
rect 244854 514163 244906 514170
rect 650922 512588 650928 512640
rect 650980 512628 650986 512640
rect 659754 512628 659760 512640
rect 650980 512600 659760 512628
rect 650980 512588 650986 512600
rect 659754 512588 659760 512600
rect 659812 512588 659818 512640
rect 658650 509256 658656 509308
rect 658708 509296 658714 509308
rect 675762 509296 675768 509308
rect 658708 509268 675768 509296
rect 658708 509256 658714 509268
rect 675762 509256 675768 509268
rect 675820 509256 675826 509308
rect 619458 506196 619464 506248
rect 619516 506236 619522 506248
rect 623322 506236 623328 506248
rect 619516 506208 623328 506236
rect 619516 506196 619522 506208
rect 623322 506196 623328 506208
rect 623380 506196 623386 506248
rect 243546 505380 243552 505432
rect 243604 505420 243610 505432
rect 246858 505420 246864 505432
rect 243604 505392 246864 505420
rect 243604 505380 243610 505392
rect 246858 505380 246864 505392
rect 246916 505380 246922 505432
rect 675854 504836 675860 504888
rect 675912 504876 675918 504888
rect 676222 504876 676228 504888
rect 675912 504848 676228 504876
rect 675912 504836 675918 504848
rect 676222 504836 676228 504848
rect 676280 504836 676286 504888
rect 208494 503748 208500 503800
rect 208552 503788 208558 503800
rect 208770 503788 208776 503800
rect 208552 503760 208776 503788
rect 208552 503748 208558 503760
rect 208770 503748 208776 503760
rect 208828 503748 208834 503800
rect 675486 502660 675492 502712
rect 675544 502700 675550 502712
rect 676130 502700 676136 502712
rect 675544 502672 676136 502700
rect 675544 502660 675550 502672
rect 676130 502660 676136 502672
rect 676188 502660 676194 502712
rect 676222 502660 676228 502712
rect 676280 502700 676286 502712
rect 676682 502700 676688 502712
rect 676280 502672 676688 502700
rect 676280 502660 676286 502672
rect 676682 502660 676688 502672
rect 676740 502660 676746 502712
rect 666378 502320 666384 502372
rect 666436 502360 666442 502372
rect 668586 502360 668592 502372
rect 666436 502332 668592 502360
rect 666436 502320 666442 502332
rect 668586 502320 668592 502332
rect 668644 502320 668650 502372
rect 676130 502116 676136 502168
rect 676188 502156 676194 502168
rect 676498 502156 676504 502168
rect 676188 502128 676504 502156
rect 676188 502116 676194 502128
rect 676498 502116 676504 502128
rect 676556 502116 676562 502168
rect 675762 502048 675768 502100
rect 675820 502088 675826 502100
rect 676314 502088 676320 502100
rect 675820 502060 676320 502088
rect 675820 502048 675826 502060
rect 676314 502048 676320 502060
rect 676372 502048 676378 502100
rect 208170 501708 208176 501760
rect 208228 501748 208234 501760
rect 208514 501748 208520 501760
rect 208228 501720 208520 501748
rect 208228 501708 208234 501720
rect 208514 501708 208520 501720
rect 208572 501708 208578 501760
rect 208004 501640 208010 501692
rect 208062 501680 208068 501692
rect 208770 501680 208776 501692
rect 208062 501652 208776 501680
rect 208062 501640 208068 501652
rect 208770 501640 208776 501652
rect 208828 501640 208834 501692
rect 675762 501572 675768 501624
rect 675820 501612 675826 501624
rect 676590 501612 676596 501624
rect 675820 501584 676596 501612
rect 675820 501572 675826 501584
rect 676590 501572 676596 501584
rect 676648 501572 676654 501624
rect 675670 500416 675676 500468
rect 675728 500456 675734 500468
rect 676130 500456 676136 500468
rect 675728 500428 676136 500456
rect 675728 500416 675734 500428
rect 676130 500416 676136 500428
rect 676188 500416 676194 500468
rect 676130 499940 676136 499992
rect 676188 499980 676194 499992
rect 676406 499980 676412 499992
rect 676188 499952 676412 499980
rect 676188 499940 676194 499952
rect 676406 499940 676412 499952
rect 676464 499940 676470 499992
rect 208218 499736 208224 499788
rect 208276 499776 208282 499788
rect 208770 499776 208776 499788
rect 208276 499748 208776 499776
rect 208276 499736 208282 499748
rect 208770 499736 208776 499748
rect 208828 499736 208834 499788
rect 208126 499668 208132 499720
rect 208184 499708 208190 499720
rect 208494 499708 208500 499720
rect 208184 499680 208500 499708
rect 208184 499668 208190 499680
rect 208494 499668 208500 499680
rect 208552 499668 208558 499720
rect 662054 499124 662060 499176
rect 662112 499164 662118 499176
rect 666378 499164 666384 499176
rect 662112 499136 666384 499164
rect 662112 499124 662118 499136
rect 666378 499124 666384 499136
rect 666436 499124 666442 499176
rect 676314 498920 676320 498972
rect 676372 498920 676378 498972
rect 675578 498852 675584 498904
rect 675636 498892 675642 498904
rect 676222 498892 676228 498904
rect 675636 498864 676228 498892
rect 675636 498852 675642 498864
rect 676222 498852 676228 498864
rect 676280 498852 676286 498904
rect 676332 498836 676360 498920
rect 676314 498784 676320 498836
rect 676372 498784 676378 498836
rect 675762 498716 675768 498768
rect 675820 498756 675826 498768
rect 676222 498756 676228 498768
rect 675820 498728 676228 498756
rect 675820 498716 675826 498728
rect 676222 498716 676228 498728
rect 676280 498716 676286 498768
rect 207962 498592 208080 498620
rect 208052 498416 208080 498592
rect 208126 498512 208132 498564
rect 208184 498552 208190 498564
rect 208402 498552 208408 498564
rect 208184 498524 208408 498552
rect 208184 498512 208190 498524
rect 208402 498512 208408 498524
rect 208460 498512 208466 498564
rect 208402 498416 208408 498428
rect 208052 498388 208408 498416
rect 208402 498376 208408 498388
rect 208460 498416 208466 498428
rect 208678 498416 208684 498428
rect 208460 498388 208684 498416
rect 208460 498376 208466 498388
rect 208678 498376 208684 498388
rect 208736 498376 208742 498428
rect 676314 498376 676320 498428
rect 676372 498376 676378 498428
rect 676332 498292 676360 498376
rect 676130 498240 676136 498292
rect 676188 498280 676194 498292
rect 676314 498280 676320 498292
rect 676188 498252 676320 498280
rect 676188 498240 676194 498252
rect 676314 498240 676320 498252
rect 676372 498240 676378 498292
rect 661962 497084 661968 497136
rect 662020 497124 662026 497136
rect 669690 497124 669696 497136
rect 662020 497096 669696 497124
rect 662020 497084 662026 497096
rect 669690 497084 669696 497096
rect 669748 497084 669754 497136
rect 675762 496880 675768 496932
rect 675820 496920 675826 496932
rect 676314 496920 676320 496932
rect 675820 496892 676320 496920
rect 675820 496880 675826 496892
rect 676314 496880 676320 496892
rect 676372 496880 676378 496932
rect 208310 496268 208316 496320
rect 208368 496308 208374 496320
rect 208586 496308 208592 496320
rect 208368 496280 208592 496308
rect 208368 496268 208374 496280
rect 208586 496268 208592 496280
rect 208644 496268 208650 496320
rect 675670 496200 675676 496252
rect 675728 496240 675734 496252
rect 676130 496240 676136 496252
rect 675728 496212 676136 496240
rect 675728 496200 675734 496212
rect 676130 496200 676136 496212
rect 676188 496240 676194 496252
rect 676314 496240 676320 496252
rect 676188 496212 676320 496240
rect 676188 496200 676194 496212
rect 676314 496200 676320 496212
rect 676372 496200 676378 496252
rect 208034 495928 208040 495980
rect 208092 495968 208098 495980
rect 208494 495968 208500 495980
rect 208092 495940 208500 495968
rect 208092 495928 208098 495940
rect 208494 495928 208500 495940
rect 208552 495928 208558 495980
rect 675394 495452 675400 495504
rect 675452 495492 675458 495504
rect 675854 495492 675860 495504
rect 675452 495464 675860 495492
rect 675452 495452 675458 495464
rect 675854 495452 675860 495464
rect 675912 495452 675918 495504
rect 675854 495316 675860 495368
rect 675912 495356 675918 495368
rect 676038 495356 676044 495368
rect 675912 495328 676044 495356
rect 675912 495316 675918 495328
rect 676038 495316 676044 495328
rect 676096 495316 676102 495368
rect 673370 495112 673376 495164
rect 673428 495152 673434 495164
rect 676130 495152 676136 495164
rect 673428 495124 676136 495152
rect 673428 495112 673434 495124
rect 676130 495112 676136 495124
rect 676188 495112 676194 495164
rect 645402 494432 645408 494484
rect 645460 494472 645466 494484
rect 673370 494472 673376 494484
rect 645460 494444 673376 494472
rect 645460 494432 645466 494444
rect 673370 494432 673376 494444
rect 673428 494432 673434 494484
rect 675302 494160 675308 494212
rect 675360 494200 675366 494212
rect 675670 494200 675676 494212
rect 675360 494172 675676 494200
rect 675360 494160 675366 494172
rect 675670 494160 675676 494172
rect 675728 494200 675734 494212
rect 676222 494200 676228 494212
rect 675728 494172 676228 494200
rect 675728 494160 675734 494172
rect 676222 494160 676228 494172
rect 676280 494160 676286 494212
rect 675670 493752 675676 493804
rect 675728 493792 675734 493804
rect 676314 493792 676320 493804
rect 675728 493764 676320 493792
rect 675728 493752 675734 493764
rect 676314 493752 676320 493764
rect 676372 493752 676378 493804
rect 669690 493276 669696 493328
rect 669748 493316 669754 493328
rect 675670 493316 675676 493328
rect 669748 493288 675676 493316
rect 669748 493276 669754 493288
rect 675670 493276 675676 493288
rect 675728 493276 675734 493328
rect 208126 493208 208132 493260
rect 208184 493248 208190 493260
rect 208678 493248 208684 493260
rect 208184 493220 208684 493248
rect 208184 493208 208190 493220
rect 208678 493208 208684 493220
rect 208736 493208 208742 493260
rect 675394 493072 675400 493124
rect 675452 493112 675458 493124
rect 676314 493112 676320 493124
rect 675452 493084 676320 493112
rect 675452 493072 675458 493084
rect 676314 493072 676320 493084
rect 676372 493072 676378 493124
rect 208034 492596 208040 492648
rect 208092 492636 208098 492648
rect 208678 492636 208684 492648
rect 208092 492608 208684 492636
rect 208092 492596 208098 492608
rect 208678 492596 208684 492608
rect 208736 492596 208742 492648
rect 660858 492188 660864 492240
rect 660916 492228 660922 492240
rect 675762 492228 675768 492240
rect 660916 492200 675768 492228
rect 660916 492188 660922 492200
rect 675762 492188 675768 492200
rect 675820 492228 675826 492240
rect 676130 492228 676136 492240
rect 675820 492200 676136 492228
rect 675820 492188 675826 492200
rect 676130 492188 676136 492200
rect 676188 492188 676194 492240
rect 675578 491780 675584 491832
rect 675636 491820 675642 491832
rect 676314 491820 676320 491832
rect 675636 491792 676320 491820
rect 675636 491780 675642 491792
rect 676314 491780 676320 491792
rect 676372 491780 676378 491832
rect 645402 491576 645408 491628
rect 645460 491616 645466 491628
rect 650922 491616 650928 491628
rect 645460 491588 650928 491616
rect 645460 491576 645466 491588
rect 650922 491576 650928 491588
rect 650980 491576 650986 491628
rect 675486 491576 675492 491628
rect 675544 491616 675550 491628
rect 676130 491616 676136 491628
rect 675544 491588 676136 491616
rect 675544 491576 675550 491588
rect 676130 491576 676136 491588
rect 676188 491576 676194 491628
rect 208034 490556 208040 490608
rect 208092 490556 208098 490608
rect 208052 489452 208080 490556
rect 675854 490420 675860 490472
rect 675912 490460 675918 490472
rect 676314 490460 676320 490472
rect 675912 490432 676320 490460
rect 675912 490420 675918 490432
rect 676314 490420 676320 490432
rect 676372 490420 676378 490472
rect 208126 490352 208132 490404
rect 208184 490392 208190 490404
rect 208494 490392 208500 490404
rect 208184 490364 208500 490392
rect 208184 490352 208190 490364
rect 208494 490352 208500 490364
rect 208552 490352 208558 490404
rect 208218 490284 208224 490336
rect 208276 490324 208282 490336
rect 208770 490324 208776 490336
rect 208276 490296 208776 490324
rect 208276 490284 208282 490296
rect 208770 490284 208776 490296
rect 208828 490284 208834 490336
rect 208034 489400 208040 489452
rect 208092 489400 208098 489452
rect 675762 489400 675768 489452
rect 675820 489440 675826 489452
rect 676314 489440 676320 489452
rect 675820 489412 676320 489440
rect 675820 489400 675826 489412
rect 676314 489400 676320 489412
rect 676372 489400 676378 489452
rect 208034 488652 208040 488704
rect 208092 488692 208098 488704
rect 208678 488692 208684 488704
rect 208092 488664 208684 488692
rect 208092 488652 208098 488664
rect 208678 488652 208684 488664
rect 208736 488652 208742 488704
rect 208034 487156 208040 487208
rect 208092 487196 208098 487208
rect 208954 487196 208960 487208
rect 208092 487168 208960 487196
rect 208092 487156 208098 487168
rect 208954 487156 208960 487168
rect 209012 487156 209018 487208
rect 675854 486952 675860 487004
rect 675912 486992 675918 487004
rect 676038 486992 676044 487004
rect 675912 486964 676044 486992
rect 675912 486952 675918 486964
rect 676038 486952 676044 486964
rect 676096 486992 676102 487004
rect 676096 486964 676437 486992
rect 676096 486952 676102 486964
rect 675670 486068 675676 486120
rect 675728 486108 675734 486120
rect 676314 486108 676320 486120
rect 675728 486080 676320 486108
rect 675728 486068 675734 486080
rect 676314 486068 676320 486080
rect 676372 486068 676378 486120
rect 208678 485796 208684 485848
rect 208736 485796 208742 485848
rect 208402 485728 208408 485780
rect 208460 485768 208466 485780
rect 208696 485768 208724 485796
rect 208460 485740 208724 485768
rect 208460 485728 208466 485740
rect 675854 483960 675860 484012
rect 675912 484000 675918 484012
rect 676314 484000 676320 484012
rect 675912 483972 676320 484000
rect 675912 483960 675918 483972
rect 676314 483960 676320 483972
rect 676372 483960 676378 484012
rect 675486 483552 675492 483604
rect 675544 483592 675550 483604
rect 676222 483592 676228 483604
rect 675544 483564 676228 483592
rect 675544 483552 675550 483564
rect 676222 483552 676228 483564
rect 676280 483552 676286 483604
rect 675762 483416 675768 483468
rect 675820 483456 675826 483468
rect 676222 483456 676228 483468
rect 675820 483428 676228 483456
rect 675820 483416 675826 483428
rect 676222 483416 676228 483428
rect 676280 483416 676286 483468
rect 659754 483348 659760 483400
rect 659812 483388 659818 483400
rect 675854 483388 675860 483400
rect 659812 483360 675860 483388
rect 659812 483348 659818 483360
rect 675854 483348 675860 483360
rect 675912 483348 675918 483400
rect 641078 483212 641084 483264
rect 641136 483252 641142 483264
rect 645402 483252 645408 483264
rect 641136 483224 645408 483252
rect 641136 483212 641142 483224
rect 645402 483212 645408 483224
rect 645460 483212 645466 483264
rect 208218 481716 208224 481768
rect 208276 481716 208282 481768
rect 208236 481496 208264 481716
rect 676038 481648 676044 481700
rect 676096 481688 676102 481700
rect 676570 481688 676576 481700
rect 676096 481660 676576 481688
rect 676096 481648 676102 481660
rect 676570 481648 676576 481660
rect 676628 481648 676634 481700
rect 675486 481512 675492 481564
rect 675544 481552 675550 481564
rect 676038 481552 676044 481564
rect 675544 481524 676044 481552
rect 675544 481512 675550 481524
rect 676038 481512 676044 481524
rect 676096 481512 676102 481564
rect 208218 481444 208224 481496
rect 208276 481444 208282 481496
rect 221466 478928 221472 478980
rect 221524 478968 221530 478980
rect 250814 478968 250820 478980
rect 221524 478940 250820 478968
rect 221524 478928 221530 478940
rect 250814 478928 250820 478940
rect 250872 478928 250878 478980
rect 657546 475528 657552 475580
rect 657604 475568 657610 475580
rect 661962 475568 661968 475580
rect 657604 475540 661968 475568
rect 657604 475528 657610 475540
rect 661962 475528 661968 475540
rect 662020 475528 662026 475580
rect 671898 475392 671904 475444
rect 671956 475432 671962 475444
rect 676222 475432 676228 475444
rect 671956 475404 676228 475432
rect 671956 475392 671962 475404
rect 676222 475392 676228 475404
rect 676280 475392 676286 475444
rect 211162 475052 211168 475104
rect 211220 475092 211226 475104
rect 219258 475092 219264 475104
rect 211220 475064 219264 475092
rect 211220 475052 211226 475064
rect 219258 475052 219264 475064
rect 219316 475052 219322 475104
rect 207942 474616 207948 474668
rect 208000 474656 208006 474668
rect 208402 474656 208408 474668
rect 208000 474628 208408 474656
rect 208000 474616 208006 474628
rect 208402 474616 208408 474628
rect 208460 474616 208466 474668
rect 208034 474236 208040 474288
rect 208092 474276 208098 474288
rect 208862 474276 208868 474288
rect 208092 474248 208868 474276
rect 208092 474236 208098 474248
rect 208862 474236 208868 474248
rect 208920 474236 208926 474288
rect 638870 473828 638876 473880
rect 638928 473868 638934 473880
rect 641078 473868 641084 473880
rect 638928 473840 641084 473868
rect 638928 473828 638934 473840
rect 641078 473828 641084 473840
rect 641136 473828 641142 473880
rect 208034 471026 208040 471038
rect 207962 470998 208040 471026
rect 208034 470986 208040 470998
rect 208092 471012 208098 471038
rect 209046 471012 209052 471024
rect 208092 470986 209052 471012
rect 208052 470984 209052 470986
rect 209046 470972 209052 470984
rect 209104 470972 209110 471024
rect 208218 470904 208224 470956
rect 208276 470944 208282 470956
rect 208770 470944 208776 470956
rect 208276 470916 208776 470944
rect 208276 470904 208282 470916
rect 208770 470904 208776 470916
rect 208828 470904 208834 470956
rect 208310 470836 208316 470888
rect 208368 470836 208374 470888
rect 208218 470632 208224 470684
rect 208276 470672 208282 470684
rect 208328 470672 208356 470836
rect 208276 470644 208356 470672
rect 208276 470632 208282 470644
rect 208126 470360 208132 470412
rect 208184 470400 208190 470412
rect 208494 470400 208500 470412
rect 208184 470372 208500 470400
rect 208184 470360 208190 470372
rect 208494 470360 208500 470372
rect 208552 470360 208558 470412
rect 208034 467640 208040 467692
rect 208092 467680 208098 467692
rect 208862 467680 208868 467692
rect 208092 467652 208868 467680
rect 208092 467640 208098 467652
rect 208862 467640 208868 467652
rect 208920 467640 208926 467692
rect 208402 466348 208408 466400
rect 208460 466388 208466 466400
rect 208460 466360 208632 466388
rect 208460 466348 208466 466360
rect 208034 466280 208040 466332
rect 208092 466320 208098 466332
rect 208092 466292 208540 466320
rect 208092 466280 208098 466292
rect 208512 466196 208540 466292
rect 208494 466144 208500 466196
rect 208552 466144 208558 466196
rect 208604 466128 208632 466360
rect 208034 466076 208040 466128
rect 208092 466116 208098 466128
rect 208586 466116 208592 466128
rect 208092 466088 208592 466116
rect 208092 466076 208098 466088
rect 208586 466076 208592 466088
rect 208644 466076 208650 466128
rect 208034 465464 208040 465516
rect 208092 465504 208098 465516
rect 208770 465504 208776 465516
rect 208092 465476 208776 465504
rect 208092 465464 208098 465476
rect 208770 465464 208776 465476
rect 208828 465464 208834 465516
rect 208034 464784 208040 464836
rect 208092 464824 208098 464836
rect 209046 464824 209052 464836
rect 208092 464796 209052 464824
rect 208092 464784 208098 464796
rect 209046 464784 209052 464796
rect 209104 464784 209110 464836
rect 620194 464036 620200 464088
rect 620252 464076 620258 464088
rect 621298 464076 621304 464088
rect 620252 464048 621304 464076
rect 620252 464036 620258 464048
rect 621298 464036 621304 464048
rect 621356 464036 621362 464088
rect 656442 462880 656448 462932
rect 656500 462920 656506 462932
rect 671898 462920 671904 462932
rect 656500 462892 671904 462920
rect 656500 462880 656506 462892
rect 671898 462880 671904 462892
rect 671956 462880 671962 462932
rect 208034 462812 208040 462864
rect 208092 462852 208098 462864
rect 208862 462852 208868 462864
rect 208092 462824 208868 462852
rect 208092 462812 208098 462824
rect 208862 462812 208868 462824
rect 208920 462812 208926 462864
rect 208218 461792 208224 461844
rect 208276 461832 208282 461844
rect 208586 461832 208592 461844
rect 208276 461804 208592 461832
rect 208276 461792 208282 461804
rect 208586 461792 208592 461804
rect 208644 461792 208650 461844
rect 208126 459140 208132 459192
rect 208184 459140 208190 459192
rect 208494 459180 208500 459192
rect 208328 459152 208500 459180
rect 208144 459044 208172 459140
rect 208328 459124 208356 459152
rect 208494 459140 208500 459152
rect 208552 459140 208558 459192
rect 208310 459072 208316 459124
rect 208368 459072 208374 459124
rect 208494 459044 208500 459056
rect 208144 459016 208500 459044
rect 208494 459004 208500 459016
rect 208552 459044 208558 459056
rect 208770 459044 208776 459056
rect 208552 459016 208776 459044
rect 208552 459004 208558 459016
rect 208770 459004 208776 459016
rect 208828 459004 208834 459056
rect 644482 458460 644488 458512
rect 644540 458500 644546 458512
rect 656442 458500 656448 458512
rect 644540 458472 656448 458500
rect 644540 458460 644546 458472
rect 656442 458460 656448 458472
rect 656500 458460 656506 458512
rect 208034 457440 208040 457492
rect 208092 457480 208098 457492
rect 208402 457480 208408 457492
rect 208092 457452 208408 457480
rect 208092 457440 208098 457452
rect 208402 457440 208408 457452
rect 208460 457440 208466 457492
rect 623322 454652 623328 454704
rect 623380 454692 623386 454704
rect 644482 454692 644488 454704
rect 623380 454664 644488 454692
rect 623380 454652 623386 454664
rect 644482 454652 644488 454664
rect 644540 454652 644546 454704
rect 208126 447512 208132 447564
rect 208184 447552 208190 447564
rect 208862 447552 208868 447564
rect 208184 447524 208868 447552
rect 208184 447512 208190 447524
rect 208862 447512 208868 447524
rect 208920 447512 208926 447564
rect 207942 447202 207948 447254
rect 208000 447242 208006 447254
rect 208402 447242 208408 447254
rect 208000 447214 208408 447242
rect 208000 447202 208006 447214
rect 208402 447202 208408 447214
rect 208460 447202 208466 447254
rect 208218 447104 208224 447156
rect 208276 447104 208282 447156
rect 208236 446884 208264 447104
rect 208218 446832 208224 446884
rect 208276 446832 208282 446884
rect 208034 446628 208040 446680
rect 208092 446668 208098 446680
rect 208678 446668 208684 446680
rect 208092 446640 208684 446668
rect 208092 446628 208098 446640
rect 208678 446628 208684 446640
rect 208736 446628 208742 446680
rect 627830 446288 627836 446340
rect 627888 446328 627894 446340
rect 638870 446328 638876 446340
rect 627888 446300 638876 446328
rect 627888 446288 627894 446300
rect 638870 446288 638876 446300
rect 638928 446288 638934 446340
rect 208034 444384 208040 444436
rect 208092 444424 208098 444436
rect 208770 444424 208776 444436
rect 208092 444396 208776 444424
rect 208092 444384 208098 444396
rect 208770 444384 208776 444396
rect 208828 444384 208834 444436
rect 645402 444112 645408 444164
rect 645460 444152 645466 444164
rect 657546 444152 657552 444164
rect 645460 444124 657552 444152
rect 645460 444112 645466 444124
rect 657546 444112 657552 444124
rect 657604 444112 657610 444164
rect 207962 443608 208080 443626
rect 208770 443608 208776 443620
rect 207962 443598 208776 443608
rect 208052 443580 208776 443598
rect 208770 443568 208776 443580
rect 208828 443568 208834 443620
rect 208126 441596 208132 441648
rect 208184 441636 208190 441648
rect 208494 441636 208500 441648
rect 208184 441608 208500 441636
rect 208184 441596 208190 441608
rect 208494 441596 208500 441608
rect 208552 441596 208558 441648
rect 208218 441528 208224 441580
rect 208276 441568 208282 441580
rect 208276 441540 208540 441568
rect 208276 441528 208282 441540
rect 208512 441444 208540 441540
rect 208586 441528 208592 441580
rect 208644 441528 208650 441580
rect 208604 441444 208632 441528
rect 208494 441392 208500 441444
rect 208552 441392 208558 441444
rect 208586 441392 208592 441444
rect 208644 441392 208650 441444
rect 208034 438196 208040 438248
rect 208092 438236 208098 438248
rect 208494 438236 208500 438248
rect 208092 438208 208500 438236
rect 208092 438196 208098 438208
rect 208494 438196 208500 438208
rect 208552 438236 208558 438248
rect 208862 438236 208868 438248
rect 208552 438208 208868 438236
rect 208552 438196 208558 438208
rect 208862 438196 208868 438208
rect 208920 438196 208926 438248
rect 208034 437380 208040 437432
rect 208092 437420 208098 437432
rect 208678 437420 208684 437432
rect 208092 437392 208684 437420
rect 208092 437380 208098 437392
rect 208678 437380 208684 437392
rect 208736 437420 208742 437432
rect 208954 437420 208960 437432
rect 208736 437392 208960 437420
rect 208736 437380 208742 437392
rect 208954 437380 208960 437392
rect 209012 437380 209018 437432
rect 208126 437312 208132 437364
rect 208184 437352 208190 437364
rect 208402 437352 208408 437364
rect 208184 437324 208408 437352
rect 208184 437312 208190 437324
rect 208402 437312 208408 437324
rect 208460 437312 208466 437364
rect 625622 437108 625628 437160
rect 625680 437148 625686 437160
rect 627830 437148 627836 437160
rect 625680 437120 627836 437148
rect 625680 437108 625686 437120
rect 627830 437108 627836 437120
rect 627888 437108 627894 437160
rect 641078 436836 641084 436888
rect 641136 436876 641142 436888
rect 645402 436876 645408 436888
rect 641136 436848 645408 436876
rect 641136 436836 641142 436848
rect 645402 436836 645408 436848
rect 645460 436836 645466 436888
rect 208034 433640 208040 433692
rect 208092 433680 208098 433692
rect 208770 433680 208776 433692
rect 208092 433652 208776 433680
rect 208092 433640 208098 433652
rect 208770 433640 208776 433652
rect 208828 433680 208834 433692
rect 209506 433680 209512 433692
rect 208828 433652 209512 433680
rect 208828 433640 208834 433652
rect 209506 433640 209512 433652
rect 209564 433640 209570 433692
rect 208954 432008 208960 432060
rect 209012 432048 209018 432060
rect 210150 432048 210156 432060
rect 209012 432020 210156 432048
rect 209012 432008 209018 432020
rect 210150 432008 210156 432020
rect 210208 432008 210214 432060
rect 208126 431736 208132 431788
rect 208184 431736 208190 431788
rect 208144 431516 208172 431736
rect 208126 431464 208132 431516
rect 208184 431464 208190 431516
rect 208126 427384 208132 427436
rect 208184 427424 208190 427436
rect 209966 427424 209972 427436
rect 208184 427396 209972 427424
rect 208184 427384 208190 427396
rect 209966 427384 209972 427396
rect 210024 427384 210030 427436
rect 635466 426636 635472 426688
rect 635524 426676 635530 426688
rect 641078 426676 641084 426688
rect 635524 426648 641084 426676
rect 635524 426636 635530 426648
rect 641078 426636 641084 426648
rect 641136 426636 641142 426688
rect 620102 425276 620108 425328
rect 620160 425316 620166 425328
rect 625622 425316 625628 425328
rect 620160 425288 625628 425316
rect 620160 425276 620166 425288
rect 625622 425276 625628 425288
rect 625680 425276 625686 425328
rect 620194 425004 620200 425056
rect 620252 425044 620258 425056
rect 621114 425044 621120 425056
rect 620252 425016 621120 425044
rect 620252 425004 620258 425016
rect 621114 425004 621120 425016
rect 621172 425004 621178 425056
rect 620286 423168 620292 423220
rect 620344 423208 620350 423220
rect 635466 423208 635472 423220
rect 620344 423180 635472 423208
rect 620344 423168 620350 423180
rect 635466 423168 635472 423180
rect 635524 423168 635530 423220
rect 208310 422080 208316 422132
rect 208368 422120 208374 422132
rect 226986 422120 226992 422132
rect 208368 422092 226992 422120
rect 208368 422080 208374 422092
rect 226986 422080 226992 422092
rect 227044 422080 227050 422132
rect 208034 422012 208040 422064
rect 208092 422052 208098 422064
rect 228090 422052 228096 422064
rect 208092 422024 228096 422052
rect 208092 422012 208098 422024
rect 228090 422012 228096 422024
rect 228148 422012 228154 422064
rect 232230 421536 232236 421588
rect 232288 421576 232294 421588
rect 250814 421576 250820 421588
rect 232288 421548 250820 421576
rect 232288 421536 232294 421548
rect 250814 421536 250820 421548
rect 250872 421536 250878 421588
rect 618998 414600 619004 414652
rect 619056 414640 619062 414652
rect 619182 414640 619188 414652
rect 619056 414612 619188 414640
rect 619056 414600 619062 414612
rect 619182 414600 619188 414612
rect 619240 414600 619246 414652
rect 208126 411200 208132 411252
rect 208184 411240 208190 411252
rect 209966 411240 209972 411252
rect 208184 411212 209972 411240
rect 208184 411200 208190 411212
rect 209966 411200 209972 411212
rect 210024 411200 210030 411252
rect 208034 410520 208040 410572
rect 208092 410560 208098 410572
rect 209506 410560 209512 410572
rect 208092 410532 209512 410560
rect 208092 410520 208098 410532
rect 209506 410520 209512 410532
rect 209564 410560 209570 410572
rect 210058 410560 210064 410572
rect 209564 410532 210064 410560
rect 209564 410520 209570 410532
rect 210058 410520 210064 410532
rect 210116 410520 210122 410572
rect 208034 409710 208040 409722
rect 207968 409682 208040 409710
rect 208034 409670 208040 409682
rect 208092 409670 208098 409722
rect 208034 408276 208040 408328
rect 208092 408316 208098 408328
rect 208310 408316 208316 408328
rect 208092 408288 208316 408316
rect 208092 408276 208098 408288
rect 208310 408276 208316 408288
rect 208368 408276 208374 408328
rect 208034 407528 208040 407580
rect 208092 407568 208098 407580
rect 210242 407568 210248 407580
rect 208092 407540 210248 407568
rect 208092 407528 208098 407540
rect 210242 407528 210248 407540
rect 210300 407528 210306 407580
rect 208126 407188 208132 407240
rect 208184 407228 208190 407240
rect 210150 407228 210156 407240
rect 208184 407200 210156 407228
rect 208184 407188 208190 407200
rect 210150 407188 210156 407200
rect 210208 407188 210214 407240
rect 208034 405488 208040 405540
rect 208092 405528 208098 405540
rect 208862 405528 208868 405540
rect 208092 405500 208868 405528
rect 208092 405488 208098 405500
rect 208862 405488 208868 405500
rect 208920 405488 208926 405540
rect 248146 396580 248152 396632
rect 248204 396620 248210 396632
rect 252194 396620 252200 396632
rect 248204 396592 252200 396620
rect 248204 396580 248210 396592
rect 252194 396580 252200 396592
rect 252252 396580 252258 396632
rect 208126 390664 208132 390716
rect 208184 390704 208190 390716
rect 210242 390704 210248 390716
rect 208184 390676 210248 390704
rect 208184 390664 208190 390676
rect 210242 390664 210248 390676
rect 210300 390664 210306 390716
rect 208310 390392 208316 390444
rect 208368 390432 208374 390444
rect 210058 390432 210064 390444
rect 208368 390404 210064 390432
rect 208368 390392 208374 390404
rect 210058 390392 210064 390404
rect 210116 390392 210122 390444
rect 208034 389820 208040 389832
rect 207962 389792 208040 389820
rect 208034 389780 208040 389792
rect 208092 389820 208098 389832
rect 208862 389820 208868 389832
rect 208092 389792 208868 389820
rect 208092 389780 208098 389792
rect 208862 389780 208868 389792
rect 208920 389780 208926 389832
rect 208005 387271 208011 387323
rect 208063 387318 208069 387323
rect 208215 387318 208221 387327
rect 208063 387282 208221 387318
rect 208063 387271 208069 387282
rect 208215 387275 208221 387282
rect 208273 387275 208279 387327
rect 208034 386312 208040 386364
rect 208092 386352 208098 386364
rect 208402 386352 208408 386364
rect 208092 386324 208408 386352
rect 208092 386312 208098 386324
rect 208402 386312 208408 386324
rect 208460 386312 208466 386364
rect 228090 386244 228096 386296
rect 228148 386284 228154 386296
rect 250078 386284 250084 386296
rect 228148 386256 250084 386284
rect 228148 386244 228154 386256
rect 250078 386244 250084 386256
rect 250136 386244 250142 386296
rect 227630 385428 227636 385480
rect 227688 385468 227694 385480
rect 228090 385468 228096 385480
rect 227688 385440 228096 385468
rect 227688 385428 227694 385440
rect 228090 385428 228096 385440
rect 228148 385428 228154 385480
rect 208126 385088 208132 385140
rect 208184 385128 208190 385140
rect 208586 385128 208592 385140
rect 208184 385100 208592 385128
rect 208184 385088 208190 385100
rect 208586 385088 208592 385100
rect 208644 385088 208650 385140
rect 208034 383456 208040 383508
rect 208092 383496 208098 383508
rect 208402 383496 208408 383508
rect 208092 383468 208408 383496
rect 208092 383456 208098 383468
rect 208402 383456 208408 383468
rect 208460 383456 208466 383508
rect 208034 383048 208040 383100
rect 208092 383088 208098 383100
rect 208586 383088 208592 383100
rect 208092 383060 208592 383088
rect 208092 383048 208098 383060
rect 208586 383048 208592 383060
rect 208644 383048 208650 383100
rect 208402 380600 208408 380652
rect 208460 380640 208466 380652
rect 210426 380640 210432 380652
rect 208460 380612 210432 380640
rect 208460 380600 208466 380612
rect 210426 380600 210432 380612
rect 210484 380600 210490 380652
rect 208026 379854 208032 379906
rect 208084 379902 208090 379906
rect 208230 379902 208236 379908
rect 208084 379862 208236 379902
rect 208084 379854 208090 379862
rect 208230 379856 208236 379862
rect 208288 379896 208294 379908
rect 208288 379868 208298 379896
rect 208288 379856 208294 379868
rect 209414 372032 209420 372084
rect 209472 372072 209478 372084
rect 210518 372072 210524 372084
rect 209472 372044 210524 372072
rect 209472 372032 209478 372044
rect 210518 372032 210524 372044
rect 210576 372032 210582 372084
rect 210518 367680 210524 367732
rect 210576 367720 210582 367732
rect 217050 367720 217056 367732
rect 210576 367692 217056 367720
rect 210576 367680 210582 367692
rect 217050 367680 217056 367692
rect 217108 367680 217114 367732
rect 217050 357616 217056 357668
rect 217108 357656 217114 357668
rect 221466 357656 221472 357668
rect 217108 357628 221472 357656
rect 217108 357616 217114 357628
rect 221466 357616 221472 357628
rect 221524 357616 221530 357668
rect 221466 329260 221472 329312
rect 221524 329300 221530 329312
rect 222386 329300 222392 329312
rect 221524 329272 222392 329300
rect 221524 329260 221530 329272
rect 222386 329260 222392 329272
rect 222444 329260 222450 329312
rect 222386 320488 222392 320540
rect 222444 320528 222450 320540
rect 233702 320528 233708 320540
rect 222444 320500 233708 320528
rect 222444 320488 222450 320500
rect 233702 320488 233708 320500
rect 233760 320488 233766 320540
rect 209322 316068 209328 316120
rect 209380 316108 209386 316120
rect 217050 316108 217056 316120
rect 209380 316080 217056 316108
rect 209380 316068 209386 316080
rect 217050 316068 217056 316080
rect 217108 316068 217114 316120
rect 217050 302808 217056 302860
rect 217108 302848 217114 302860
rect 229194 302848 229200 302860
rect 217108 302820 229200 302848
rect 217108 302808 217114 302820
rect 229194 302808 229200 302820
rect 229252 302808 229258 302860
rect 233702 297436 233708 297488
rect 233760 297476 233766 297488
rect 238026 297476 238032 297488
rect 233760 297448 238032 297476
rect 233760 297436 233766 297448
rect 238026 297436 238032 297448
rect 238084 297436 238090 297488
rect 229194 293968 229200 294020
rect 229252 294008 229258 294020
rect 233702 294008 233708 294020
rect 229252 293980 233708 294008
rect 229252 293968 229258 293980
rect 233702 293968 233708 293980
rect 233760 293968 233766 294020
rect 238026 290976 238032 291028
rect 238084 291016 238090 291028
rect 240234 291016 240240 291028
rect 238084 290988 240240 291016
rect 238084 290976 238090 290988
rect 240234 290976 240240 290988
rect 240292 290976 240298 291028
rect 233702 287508 233708 287560
rect 233760 287548 233766 287560
rect 244650 287548 244656 287560
rect 233760 287520 244656 287548
rect 233760 287508 233766 287520
rect 244650 287508 244656 287520
rect 244708 287508 244714 287560
rect 621114 285400 621120 285452
rect 621172 285440 621178 285452
rect 623046 285440 623052 285452
rect 621172 285412 623052 285440
rect 621172 285400 621178 285412
rect 623046 285400 623052 285412
rect 623104 285400 623110 285452
rect 229746 284516 229752 284568
rect 229804 284556 229810 284568
rect 232322 284556 232328 284568
rect 229804 284528 232328 284556
rect 229804 284516 229810 284528
rect 232322 284516 232328 284528
rect 232380 284516 232386 284568
rect 232322 284040 232328 284092
rect 232380 284080 232386 284092
rect 250170 284080 250176 284092
rect 232380 284052 250176 284080
rect 232380 284040 232386 284052
rect 250170 284040 250176 284052
rect 250228 284040 250234 284092
rect 634912 281126 636294 281152
rect 634912 281046 634944 281126
rect 634910 280950 634944 281046
rect 634912 280890 634944 280950
rect 636264 281046 636294 281126
rect 636264 280950 638626 281046
rect 636264 280890 636294 280950
rect 634912 280868 636294 280890
rect 638530 280892 638626 280950
rect 642298 280916 643130 280936
rect 638530 280796 639454 280892
rect 642298 280880 642326 280916
rect 640222 280784 642326 280880
rect 639514 280748 639520 280760
rect 639475 280720 639520 280748
rect 639514 280708 639520 280720
rect 639572 280708 639578 280760
rect 248422 280504 248428 280556
rect 248480 280544 248486 280556
rect 257438 280544 257444 280556
rect 248480 280516 257444 280544
rect 248480 280504 248486 280516
rect 257438 280504 257444 280516
rect 257496 280504 257502 280556
rect 617158 280504 617164 280556
rect 617216 280544 617222 280556
rect 625070 280544 625076 280556
rect 617216 280516 625076 280544
rect 617216 280504 617222 280516
rect 625070 280504 625076 280516
rect 625128 280504 625134 280556
rect 250630 280436 250636 280488
rect 250688 280476 250694 280488
rect 262222 280476 262228 280488
rect 250688 280448 262228 280476
rect 250688 280436 250694 280448
rect 262222 280436 262228 280448
rect 262280 280436 262286 280488
rect 607590 280436 607596 280488
rect 607648 280476 607654 280488
rect 619826 280476 619832 280488
rect 607648 280448 619832 280476
rect 607648 280436 607654 280448
rect 619826 280436 619832 280448
rect 619884 280436 619890 280488
rect 251182 280368 251188 280420
rect 251240 280408 251246 280420
rect 362870 280408 362876 280420
rect 251240 280380 362876 280408
rect 251240 280368 251246 280380
rect 362870 280368 362876 280380
rect 362928 280368 362934 280420
rect 588270 280368 588276 280420
rect 588328 280408 588334 280420
rect 622034 280408 622040 280420
rect 588328 280380 622040 280408
rect 588328 280368 588334 280380
rect 622034 280368 622040 280380
rect 622092 280368 622098 280420
rect 250538 280300 250544 280352
rect 250596 280340 250602 280352
rect 420278 280340 420284 280352
rect 250596 280312 420284 280340
rect 250596 280300 250602 280312
rect 420278 280300 420284 280312
rect 420336 280300 420342 280352
rect 434998 280300 435004 280352
rect 435056 280340 435062 280352
rect 621114 280340 621120 280352
rect 435056 280312 621120 280340
rect 435056 280300 435062 280312
rect 621114 280300 621120 280312
rect 621172 280300 621178 280352
rect 640222 280348 640318 280784
rect 642298 280712 642326 280784
rect 643110 280880 643130 280916
rect 643110 280784 643140 280880
rect 643110 280712 643130 280784
rect 642298 280692 643130 280712
rect 251366 280232 251372 280284
rect 251424 280272 251430 280284
rect 271882 280272 271888 280284
rect 251424 280244 271888 280272
rect 251424 280232 251430 280244
rect 271882 280232 271888 280244
rect 271940 280232 271946 280284
rect 360570 280232 360576 280284
rect 360628 280272 360634 280284
rect 549906 280272 549912 280284
rect 360628 280244 549912 280272
rect 360628 280232 360634 280244
rect 549906 280232 549912 280244
rect 549964 280232 549970 280284
rect 573918 280232 573924 280284
rect 573976 280272 573982 280284
rect 621942 280272 621948 280284
rect 573976 280244 621948 280272
rect 573976 280232 573982 280244
rect 621942 280232 621948 280244
rect 622000 280232 622006 280284
rect 639358 280254 640318 280348
rect 639358 280252 640298 280254
rect 252102 280164 252108 280216
rect 252160 280204 252166 280216
rect 675946 280204 675952 280216
rect 252160 280176 675952 280204
rect 252160 280164 252166 280176
rect 675946 280164 675952 280176
rect 676004 280164 676010 280216
rect 252378 280096 252384 280148
rect 252436 280136 252442 280148
rect 643194 280136 643200 280148
rect 252436 280108 643200 280136
rect 252436 280096 252442 280108
rect 643194 280096 643200 280108
rect 643252 280096 643258 280148
rect 250722 280028 250728 280080
rect 250780 280068 250786 280080
rect 310338 280068 310344 280080
rect 250780 280040 310344 280068
rect 250780 280028 250786 280040
rect 310338 280028 310344 280040
rect 310396 280028 310402 280080
rect 612466 280028 612472 280080
rect 612524 280068 612530 280080
rect 633258 280068 633264 280080
rect 612524 280040 633264 280068
rect 612524 280028 612530 280040
rect 633258 280028 633264 280040
rect 633316 280028 633322 280080
rect 249158 279960 249164 280012
rect 249216 280000 249222 280012
rect 511634 280000 511640 280012
rect 249216 279972 511640 280000
rect 249216 279960 249222 279972
rect 511634 279960 511640 279972
rect 511692 279960 511698 280012
rect 554874 279960 554880 280012
rect 554932 280000 554938 280012
rect 646506 280000 646512 280012
rect 554932 279972 646512 280000
rect 554932 279960 554938 279972
rect 646506 279960 646512 279972
rect 646564 279960 646570 280012
rect 367930 279892 367936 279944
rect 367988 279932 367994 279944
rect 624426 279932 624432 279944
rect 367988 279904 624432 279932
rect 367988 279892 367994 279904
rect 624426 279892 624432 279904
rect 624484 279892 624490 279944
rect 211530 279824 211536 279876
rect 211588 279864 211594 279876
rect 463794 279864 463800 279876
rect 211588 279836 463800 279864
rect 211588 279824 211594 279836
rect 463794 279824 463800 279836
rect 463852 279824 463858 279876
rect 487714 279824 487720 279876
rect 487772 279864 487778 279876
rect 637674 279864 637680 279876
rect 487772 279836 637680 279864
rect 487772 279824 487778 279836
rect 637674 279824 637680 279836
rect 637732 279824 637738 279876
rect 232506 279756 232512 279808
rect 232564 279796 232570 279808
rect 473362 279796 473368 279808
rect 232564 279768 473368 279796
rect 232564 279756 232570 279768
rect 473362 279756 473368 279768
rect 473420 279756 473426 279808
rect 497282 279756 497288 279808
rect 497340 279796 497346 279808
rect 625530 279796 625536 279808
rect 497340 279768 625536 279796
rect 497340 279756 497346 279768
rect 625530 279756 625536 279768
rect 625588 279756 625594 279808
rect 252746 279688 252752 279740
rect 252804 279728 252810 279740
rect 430306 279728 430312 279740
rect 252804 279700 430312 279728
rect 252804 279688 252810 279700
rect 430306 279688 430312 279700
rect 430364 279688 430370 279740
rect 454226 279688 454232 279740
rect 454284 279728 454290 279740
rect 675210 279728 675216 279740
rect 454284 279700 675216 279728
rect 454284 279688 454290 279700
rect 675210 279688 675216 279700
rect 675268 279688 675274 279740
rect 249434 279620 249440 279672
rect 249492 279660 249498 279672
rect 415770 279660 415776 279672
rect 249492 279632 415776 279660
rect 249492 279620 249498 279632
rect 415770 279620 415776 279632
rect 415828 279620 415834 279672
rect 251550 279552 251556 279604
rect 251608 279592 251614 279604
rect 387066 279592 387072 279604
rect 251608 279564 387072 279592
rect 251608 279552 251614 279564
rect 387066 279552 387072 279564
rect 387124 279552 387130 279604
rect 251458 279484 251464 279536
rect 251516 279524 251522 279536
rect 286418 279524 286424 279536
rect 251516 279496 286424 279524
rect 251516 279484 251522 279496
rect 286418 279484 286424 279496
rect 286476 279484 286482 279536
rect 344010 279484 344016 279536
rect 344068 279524 344074 279536
rect 620010 279524 620016 279536
rect 344068 279496 620016 279524
rect 344068 279484 344074 279496
rect 620010 279484 620016 279496
rect 620068 279484 620074 279536
rect 248238 279416 248244 279468
rect 248296 279456 248302 279468
rect 377498 279456 377504 279468
rect 248296 279428 377504 279456
rect 248296 279416 248302 279428
rect 377498 279416 377504 279428
rect 377556 279416 377562 279468
rect 232322 279076 232328 279128
rect 232380 279116 232386 279128
rect 248146 279116 248152 279128
rect 232380 279088 248152 279116
rect 232380 279076 232386 279088
rect 248146 279076 248152 279088
rect 248204 279116 248210 279128
rect 248514 279116 248520 279128
rect 248204 279088 248520 279116
rect 248204 279076 248210 279088
rect 248514 279076 248520 279088
rect 248572 279076 248578 279128
rect 251918 279076 251924 279128
rect 251976 279116 251982 279128
rect 676130 279116 676136 279128
rect 251976 279088 676136 279116
rect 251976 279076 251982 279088
rect 676130 279076 676136 279088
rect 676188 279076 676194 279128
rect 252194 279008 252200 279060
rect 252252 279048 252258 279060
rect 676294 279048 676300 279060
rect 252252 279020 676300 279048
rect 252252 279008 252258 279020
rect 676294 279008 676300 279020
rect 676352 279008 676358 279060
rect 249066 278940 249072 278992
rect 249124 278980 249130 278992
rect 564442 278980 564448 278992
rect 249124 278952 564448 278980
rect 249124 278940 249130 278952
rect 564442 278940 564448 278952
rect 564500 278940 564506 278992
rect 569226 278940 569232 278992
rect 569284 278980 569290 278992
rect 619642 278980 619648 278992
rect 569284 278952 619648 278980
rect 569284 278940 569290 278952
rect 619642 278940 619648 278952
rect 619700 278940 619706 278992
rect 535738 278872 535744 278924
rect 535796 278912 535802 278924
rect 621666 278912 621672 278924
rect 535796 278884 621672 278912
rect 535796 278872 535802 278884
rect 621666 278872 621672 278884
rect 621724 278872 621730 278924
rect 251734 278804 251740 278856
rect 251792 278844 251798 278856
rect 516602 278844 516608 278856
rect 251792 278816 516608 278844
rect 251792 278804 251798 278816
rect 516602 278804 516608 278816
rect 516660 278804 516666 278856
rect 526170 278804 526176 278856
rect 526228 278844 526234 278856
rect 619734 278844 619740 278856
rect 526228 278816 619740 278844
rect 526228 278804 526234 278816
rect 619734 278804 619740 278816
rect 619792 278804 619798 278856
rect 250446 278736 250452 278788
rect 250504 278776 250510 278788
rect 502486 278776 502492 278788
rect 250504 278748 502492 278776
rect 250504 278736 250510 278748
rect 502486 278736 502492 278748
rect 502544 278736 502550 278788
rect 506850 278736 506856 278788
rect 506908 278776 506914 278788
rect 619550 278776 619556 278788
rect 506908 278748 619556 278776
rect 506908 278736 506914 278748
rect 619550 278736 619556 278748
rect 619608 278736 619614 278788
rect 249526 278668 249532 278720
rect 249584 278708 249590 278720
rect 492498 278708 492504 278720
rect 249584 278680 492504 278708
rect 249584 278668 249590 278680
rect 492498 278668 492504 278680
rect 492556 278668 492562 278720
rect 578794 278668 578800 278720
rect 578852 278708 578858 278720
rect 622954 278708 622960 278720
rect 578852 278680 622960 278708
rect 578852 278668 578858 278680
rect 622954 278668 622960 278680
rect 623012 278668 623018 278720
rect 250906 278600 250912 278652
rect 250964 278640 250970 278652
rect 382282 278640 382288 278652
rect 250964 278612 382288 278640
rect 250964 278600 250970 278612
rect 382282 278600 382288 278612
rect 382340 278600 382346 278652
rect 401418 278600 401424 278652
rect 401476 278640 401482 278652
rect 621758 278640 621764 278652
rect 401476 278612 621764 278640
rect 401476 278600 401482 278612
rect 621758 278600 621764 278612
rect 621816 278600 621822 278652
rect 248330 278532 248336 278584
rect 248388 278572 248394 278584
rect 410986 278572 410992 278584
rect 248388 278544 410992 278572
rect 248388 278532 248394 278544
rect 410986 278532 410992 278544
rect 411044 278532 411050 278584
rect 248146 278464 248152 278516
rect 248204 278504 248210 278516
rect 360570 278504 360576 278516
rect 248204 278476 360576 278504
rect 248204 278464 248210 278476
rect 360570 278464 360576 278476
rect 360628 278464 360634 278516
rect 249618 278396 249624 278448
rect 249676 278436 249682 278448
rect 315122 278436 315128 278448
rect 249676 278408 315128 278436
rect 249676 278396 249682 278408
rect 315122 278396 315128 278408
rect 315180 278396 315186 278448
rect 252838 278328 252844 278380
rect 252896 278368 252902 278380
rect 300770 278368 300776 278380
rect 252896 278340 300776 278368
rect 252896 278328 252902 278340
rect 300770 278328 300776 278340
rect 300828 278328 300834 278380
rect 251642 278260 251648 278312
rect 251700 278300 251706 278312
rect 540522 278300 540528 278312
rect 251700 278272 540528 278300
rect 251700 278260 251706 278272
rect 540522 278260 540528 278272
rect 540580 278260 540586 278312
rect 244853 278071 244905 278077
rect 449467 278072 449520 278079
rect 449467 278060 449468 278072
rect 244905 278032 449468 278060
rect 244853 278013 244905 278019
rect 449467 278020 449468 278032
rect 449467 278014 449520 278020
rect 281645 277962 281697 277968
rect 673318 277960 673370 277967
rect 281697 277921 673318 277949
rect 281645 277903 281697 277909
rect 673318 277902 673370 277908
rect 611178 276288 611184 276340
rect 611236 276328 611242 276340
rect 619090 276328 619096 276340
rect 611236 276300 619096 276328
rect 611236 276288 611242 276300
rect 619090 276288 619096 276300
rect 619148 276288 619154 276340
rect 609706 274112 609712 274164
rect 609764 274152 609770 274164
rect 620746 274152 620752 274164
rect 609764 274124 620752 274152
rect 609764 274112 609770 274124
rect 620746 274112 620752 274124
rect 620804 274112 620810 274164
rect 229838 266360 229844 266412
rect 229896 266400 229902 266412
rect 576954 266400 576960 266412
rect 229896 266372 576960 266400
rect 229896 266360 229902 266372
rect 576954 266360 576960 266372
rect 577012 266360 577018 266412
rect 339042 265272 339048 265324
rect 339100 265312 339106 265324
rect 611730 265312 611736 265324
rect 339100 265284 611736 265312
rect 339100 265272 339106 265284
rect 611730 265272 611736 265284
rect 611788 265272 611794 265324
rect 324690 264184 324696 264236
rect 324748 264224 324754 264236
rect 604554 264224 604560 264236
rect 324748 264196 604560 264224
rect 324748 264184 324754 264196
rect 604554 264184 604560 264196
rect 604612 264184 604618 264236
rect 610258 263164 610264 263216
rect 610316 263204 610322 263216
rect 611178 263204 611184 263216
rect 610316 263176 611184 263204
rect 610316 263164 610322 263176
rect 611178 263164 611184 263176
rect 611236 263164 611242 263216
rect 208034 263028 208040 263080
rect 208092 263068 208098 263080
rect 384306 263068 384312 263080
rect 208092 263040 384312 263068
rect 208092 263028 208098 263040
rect 384306 263028 384312 263040
rect 384364 263028 384370 263080
rect 391850 263028 391856 263080
rect 391908 263068 391914 263080
rect 601978 263068 601984 263080
rect 391908 263040 601984 263068
rect 391908 263028 391914 263040
rect 601978 263028 601984 263040
rect 602036 263028 602042 263080
rect 577598 262076 577604 262128
rect 577656 262116 577662 262128
rect 622862 262116 622868 262128
rect 577656 262088 622868 262116
rect 577656 262076 577662 262088
rect 622862 262076 622868 262088
rect 622920 262076 622926 262128
rect 565914 262008 565920 262060
rect 565972 262048 565978 262060
rect 621850 262048 621856 262060
rect 565972 262020 621856 262048
rect 565972 262008 565978 262020
rect 621850 262008 621856 262020
rect 621908 262008 621914 262060
rect 252010 261940 252016 261992
rect 252068 261980 252074 261992
rect 640250 261980 640256 261992
rect 252068 261952 640256 261980
rect 252068 261940 252074 261952
rect 640250 261940 640256 261952
rect 640308 261940 640314 261992
rect 583578 260852 583584 260904
rect 583636 260892 583642 260904
rect 638870 260892 638876 260904
rect 583636 260864 638876 260892
rect 583636 260852 583642 260864
rect 638870 260852 638876 260864
rect 638928 260852 638934 260904
rect 587350 260240 587356 260292
rect 587408 260280 587414 260292
rect 620010 260280 620016 260292
rect 587408 260252 620016 260280
rect 587408 260240 587414 260252
rect 620010 260240 620016 260252
rect 620068 260280 620074 260292
rect 652578 260280 652584 260292
rect 620068 260252 652584 260280
rect 620068 260240 620074 260252
rect 652578 260240 652584 260252
rect 652636 260240 652642 260292
rect 590478 260104 590484 260156
rect 590536 260144 590542 260156
rect 592686 260144 592692 260156
rect 590536 260116 592692 260144
rect 590536 260104 590542 260116
rect 592686 260104 592692 260116
rect 592744 260144 592750 260156
rect 610810 260144 610816 260156
rect 592744 260116 610816 260144
rect 592744 260104 592750 260116
rect 610810 260104 610816 260116
rect 610868 260104 610874 260156
rect 625254 260104 625260 260156
rect 625312 260144 625318 260156
rect 643378 260144 643384 260156
rect 625312 260116 643384 260144
rect 625312 260104 625318 260116
rect 643378 260104 643384 260116
rect 643436 260104 643442 260156
rect 645786 260108 647118 260136
rect 587350 260076 587356 260088
rect 557698 260048 587356 260076
rect 522214 260008 522220 260020
rect 519058 259980 522220 260008
rect 397554 259900 397560 259952
rect 397612 259940 397618 259952
rect 423866 259940 423872 259952
rect 397612 259912 423872 259940
rect 397612 259900 397618 259912
rect 423866 259900 423872 259912
rect 423924 259900 423930 259952
rect 424602 259900 424608 259952
rect 424660 259940 424666 259952
rect 456986 259940 456992 259952
rect 424660 259912 456992 259940
rect 424660 259900 424666 259912
rect 456986 259900 456992 259912
rect 457044 259940 457050 259952
rect 489554 259940 489560 259952
rect 457044 259912 489560 259940
rect 457044 259900 457050 259912
rect 489554 259900 489560 259912
rect 489612 259940 489618 259952
rect 519058 259940 519086 259980
rect 522214 259968 522220 259980
rect 522272 260008 522278 260020
rect 554782 260008 554788 260020
rect 522272 259980 554788 260008
rect 522272 259968 522278 259980
rect 554782 259968 554788 259980
rect 554840 260008 554846 260020
rect 557698 260008 557726 260048
rect 587350 260036 587356 260048
rect 587408 260036 587414 260088
rect 610442 260036 610448 260088
rect 610500 260076 610506 260088
rect 618630 260076 618636 260088
rect 610500 260048 618636 260076
rect 610500 260036 610506 260048
rect 618630 260036 618636 260048
rect 618688 260076 618694 260088
rect 618688 260048 619550 260076
rect 618688 260036 618694 260048
rect 554840 259980 557726 260008
rect 554840 259968 554846 259980
rect 610258 259960 610264 260012
rect 610316 260000 610322 260012
rect 611592 260000 611621 260002
rect 610316 259972 611621 260000
rect 610316 259960 610322 259972
rect 489612 259912 519086 259940
rect 489612 259900 489618 259912
rect 545582 259900 545588 259952
rect 545640 259940 545646 259952
rect 548434 259940 548440 259952
rect 545640 259912 548440 259940
rect 545640 259900 545646 259912
rect 548434 259900 548440 259912
rect 548492 259940 548498 259952
rect 548492 259912 549998 259940
rect 548492 259900 548498 259912
rect 395070 259832 395076 259884
rect 395128 259872 395134 259884
rect 397278 259872 397284 259884
rect 395128 259844 397284 259872
rect 395128 259832 395134 259844
rect 397278 259832 397284 259844
rect 397336 259872 397342 259884
rect 415402 259872 415408 259884
rect 397336 259844 415408 259872
rect 397336 259832 397342 259844
rect 415402 259832 415408 259844
rect 415460 259832 415466 259884
rect 423682 259832 423688 259884
rect 423740 259872 423746 259884
rect 424620 259872 424648 259900
rect 513014 259872 513020 259884
rect 423740 259844 424648 259872
rect 511330 259844 513020 259872
rect 423740 259832 423746 259844
rect 384975 259756 384981 259768
rect 382820 259696 382826 259748
rect 382878 259736 382884 259748
rect 383788 259736 384981 259756
rect 382878 259728 384981 259736
rect 382878 259708 383828 259728
rect 384975 259716 384981 259728
rect 385033 259756 385039 259768
rect 385033 259736 385528 259756
rect 388371 259736 388377 259748
rect 385033 259728 388377 259736
rect 385033 259716 385039 259728
rect 385485 259708 388377 259728
rect 382878 259696 382884 259708
rect 388371 259696 388377 259708
rect 388429 259696 388435 259748
rect 389293 259716 389299 259768
rect 389351 259756 389357 259768
rect 395420 259763 396172 259791
rect 414850 259764 414856 259816
rect 414908 259804 414914 259816
rect 418062 259804 418068 259816
rect 414908 259776 418068 259804
rect 414908 259764 414914 259776
rect 418062 259764 418068 259776
rect 418120 259764 418126 259816
rect 418272 259776 418668 259804
rect 389351 259736 389758 259756
rect 391083 259736 391875 259756
rect 395420 259736 395448 259763
rect 389351 259728 395448 259736
rect 389351 259716 389357 259728
rect 389723 259708 391115 259728
rect 391843 259708 395448 259728
rect 396144 259736 396172 259763
rect 397830 259748 397836 259760
rect 397029 259736 397836 259748
rect 396144 259720 397836 259736
rect 395523 259690 396098 259718
rect 396144 259708 397063 259720
rect 397830 259708 397836 259720
rect 397888 259708 397894 259760
rect 396144 259707 396172 259708
rect 210426 259628 210432 259680
rect 210484 259668 210490 259680
rect 383891 259668 385405 259688
rect 388868 259668 389672 259688
rect 391154 259668 391804 259688
rect 391979 259668 391985 259680
rect 210484 259660 391985 259668
rect 210484 259640 383935 259660
rect 385373 259640 388901 259660
rect 389637 259640 391191 259660
rect 391772 259640 391985 259660
rect 210484 259628 210490 259640
rect 391979 259628 391985 259640
rect 392037 259668 392043 259680
rect 395523 259668 395551 259690
rect 392037 259640 395551 259668
rect 396070 259668 396098 259690
rect 397030 259668 398030 259680
rect 418272 259668 418300 259776
rect 396070 259652 418300 259668
rect 396070 259640 397063 259652
rect 397983 259640 418300 259652
rect 418364 259708 418576 259736
rect 392037 259628 392043 259640
rect 247410 259560 247416 259612
rect 247468 259600 247474 259612
rect 383967 259600 385321 259620
rect 388947 259600 389571 259620
rect 391224 259600 391744 259620
rect 395622 259612 396020 259640
rect 395622 259600 395650 259612
rect 247468 259592 395650 259600
rect 247468 259572 384011 259592
rect 385281 259572 388979 259592
rect 389537 259572 391259 259592
rect 391716 259572 395650 259592
rect 395992 259600 396020 259612
rect 397024 259600 398019 259612
rect 418364 259600 418392 259708
rect 395992 259584 418392 259600
rect 395992 259572 397063 259584
rect 397983 259572 418392 259584
rect 247468 259560 247474 259572
rect 384490 259512 384496 259564
rect 384548 259552 384554 259564
rect 389182 259552 389188 259564
rect 384548 259532 385202 259552
rect 389017 259532 389188 259552
rect 384548 259524 389188 259532
rect 384548 259512 384554 259524
rect 385167 259504 389051 259524
rect 389182 259512 389188 259524
rect 389240 259512 389246 259564
rect 391390 259512 391396 259564
rect 391448 259552 391454 259564
rect 391448 259532 391689 259552
rect 395791 259532 395797 259556
rect 391448 259524 395797 259532
rect 391448 259512 391454 259524
rect 391655 259504 395797 259524
rect 395849 259532 395855 259556
rect 397554 259544 397560 259556
rect 397015 259532 397560 259544
rect 395849 259516 397560 259532
rect 395849 259504 397063 259516
rect 397554 259504 397560 259516
rect 397612 259504 397618 259556
rect 397670 259504 397676 259556
rect 397728 259544 397734 259556
rect 397830 259544 397836 259556
rect 397728 259516 397836 259544
rect 397728 259504 397734 259516
rect 397830 259504 397836 259516
rect 397888 259544 397894 259556
rect 418442 259552 418448 259604
rect 418500 259592 418506 259604
rect 418548 259600 418576 259708
rect 418640 259668 418668 259776
rect 421888 259746 421894 259798
rect 421946 259786 421952 259798
rect 421946 259758 422224 259786
rect 426442 259764 426448 259816
rect 426500 259804 426506 259816
rect 427730 259804 427736 259816
rect 426500 259776 427736 259804
rect 426500 259764 426506 259776
rect 427730 259764 427736 259776
rect 427788 259804 427794 259816
rect 429846 259804 429852 259816
rect 427788 259776 429852 259804
rect 427788 259764 427794 259776
rect 429846 259764 429852 259776
rect 429904 259804 429910 259816
rect 429904 259776 447878 259804
rect 454410 259784 454416 259836
rect 454468 259824 454474 259836
rect 454468 259804 454935 259824
rect 457170 259804 457176 259816
rect 454468 259796 457176 259804
rect 454468 259784 454474 259796
rect 429904 259764 429910 259776
rect 421946 259746 421952 259758
rect 422196 259736 422224 259758
rect 447850 259748 447878 259776
rect 450635 259751 451345 259779
rect 454902 259776 457176 259796
rect 457170 259764 457176 259776
rect 457228 259804 457234 259816
rect 462690 259804 462696 259816
rect 457228 259776 462696 259804
rect 457228 259764 457234 259776
rect 462690 259764 462696 259776
rect 462748 259804 462754 259816
rect 480262 259804 480268 259816
rect 462748 259776 480268 259804
rect 462748 259764 462754 259776
rect 480262 259764 480268 259776
rect 480320 259804 480326 259816
rect 483466 259804 483472 259820
rect 480320 259776 483472 259804
rect 480320 259764 480326 259776
rect 483466 259768 483472 259776
rect 483524 259804 483530 259820
rect 483524 259776 483801 259804
rect 483524 259768 483530 259776
rect 430270 259736 430276 259748
rect 422196 259708 430276 259736
rect 421595 259680 422149 259708
rect 430270 259696 430276 259708
rect 430328 259696 430334 259748
rect 447832 259696 447838 259748
rect 447890 259736 447896 259748
rect 449975 259736 449981 259748
rect 447890 259708 449981 259736
rect 447890 259696 447896 259708
rect 449975 259696 449981 259708
rect 450033 259736 450039 259748
rect 450635 259736 450663 259751
rect 450033 259708 450663 259736
rect 451317 259736 451345 259751
rect 453371 259736 453377 259748
rect 450033 259696 450039 259708
rect 450746 259683 451262 259711
rect 451317 259708 453377 259736
rect 453371 259696 453377 259708
rect 453429 259736 453435 259748
rect 453728 259736 454813 259756
rect 457644 259736 457650 259748
rect 453429 259728 457650 259736
rect 453429 259708 453773 259728
rect 454778 259708 457650 259728
rect 453429 259696 453435 259708
rect 457644 259696 457650 259708
rect 457702 259736 457708 259748
rect 458022 259736 458028 259748
rect 457702 259708 458028 259736
rect 457702 259696 457708 259708
rect 458022 259696 458028 259708
rect 458080 259736 458086 259748
rect 458872 259736 458878 259748
rect 458080 259708 458878 259736
rect 458080 259696 458086 259708
rect 458872 259696 458878 259708
rect 458930 259736 458936 259748
rect 460080 259736 460086 259748
rect 458930 259708 460086 259736
rect 458930 259696 458936 259708
rect 460080 259696 460086 259708
rect 460138 259736 460144 259748
rect 462261 259736 462267 259748
rect 460138 259708 462267 259736
rect 460138 259696 460144 259708
rect 462261 259696 462267 259708
rect 462319 259736 462325 259748
rect 480420 259736 480426 259748
rect 462319 259708 480426 259736
rect 462319 259696 462325 259708
rect 480420 259696 480426 259708
rect 480478 259736 480484 259748
rect 482575 259736 482581 259748
rect 480478 259708 482581 259736
rect 480478 259696 480484 259708
rect 482575 259696 482581 259708
rect 482633 259696 482639 259748
rect 483773 259736 483801 259776
rect 494706 259764 494712 259816
rect 494764 259804 494770 259816
rect 511330 259804 511358 259844
rect 513014 259832 513020 259844
rect 513072 259832 513078 259884
rect 522398 259832 522404 259884
rect 522456 259872 522462 259884
rect 522858 259872 522864 259884
rect 522456 259844 522864 259872
rect 522456 259832 522462 259844
rect 522858 259832 522864 259844
rect 522916 259872 522922 259884
rect 523226 259872 523232 259884
rect 522916 259844 523232 259872
rect 522916 259832 522922 259844
rect 523226 259832 523232 259844
rect 523284 259872 523290 259884
rect 524054 259872 524060 259884
rect 523284 259844 524060 259872
rect 523284 259832 523290 259844
rect 524054 259832 524060 259844
rect 524112 259872 524118 259884
rect 525250 259872 525256 259884
rect 524112 259844 525256 259872
rect 524112 259832 524118 259844
rect 525250 259832 525256 259844
rect 525308 259872 525314 259884
rect 527458 259872 527464 259884
rect 525308 259844 527464 259872
rect 525308 259832 525314 259844
rect 527458 259832 527464 259844
rect 527516 259872 527522 259884
rect 527516 259844 542270 259872
rect 527516 259832 527522 259844
rect 494764 259776 511358 259804
rect 494764 259764 494770 259776
rect 512830 259764 512836 259816
rect 512888 259764 512894 259816
rect 515422 259804 516715 259824
rect 518534 259804 518540 259816
rect 515194 259796 518540 259804
rect 515194 259776 515465 259796
rect 516673 259776 518540 259796
rect 486893 259736 486899 259748
rect 483018 259699 483700 259727
rect 483773 259708 486899 259736
rect 421595 259668 421629 259680
rect 418640 259640 421629 259668
rect 422119 259668 422149 259680
rect 423682 259668 423688 259680
rect 422119 259640 423688 259668
rect 421677 259612 422045 259640
rect 423682 259628 423688 259640
rect 423740 259628 423746 259680
rect 423850 259628 423856 259680
rect 423908 259668 423914 259680
rect 428391 259668 428397 259680
rect 423908 259640 428397 259668
rect 423908 259628 423914 259640
rect 428391 259628 428397 259640
rect 428449 259668 428455 259680
rect 450746 259668 450776 259683
rect 428449 259640 450776 259668
rect 451234 259668 451262 259683
rect 453860 259668 454736 259688
rect 456250 259668 456256 259680
rect 451234 259660 456256 259668
rect 451234 259640 453891 259660
rect 454706 259640 456256 259660
rect 428449 259628 428455 259640
rect 421677 259600 421707 259612
rect 418500 259552 418514 259592
rect 418548 259572 421707 259600
rect 422009 259600 422045 259612
rect 450822 259605 451188 259633
rect 456250 259628 456256 259640
rect 456308 259668 456314 259680
rect 460791 259668 460797 259680
rect 456308 259640 460797 259668
rect 456308 259628 456314 259640
rect 460791 259628 460797 259640
rect 460849 259668 460855 259680
rect 483018 259668 483046 259699
rect 460849 259640 483046 259668
rect 483672 259668 483700 259699
rect 486893 259696 486899 259708
rect 486951 259736 486957 259748
rect 495270 259736 495276 259748
rect 486951 259708 495276 259736
rect 486951 259696 486957 259708
rect 495270 259696 495276 259708
rect 495328 259736 495334 259748
rect 512848 259736 512876 259764
rect 515194 259748 515222 259776
rect 495328 259708 512876 259736
rect 495328 259696 495334 259708
rect 513014 259696 513020 259748
rect 513072 259736 513078 259748
rect 515176 259736 515182 259748
rect 513072 259708 515182 259736
rect 513072 259696 513078 259708
rect 515176 259696 515182 259708
rect 515234 259696 515240 259748
rect 516142 259716 516148 259768
rect 516200 259756 516206 259768
rect 518534 259764 518540 259776
rect 518592 259764 518598 259816
rect 542242 259804 542270 259844
rect 545306 259832 545312 259884
rect 545364 259872 545370 259884
rect 549970 259872 549998 259912
rect 558646 259900 558652 259952
rect 558704 259940 558710 259952
rect 586614 259940 586620 259952
rect 558704 259912 586620 259940
rect 558704 259900 558710 259912
rect 586614 259900 586620 259912
rect 586672 259900 586678 259952
rect 611592 259940 611621 259972
rect 611730 259968 611736 260020
rect 611788 260008 611794 260020
rect 617250 260008 617256 260020
rect 611788 259980 617256 260008
rect 611788 259968 611794 259980
rect 617250 259968 617256 259980
rect 617308 259968 617314 260020
rect 619522 260008 619550 260048
rect 638778 260036 638784 260088
rect 638836 260076 638842 260088
rect 645586 260076 645592 260088
rect 638836 260048 645592 260076
rect 638836 260036 638842 260048
rect 645586 260036 645592 260048
rect 645644 260076 645650 260088
rect 645786 260076 645814 260108
rect 645644 260048 645814 260076
rect 647090 260076 647118 260108
rect 653222 260076 653228 260088
rect 645644 260036 645650 260048
rect 645884 260040 647034 260068
rect 647090 260048 653228 260076
rect 643010 260008 643016 260020
rect 619522 259980 643016 260008
rect 643010 259968 643016 259980
rect 643068 260008 643074 260020
rect 645884 260008 645912 260040
rect 643068 259980 645912 260008
rect 647006 260008 647034 260040
rect 653222 260036 653228 260048
rect 653280 260036 653286 260088
rect 643068 259968 643074 259980
rect 645960 259972 646970 260000
rect 647006 259980 650462 260008
rect 613018 259940 613024 259952
rect 611592 259912 613024 259940
rect 610357 259901 611313 259902
rect 551194 259872 551200 259884
rect 545364 259844 549860 259872
rect 549970 259844 551200 259872
rect 545364 259832 545370 259844
rect 545582 259804 545588 259816
rect 542242 259776 545588 259804
rect 545582 259764 545588 259776
rect 545640 259764 545646 259816
rect 549832 259804 549860 259844
rect 551194 259832 551200 259844
rect 551252 259832 551258 259884
rect 555426 259872 555432 259884
rect 553696 259844 555432 259872
rect 553494 259804 553500 259816
rect 549832 259776 553500 259804
rect 553494 259764 553500 259776
rect 553552 259764 553558 259816
rect 516200 259736 516628 259756
rect 519500 259736 519506 259748
rect 516200 259728 519506 259736
rect 516200 259716 516206 259728
rect 516600 259708 519506 259728
rect 519500 259696 519506 259708
rect 519558 259736 519564 259748
rect 527872 259736 527878 259748
rect 519558 259708 527878 259736
rect 519558 259696 519564 259708
rect 527872 259696 527878 259708
rect 527930 259736 527936 259748
rect 545030 259736 545036 259748
rect 527930 259708 545036 259736
rect 527930 259696 527936 259708
rect 545030 259696 545036 259708
rect 545088 259736 545094 259748
rect 547775 259736 547781 259748
rect 545088 259708 547781 259736
rect 545088 259696 545094 259708
rect 547775 259696 547781 259708
rect 547833 259736 547839 259748
rect 548150 259736 548950 259756
rect 552093 259736 552099 259748
rect 547833 259728 552099 259736
rect 547833 259708 548183 259728
rect 548913 259708 552099 259728
rect 547833 259696 547839 259708
rect 552093 259696 552099 259708
rect 552151 259736 552157 259748
rect 553696 259736 553724 259844
rect 555426 259832 555432 259844
rect 555484 259872 555490 259884
rect 578058 259872 578064 259884
rect 555484 259844 578064 259872
rect 555484 259832 555490 259844
rect 578058 259832 578064 259844
rect 578116 259872 578122 259884
rect 580818 259872 580824 259884
rect 578116 259844 580824 259872
rect 578116 259832 578122 259844
rect 580818 259832 580824 259844
rect 580876 259832 580882 259884
rect 585284 259864 585312 259865
rect 583709 259836 585312 259864
rect 558646 259804 558652 259816
rect 552151 259708 553724 259736
rect 554064 259776 558652 259804
rect 552151 259696 552157 259708
rect 488850 259668 488856 259680
rect 460849 259628 460855 259640
rect 483292 259622 483615 259650
rect 483672 259640 488856 259668
rect 488850 259628 488856 259640
rect 488908 259668 488914 259680
rect 493391 259668 493397 259680
rect 488908 259640 493397 259668
rect 488908 259628 488914 259640
rect 493391 259628 493397 259640
rect 493449 259668 493455 259680
rect 515632 259668 516550 259688
rect 521450 259668 521456 259680
rect 493449 259660 521456 259668
rect 493449 259640 515675 259660
rect 516515 259640 521456 259660
rect 493449 259628 493455 259640
rect 521450 259628 521456 259640
rect 521508 259668 521514 259680
rect 525986 259668 525992 259680
rect 521508 259640 525992 259668
rect 521508 259628 521514 259640
rect 525986 259628 525992 259640
rect 526044 259668 526050 259680
rect 548221 259668 548866 259688
rect 554064 259680 554092 259776
rect 558646 259764 558652 259776
rect 558704 259764 558710 259816
rect 577782 259764 577788 259816
rect 577840 259804 577846 259816
rect 583709 259804 583737 259836
rect 577840 259776 583737 259804
rect 585284 259804 585312 259836
rect 601978 259832 601984 259884
rect 602036 259872 602042 259884
rect 610353 259874 611313 259901
rect 613018 259900 613024 259912
rect 613076 259940 613082 259952
rect 620654 259940 620660 259952
rect 613076 259912 620660 259940
rect 613076 259900 613082 259912
rect 620654 259900 620660 259912
rect 620712 259900 620718 259952
rect 642090 259900 642096 259952
rect 642148 259940 642154 259952
rect 645960 259940 645988 259972
rect 642148 259912 645988 259940
rect 646942 259940 646970 259972
rect 649910 259940 649916 259952
rect 642148 259900 642154 259912
rect 646044 259904 646902 259932
rect 646942 259912 649916 259940
rect 610353 259872 610381 259874
rect 602036 259844 610381 259872
rect 611285 259872 611313 259874
rect 616330 259872 616336 259884
rect 611285 259844 616336 259872
rect 602036 259832 602042 259844
rect 610463 259833 611239 259834
rect 586062 259804 586068 259816
rect 584682 259786 584688 259798
rect 577840 259764 577846 259776
rect 584010 259758 584688 259786
rect 556671 259696 556677 259748
rect 556729 259736 556735 259748
rect 565914 259736 565920 259748
rect 556729 259708 565920 259736
rect 556729 259696 556735 259708
rect 565914 259696 565920 259708
rect 565972 259696 565978 259748
rect 576954 259696 576960 259748
rect 577012 259736 577018 259748
rect 584010 259736 584038 259758
rect 584682 259746 584688 259758
rect 584740 259746 584746 259798
rect 585284 259776 586068 259804
rect 586062 259764 586068 259776
rect 586120 259764 586126 259816
rect 604554 259764 604560 259816
rect 604612 259804 604618 259816
rect 610459 259806 611239 259833
rect 616330 259832 616336 259844
rect 616388 259832 616394 259884
rect 640986 259832 640992 259884
rect 641044 259872 641050 259884
rect 646044 259872 646072 259904
rect 641044 259844 646072 259872
rect 646874 259872 646902 259904
rect 649910 259900 649916 259912
rect 649968 259900 649974 259952
rect 648990 259872 648996 259884
rect 641044 259832 641050 259844
rect 646128 259836 646840 259864
rect 646874 259844 648996 259872
rect 610459 259804 610487 259806
rect 604612 259776 610487 259804
rect 611209 259804 611239 259806
rect 621850 259804 621856 259816
rect 611209 259776 621856 259804
rect 604612 259764 604618 259776
rect 577012 259708 584038 259736
rect 585154 259708 585182 259709
rect 577012 259696 577018 259708
rect 584155 259680 585182 259708
rect 586614 259696 586620 259748
rect 586672 259736 586678 259748
rect 591191 259736 591197 259748
rect 586672 259708 591197 259736
rect 586672 259696 586678 259708
rect 591191 259696 591197 259708
rect 591249 259736 591255 259748
rect 610546 259738 611164 259766
rect 621850 259764 621856 259776
rect 621908 259764 621914 259816
rect 638870 259764 638876 259816
rect 638928 259804 638934 259816
rect 646128 259804 646156 259836
rect 638928 259776 646156 259804
rect 646812 259804 646840 259836
rect 648990 259832 648996 259844
rect 649048 259832 649054 259884
rect 650434 259872 650462 259980
rect 651290 259872 651296 259884
rect 650434 259844 651296 259872
rect 651290 259832 651296 259844
rect 651348 259872 651354 259884
rect 657822 259872 657828 259884
rect 651348 259844 657828 259872
rect 651348 259832 651354 259844
rect 657822 259832 657828 259844
rect 657880 259832 657886 259884
rect 638928 259764 638934 259776
rect 646212 259768 646758 259796
rect 646812 259776 652625 259804
rect 610546 259736 610574 259738
rect 591249 259708 610574 259736
rect 611134 259736 611164 259738
rect 619250 259736 619256 259748
rect 611134 259708 619256 259736
rect 591249 259696 591255 259708
rect 554046 259668 554052 259680
rect 526044 259660 554052 259668
rect 526044 259640 548252 259660
rect 548833 259640 554052 259660
rect 526044 259628 526050 259640
rect 554046 259628 554052 259640
rect 554104 259628 554110 259680
rect 554992 259628 554998 259680
rect 555050 259668 555056 259680
rect 555822 259668 555828 259680
rect 555050 259640 555828 259668
rect 555050 259628 555056 259640
rect 555822 259628 555828 259640
rect 555880 259668 555886 259680
rect 557880 259668 557886 259680
rect 555880 259640 557886 259668
rect 555880 259628 555886 259640
rect 557880 259628 557886 259640
rect 557938 259668 557944 259680
rect 560061 259668 560067 259680
rect 557938 259640 560067 259668
rect 557938 259628 557944 259640
rect 560061 259628 560067 259640
rect 560119 259668 560125 259680
rect 560470 259668 560476 259680
rect 560119 259640 560476 259668
rect 560119 259628 560125 259640
rect 560470 259628 560476 259640
rect 560528 259668 560534 259680
rect 578220 259668 578226 259680
rect 560528 259640 578226 259668
rect 560528 259628 560534 259640
rect 578220 259628 578226 259640
rect 578278 259668 578284 259680
rect 580375 259668 580381 259680
rect 578278 259640 580381 259668
rect 578278 259628 578284 259640
rect 580375 259628 580381 259640
rect 580433 259628 580439 259680
rect 580488 259632 580818 259660
rect 450822 259600 450850 259605
rect 422009 259572 450850 259600
rect 451160 259600 451188 259605
rect 453932 259600 454675 259620
rect 483292 259600 483320 259622
rect 451160 259592 483320 259600
rect 451160 259572 453967 259592
rect 454642 259572 483320 259592
rect 483587 259600 483615 259622
rect 515702 259600 516488 259620
rect 548283 259600 548788 259620
rect 580488 259600 580516 259632
rect 483587 259592 580516 259600
rect 483587 259572 515735 259592
rect 516425 259572 548326 259592
rect 548751 259572 580516 259592
rect 580790 259600 580818 259632
rect 583771 259628 583777 259680
rect 583829 259668 583835 259680
rect 584155 259668 584183 259680
rect 583829 259640 584183 259668
rect 585154 259668 585182 259680
rect 593070 259668 593076 259680
rect 585071 259640 585099 259641
rect 585154 259640 593076 259668
rect 583829 259628 583835 259640
rect 584258 259612 585099 259640
rect 593070 259628 593076 259640
rect 593128 259668 593134 259680
rect 610626 259668 610632 259680
rect 593128 259640 610632 259668
rect 593128 259628 593134 259640
rect 610626 259628 610632 259640
rect 610684 259668 610690 259680
rect 610745 259670 611082 259698
rect 619250 259696 619256 259708
rect 619308 259736 619314 259748
rect 623782 259736 623788 259748
rect 619308 259708 623788 259736
rect 619308 259696 619314 259708
rect 623782 259696 623788 259708
rect 623840 259736 623846 259748
rect 646212 259736 646240 259768
rect 623840 259708 646240 259736
rect 646456 259728 646462 259740
rect 623840 259696 623846 259708
rect 646276 259700 646462 259728
rect 610745 259668 610773 259670
rect 610684 259640 610773 259668
rect 611052 259668 611082 259670
rect 615339 259668 615822 259679
rect 611052 259650 632568 259668
rect 611052 259640 615375 259650
rect 615789 259640 632568 259650
rect 610684 259628 610690 259640
rect 610816 259629 611024 259630
rect 584258 259600 584286 259612
rect 451160 259570 451188 259572
rect 421750 259552 421756 259564
rect 397888 259532 398016 259544
rect 418462 259532 418514 259552
rect 421747 259532 421756 259552
rect 397888 259516 403166 259532
rect 397888 259504 397894 259516
rect 397983 259504 403166 259516
rect 385862 259471 385914 259504
rect 385874 259470 385902 259471
rect 403138 259328 403166 259504
rect 418462 259512 421756 259532
rect 421808 259512 421814 259564
rect 418462 259504 421792 259512
rect 418462 259471 418514 259504
rect 431198 259492 431204 259544
rect 431256 259532 431262 259544
rect 446314 259532 446320 259544
rect 431256 259504 446320 259532
rect 431256 259492 431262 259504
rect 446314 259492 446320 259504
rect 446372 259492 446378 259544
rect 451006 259532 451012 259565
rect 450886 259513 451012 259532
rect 451064 259532 451070 259565
rect 454134 259552 454140 259564
rect 453994 259532 454140 259552
rect 451064 259524 454140 259532
rect 451064 259513 454030 259524
rect 450886 259504 454030 259513
rect 454134 259512 454140 259524
rect 454192 259512 454198 259564
rect 483457 259512 483463 259564
rect 483515 259512 483521 259564
rect 516142 259552 516148 259564
rect 516068 259551 516148 259552
rect 516062 259524 516148 259551
rect 418474 259470 418502 259471
rect 450886 259470 450914 259504
rect 483462 259448 483514 259512
rect 516062 259448 516114 259524
rect 516142 259512 516148 259524
rect 516200 259512 516206 259564
rect 548434 259512 548440 259564
rect 548492 259552 548498 259564
rect 548492 259548 548572 259552
rect 548492 259524 548714 259548
rect 548492 259512 548498 259524
rect 548544 259520 548714 259524
rect 580602 259522 580608 259574
rect 580660 259562 580666 259574
rect 580790 259572 584286 259600
rect 585071 259600 585099 259612
rect 610809 259602 611024 259629
rect 610809 259600 610837 259602
rect 584498 259562 584504 259574
rect 580660 259534 580751 259562
rect 580660 259522 580666 259534
rect 580723 259532 580751 259534
rect 584396 259534 584504 259562
rect 584396 259532 584424 259534
rect 548662 259446 548714 259520
rect 580723 259505 584424 259532
rect 584498 259522 584504 259534
rect 584556 259522 584562 259574
rect 585071 259572 610837 259600
rect 610996 259600 611024 259602
rect 615422 259600 615738 259622
rect 632540 259612 632568 259640
rect 643378 259628 643384 259680
rect 643436 259668 643442 259680
rect 646276 259668 646304 259700
rect 646456 259688 646462 259700
rect 646514 259728 646520 259740
rect 646730 259736 646758 259768
rect 651850 259736 651856 259748
rect 646514 259700 646686 259728
rect 646730 259708 651856 259736
rect 646514 259688 646520 259700
rect 643436 259640 646304 259668
rect 646658 259668 646686 259700
rect 651850 259696 651856 259708
rect 651908 259696 651914 259748
rect 652597 259736 652625 259776
rect 654471 259736 654477 259748
rect 652597 259708 654477 259736
rect 654471 259696 654477 259708
rect 654529 259696 654535 259748
rect 659754 259736 659760 259748
rect 657734 259708 659760 259736
rect 657734 259680 657762 259708
rect 659754 259696 659760 259708
rect 659812 259696 659818 259748
rect 649634 259668 649640 259680
rect 643436 259628 643442 259640
rect 646348 259632 646626 259660
rect 646658 259640 649640 259668
rect 625668 259600 625674 259612
rect 610996 259593 625674 259600
rect 610996 259572 615451 259593
rect 615696 259572 625674 259593
rect 610902 259512 610908 259564
rect 610960 259532 610966 259564
rect 615594 259552 615600 259564
rect 615501 259532 615600 259552
rect 610960 259524 615600 259532
rect 610960 259512 615531 259524
rect 615594 259512 615600 259524
rect 615652 259512 615658 259564
rect 625668 259560 625674 259572
rect 625726 259560 625732 259612
rect 627738 259560 627744 259612
rect 627796 259600 627802 259612
rect 627796 259572 631694 259600
rect 627796 259560 627802 259572
rect 631666 259532 631694 259572
rect 632522 259560 632528 259612
rect 632580 259560 632586 259612
rect 646348 259600 646376 259632
rect 639394 259572 646376 259600
rect 646598 259600 646626 259632
rect 649634 259628 649640 259640
rect 649692 259668 649698 259680
rect 652792 259668 652798 259680
rect 649692 259640 652798 259668
rect 649692 259628 649698 259640
rect 652792 259628 652798 259640
rect 652850 259668 652856 259680
rect 653622 259668 653628 259680
rect 652850 259640 653628 259668
rect 652850 259628 652856 259640
rect 653622 259628 653628 259640
rect 653680 259668 653686 259680
rect 655680 259668 655686 259680
rect 653680 259640 655686 259668
rect 653680 259628 653686 259640
rect 655680 259628 655686 259640
rect 655738 259668 655744 259680
rect 657716 259668 657722 259680
rect 655738 259640 657722 259668
rect 655738 259628 655744 259640
rect 657716 259628 657722 259640
rect 657774 259628 657780 259680
rect 657822 259628 657828 259680
rect 657880 259668 657886 259680
rect 676038 259668 676044 259680
rect 657880 259640 676044 259668
rect 657880 259628 657886 259640
rect 676038 259628 676044 259640
rect 676096 259628 676102 259680
rect 658270 259600 658276 259612
rect 639394 259532 639422 259572
rect 646456 259540 646462 259592
rect 646514 259540 646520 259592
rect 646598 259572 658276 259600
rect 658270 259560 658276 259572
rect 658328 259560 658334 259612
rect 580723 259504 584421 259505
rect 610936 259504 615531 259512
rect 631666 259504 639422 259532
rect 581262 259448 581314 259504
rect 613862 259448 613914 259504
rect 646474 259470 646502 259540
rect 414850 259328 414856 259340
rect 403138 259300 414856 259328
rect 414850 259288 414856 259300
rect 414908 259288 414914 259340
<< via1 >>
rect 351826 729372 351878 729424
rect 353860 729372 353912 729424
rect 355920 729372 355972 729424
rect 356750 729372 356802 729424
rect 361036 729372 361088 729424
rect 366122 729372 366174 729424
rect 379022 729372 379074 729424
rect 381062 729372 381114 729424
rect 383120 729372 383172 729424
rect 383950 729372 384002 729424
rect 386980 729372 387032 729424
rect 393328 729372 393380 729424
rect 406392 729372 406444 729424
rect 408048 729372 408100 729424
rect 410118 729372 410170 729424
rect 414304 729372 414356 729424
rect 420284 729372 420336 729424
rect 433226 729372 433278 729424
rect 435262 729372 435314 729424
rect 437320 729372 437372 729424
rect 438150 729372 438202 729424
rect 441260 729372 441312 729424
rect 447516 729372 447568 729424
rect 460426 729372 460478 729424
rect 462466 729372 462518 729424
rect 464520 729372 464572 729424
rect 465364 729372 465416 729424
rect 468584 729372 468636 729424
rect 474748 729372 474800 729424
rect 487352 729372 487404 729424
rect 489462 729372 489514 729424
rect 491520 729372 491572 729424
rect 492350 729372 492402 729424
rect 495448 729372 495500 729424
rect 501722 729372 501774 729424
rect 514626 729372 514678 729424
rect 516662 729372 516714 729424
rect 518724 729372 518776 729424
rect 519552 729372 519604 729424
rect 522680 729372 522732 729424
rect 528936 729372 528988 729424
rect 541908 729372 541960 729424
rect 543862 729372 543914 729424
rect 545910 729372 545962 729424
rect 546738 729372 546790 729424
rect 553040 729372 553092 729424
rect 556122 729372 556174 729424
rect 570336 729372 570388 729424
rect 575028 729440 575080 729492
rect 573510 729372 573562 729424
rect 573950 729372 574002 729424
rect 577052 729372 577104 729424
rect 581167 729372 581219 729424
rect 583308 729372 583360 729424
rect 594164 729372 594216 729424
rect 595881 729372 595933 729424
rect 380356 729304 380408 729356
rect 384864 729304 384916 729356
rect 434551 729304 434603 729356
rect 439144 729304 439196 729356
rect 488751 729304 488803 729356
rect 493424 729304 493476 729356
rect 515964 729304 516016 729356
rect 520472 729304 520524 729356
rect 522588 729304 522640 729356
rect 523370 729304 523422 729356
rect 352388 729236 352440 729288
rect 353151 729236 353203 729288
rect 431876 729236 431928 729288
rect 432672 729236 432724 729288
rect 516884 729236 516936 729288
rect 517871 729236 517923 729288
rect 519184 729236 519236 729288
rect 526767 729304 526819 729356
rect 543151 729304 543203 729356
rect 547704 729304 547756 729356
rect 568956 729304 569008 729356
rect 571062 729304 571114 729356
rect 572268 729304 572320 729356
rect 573120 729304 573172 729356
rect 597351 729372 597403 729424
rect 601892 729372 601944 729424
rect 604771 729372 604823 729424
rect 624432 729430 624484 729482
rect 629216 729440 629268 729492
rect 610448 729372 610500 729424
rect 623226 729372 623278 729424
rect 625262 729372 625314 729424
rect 626471 729372 626523 729424
rect 627330 729372 627382 729424
rect 627698 729372 627750 729424
rect 628158 729372 628210 729424
rect 631240 729372 631292 729424
rect 635380 729372 635432 729424
rect 637496 729372 637548 729424
rect 650192 729372 650244 729424
rect 650422 729372 650474 729424
rect 652462 729372 652514 729424
rect 654884 729372 654936 729424
rect 598062 729304 598114 729356
rect 600120 729304 600172 729356
rect 600512 729304 600564 729356
rect 603849 729304 603901 729356
rect 608167 729304 608219 729356
rect 651756 729304 651808 729356
rect 656264 729304 656316 729356
rect 659171 729372 659223 729424
rect 664728 729372 664780 729424
rect 662567 729304 662619 729356
rect 598580 729236 598632 729288
rect 599270 729236 599322 729288
rect 600950 729236 601002 729288
rect 553316 729100 553368 729152
rect 553960 729100 554012 729152
rect 465548 729032 465600 729084
rect 492688 729032 492740 729084
rect 529120 729032 529172 729084
rect 554696 729032 554748 729084
rect 555524 729032 555576 729084
rect 556536 729032 556588 729084
rect 557088 729032 557140 729084
rect 602536 729032 602588 729084
rect 610724 729032 610776 729084
rect 250912 728964 250964 729016
rect 463616 728964 463668 729016
rect 474932 728964 474984 729016
rect 500416 728964 500468 729016
rect 522496 728964 522548 729016
rect 619556 728964 619608 729016
rect 360944 728896 360996 728948
rect 568864 728896 568916 728948
rect 576500 728896 576552 728948
rect 631148 728896 631200 728948
rect 356344 728828 356396 728880
rect 363428 728828 363480 728880
rect 363980 728828 364032 728880
rect 366096 728828 366148 728880
rect 378884 728828 378936 728880
rect 393328 728828 393380 728880
rect 405748 728828 405800 728880
rect 420284 728828 420336 728880
rect 433072 728828 433124 728880
rect 447516 728828 447568 728880
rect 460304 728828 460356 728880
rect 463984 728828 464036 728880
rect 464904 728828 464956 728880
rect 472264 728828 472316 728880
rect 474748 728828 474800 728880
rect 487352 728828 487404 728880
rect 501704 728828 501756 728880
rect 514492 728828 514544 728880
rect 358184 728760 358236 728812
rect 366464 728760 366516 728812
rect 385508 728760 385560 728812
rect 393604 728760 393656 728812
rect 412464 728760 412516 728812
rect 420744 728760 420796 728812
rect 439604 728760 439656 728812
rect 447792 728760 447844 728812
rect 466928 728760 466980 728812
rect 475208 728760 475260 728812
rect 493884 728760 493936 728812
rect 502164 728760 502216 728812
rect 521392 728828 521444 728880
rect 529304 728828 529356 728880
rect 548256 728828 548308 728880
rect 555524 728828 555576 728880
rect 556260 728828 556312 728880
rect 568496 728828 568548 728880
rect 577420 728828 577472 728880
rect 583308 728828 583360 728880
rect 594164 728828 594216 728880
rect 611460 728828 611512 728880
rect 622684 728828 622736 728880
rect 631976 728828 632028 728880
rect 528936 728760 528988 728812
rect 541356 728760 541408 728812
rect 547704 728760 547756 728812
rect 570336 728760 570388 728812
rect 577604 728760 577656 728812
rect 583584 728760 583636 728812
rect 600512 728760 600564 728812
rect 610448 728760 610500 728812
rect 623052 728760 623104 728812
rect 637680 728760 637732 728812
rect 654884 728760 654936 728812
rect 353124 728692 353176 728744
rect 357632 728692 357684 728744
rect 380356 728692 380408 728744
rect 384864 728692 384916 728744
rect 407036 728692 407088 728744
rect 411912 728692 411964 728744
rect 434544 728692 434596 728744
rect 439144 728692 439196 728744
rect 461776 728692 461828 728744
rect 466284 728692 466336 728744
rect 488732 728692 488784 728744
rect 493424 728692 493476 728744
rect 515964 728692 516016 728744
rect 520472 728692 520524 728744
rect 543104 728692 543156 728744
rect 546968 728692 547020 728744
rect 287712 728420 287764 728472
rect 356988 728624 357040 728676
rect 384036 728624 384088 728676
rect 411176 728624 411228 728676
rect 438316 728624 438368 728676
rect 465548 728624 465600 728676
rect 500416 728624 500468 728676
rect 501612 728624 501664 728676
rect 529120 728624 529172 728676
rect 556168 728624 556220 728676
rect 568956 728624 569008 728676
rect 574936 728692 574988 728744
rect 597292 728692 597344 728744
rect 601892 728692 601944 728744
rect 624524 728692 624576 728744
rect 574200 728624 574252 728676
rect 601156 728624 601208 728676
rect 628388 728692 628440 728744
rect 655436 728692 655488 728744
rect 637496 728624 637548 728676
rect 649548 728624 649600 728676
rect 654884 728624 654936 728676
rect 368028 728556 368080 728608
rect 392224 728556 392276 728608
rect 420192 728556 420244 728608
rect 447700 728556 447752 728608
rect 474932 728556 474984 728608
rect 492688 728556 492740 728608
rect 519644 728556 519696 728608
rect 546968 728556 547020 728608
rect 550464 728556 550516 728608
rect 621764 728556 621816 728608
rect 664728 728556 664780 728608
rect 675952 728556 676004 728608
rect 468308 728488 468360 728540
rect 383392 728420 383444 728472
rect 391120 728420 391172 728472
rect 410716 728420 410768 728472
rect 417524 728420 417576 728472
rect 418168 728420 418220 728472
rect 437488 728420 437540 728472
rect 445308 728420 445360 728472
rect 491952 728420 492004 728472
rect 499588 728420 499640 728472
rect 629400 728488 629452 728540
rect 651756 728488 651808 728540
rect 546324 728420 546376 728472
rect 553316 728420 553368 728472
rect 575856 728420 575908 728472
rect 583676 728420 583728 728472
rect 656264 728420 656316 728472
rect 675860 728420 675912 728472
rect 597936 728352 597988 728404
rect 335828 728284 335880 728336
rect 441996 728284 442048 728336
rect 476404 728284 476456 728336
rect 610080 728284 610132 728336
rect 436384 728216 436436 728268
rect 600144 728216 600196 728268
rect 414672 728148 414724 728200
rect 584688 728148 584740 728200
rect 658248 728194 658300 728246
rect 673124 728192 673176 728244
rect 409244 728080 409296 728132
rect 600236 728080 600288 728132
rect 394524 728012 394576 728064
rect 589104 728012 589156 728064
rect 388084 727944 388136 727996
rect 600328 727944 600380 727996
rect 378792 727876 378844 727928
rect 593520 727876 593572 727928
rect 367660 727808 367712 727860
rect 585608 727808 585660 727860
rect 499588 726856 499640 726908
rect 594624 726856 594676 726908
rect 491032 726788 491084 726840
rect 596832 726788 596884 726840
rect 382288 726720 382340 726772
rect 569876 726720 569928 726772
rect 584688 726720 584740 726772
rect 595728 726720 595780 726772
rect 568864 725700 568916 725752
rect 583584 725700 583636 725752
rect 246312 725632 246364 725684
rect 578432 725632 578484 725684
rect 246817 725452 246869 725504
rect 649298 725440 649350 725492
rect 448068 724544 448120 724596
rect 464536 724544 464588 724596
rect 583584 724136 583636 724188
rect 588000 724136 588052 724188
rect 585608 723456 585660 723508
rect 594624 723456 594676 723508
rect 607320 723456 607372 723508
rect 599040 723388 599092 723440
rect 593520 722640 593572 722692
rect 594716 722640 594768 722692
rect 468308 722300 468360 722352
rect 468860 722300 468912 722352
rect 589104 722232 589156 722284
rect 594624 722232 594676 722284
rect 600236 722096 600288 722148
rect 602352 722096 602404 722148
rect 596832 721416 596884 721468
rect 603732 721416 603784 721468
rect 600328 721280 600380 721332
rect 604560 721280 604612 721332
rect 652676 721212 652728 721264
rect 653412 721212 653464 721264
rect 595728 720600 595780 720652
rect 596832 720600 596884 720652
rect 610080 720124 610132 720176
rect 616704 720124 616756 720176
rect 607320 720056 607372 720108
rect 613484 720056 613536 720108
rect 359012 719036 359064 719088
rect 359748 719036 359800 719088
rect 363428 719036 363480 719088
rect 575396 719036 575448 719088
rect 597936 719036 597988 719088
rect 605848 719036 605900 719088
rect 485972 718832 486024 718884
rect 486524 718832 486576 718884
rect 605848 717880 605900 717932
rect 613392 717880 613444 717932
rect 603732 716792 603784 716844
rect 608976 716792 609028 716844
rect 464536 715704 464588 715756
rect 468768 715704 468820 715756
rect 208132 714616 208184 714668
rect 209972 714616 210024 714668
rect 351376 714616 351428 714668
rect 596832 714480 596884 714532
rect 597936 714480 597988 714532
rect 600144 713528 600196 713580
rect 604836 713528 604888 713580
rect 613484 713528 613536 713580
rect 614588 713528 614640 713580
rect 599040 713460 599092 713512
rect 606768 713460 606820 713512
rect 602352 712712 602404 712764
rect 604652 712712 604704 712764
rect 594716 712576 594768 712628
rect 600144 712576 600196 712628
rect 208132 711284 208184 711336
rect 365636 711284 365688 711336
rect 468768 711284 468820 711336
rect 478704 711284 478756 711336
rect 588000 711284 588052 711336
rect 604744 711284 604796 711336
rect 594624 710264 594676 710316
rect 598028 710264 598080 710316
rect 600144 708292 600196 708344
rect 602352 708292 602404 708344
rect 608976 708292 609028 708344
rect 611184 708292 611236 708344
rect 320740 707952 320792 708004
rect 595268 707952 595320 708004
rect 604744 707272 604796 707324
rect 605848 707272 605900 707324
rect 606768 707000 606820 707052
rect 608056 707000 608108 707052
rect 604652 706320 604704 706372
rect 607872 706320 607924 706372
rect 351284 705776 351336 705828
rect 512468 705776 512520 705828
rect 344660 704688 344712 704740
rect 541264 704688 541316 704740
rect 257904 703668 257956 703720
rect 354596 703668 354648 703720
rect 354688 703532 354740 703584
rect 513572 703532 513624 703584
rect 675952 702512 676004 702564
rect 676228 702512 676280 702564
rect 598028 702444 598080 702496
rect 605664 702444 605716 702496
rect 646512 701968 646564 702020
rect 676044 701968 676096 702020
rect 323040 701356 323092 701408
rect 383392 701356 383444 701408
rect 675860 701084 675912 701136
rect 676320 701084 676372 701136
rect 605848 701016 605900 701068
rect 607964 701016 608016 701068
rect 604836 700472 604888 700524
rect 610080 700472 610132 700524
rect 597936 700404 597988 700456
rect 600144 700404 600196 700456
rect 605664 700336 605716 700388
rect 611276 700336 611328 700388
rect 248980 700268 249032 700320
rect 386612 700268 386664 700320
rect 614588 699996 614640 700048
rect 615600 699996 615652 700048
rect 613392 699860 613444 699912
rect 614496 699860 614548 699912
rect 321108 699792 321160 699844
rect 358736 699792 358788 699844
rect 604560 699792 604612 699844
rect 605664 699792 605716 699844
rect 288724 699724 288776 699776
rect 384956 699724 385008 699776
rect 255696 699520 255748 699572
rect 308136 699520 308188 699572
rect 287252 699452 287304 699504
rect 299856 699452 299908 699504
rect 302616 699452 302668 699504
rect 329664 699452 329716 699504
rect 250176 699384 250228 699436
rect 301144 699384 301196 699436
rect 303904 699384 303956 699436
rect 321568 699384 321620 699436
rect 210432 699316 210484 699368
rect 309424 699316 309476 699368
rect 317704 699316 317756 699368
rect 324788 699316 324840 699368
rect 288632 699248 288684 699300
rect 330768 699248 330820 699300
rect 289092 699180 289144 699232
rect 361772 699180 361824 699232
rect 249624 699112 249676 699164
rect 292864 699112 292916 699164
rect 321844 699112 321896 699164
rect 249532 699044 249584 699096
rect 295624 699044 295676 699096
rect 297280 699044 297332 699096
rect 322028 699044 322080 699096
rect 294980 698976 295032 699028
rect 301788 698976 301840 699028
rect 249348 698908 249400 698960
rect 305560 698976 305612 699028
rect 328560 698976 328612 699028
rect 306664 698908 306716 698960
rect 316600 698908 316652 698960
rect 596832 698908 596884 698960
rect 250636 698840 250688 698892
rect 301696 698840 301748 698892
rect 301788 698840 301840 698892
rect 306848 698840 306900 698892
rect 313656 698840 313708 698892
rect 320648 698840 320700 698892
rect 361680 698840 361732 698892
rect 474288 698772 474340 698824
rect 251280 698704 251332 698756
rect 314824 698702 314876 698754
rect 321200 698704 321252 698756
rect 576960 698704 577012 698756
rect 654240 698636 654292 698688
rect 676320 698704 676372 698756
rect 323684 698092 323736 698144
rect 390016 698092 390068 698144
rect 321568 698024 321620 698076
rect 508144 698024 508196 698076
rect 675952 697948 676004 698000
rect 676326 697950 676378 698002
rect 675676 697480 675728 697532
rect 676044 697480 676096 697532
rect 478704 696936 478756 696988
rect 489744 696936 489796 696988
rect 664820 696936 664872 696988
rect 667488 696936 667540 696988
rect 675584 696528 675636 696580
rect 675860 696528 675912 696580
rect 676320 696528 676372 696580
rect 654884 696460 654936 696512
rect 676044 696460 676096 696512
rect 675768 696052 675820 696104
rect 676044 696052 676096 696104
rect 320556 695780 320608 695832
rect 321200 695780 321252 695832
rect 557088 695372 557140 695424
rect 675860 695372 675912 695424
rect 676044 695372 676096 695424
rect 384956 695304 385008 695356
rect 387164 695304 387216 695356
rect 619648 695304 619700 695356
rect 320648 695100 320700 695152
rect 322580 695100 322632 695152
rect 321936 694760 321988 694812
rect 370788 694760 370840 694812
rect 361864 694692 361916 694744
rect 376676 694692 376728 694744
rect 358736 694624 358788 694676
rect 372812 694624 372864 694676
rect 381276 694624 381328 694676
rect 460580 694624 460632 694676
rect 321844 694556 321896 694608
rect 388820 694556 388872 694608
rect 321016 694488 321068 694540
rect 375204 694488 375256 694540
rect 625076 694488 625128 694540
rect 675676 694488 675728 694540
rect 676136 694488 676188 694540
rect 624432 694216 624484 694268
rect 676044 694216 676096 694268
rect 675860 694012 675912 694064
rect 676136 694012 676188 694064
rect 208132 693944 208184 693996
rect 208316 693944 208368 693996
rect 324788 693128 324840 693180
rect 356988 693128 357040 693180
rect 450736 693128 450788 693180
rect 676320 693128 676372 693180
rect 208132 692516 208184 692568
rect 208960 692516 209012 692568
rect 226265 692383 226757 692698
rect 287712 692516 287764 692568
rect 608056 692040 608108 692092
rect 611460 692040 611512 692092
rect 320648 691428 320700 691480
rect 321108 691428 321160 691480
rect 676228 691162 676280 691214
rect 611184 690612 611236 690664
rect 612288 690612 612340 690664
rect 675860 690272 675912 690324
rect 676320 690272 676372 690324
rect 506304 689796 506356 689848
rect 675860 689796 675912 689848
rect 576960 689184 577012 689236
rect 590208 689184 590260 689236
rect 676044 688096 676096 688148
rect 676320 688096 676372 688148
rect 251740 687620 251792 687672
rect 279892 687620 279944 687672
rect 667488 687620 667540 687672
rect 675952 687620 676004 687672
rect 675676 687076 675728 687128
rect 676320 687076 676372 687128
rect 489744 687008 489796 687060
rect 496368 687008 496420 687060
rect 675768 687008 675820 687060
rect 676228 687008 676280 687060
rect 602352 684764 602404 684816
rect 611184 684764 611236 684816
rect 614496 684560 614548 684612
rect 615692 684560 615744 684612
rect 596832 684492 596884 684544
rect 603548 684492 603600 684544
rect 322028 684288 322080 684340
rect 360668 684288 360720 684340
rect 616704 684084 616756 684136
rect 617900 684084 617952 684136
rect 600144 683064 600196 683116
rect 603456 683064 603508 683116
rect 330768 682112 330820 682164
rect 359840 682112 359892 682164
rect 496368 682112 496420 682164
rect 506396 682112 506448 682164
rect 590208 681500 590260 681552
rect 600144 681500 600196 681552
rect 607964 681432 608016 681484
rect 612564 681432 612616 681484
rect 611276 681092 611328 681144
rect 612472 681092 612524 681144
rect 611460 681024 611512 681076
rect 614588 681024 614640 681076
rect 610080 680956 610132 681008
rect 613392 680956 613444 681008
rect 650928 680956 650980 681008
rect 654240 680956 654292 681008
rect 328560 678780 328612 678832
rect 362600 678780 362652 678832
rect 612564 677760 612616 677812
rect 614496 677760 614548 677812
rect 208132 677556 208184 677608
rect 209972 677556 210024 677608
rect 390200 676604 390252 676656
rect 390660 676604 390712 676656
rect 607872 676604 607924 676656
rect 608976 676604 609028 676656
rect 605664 676468 605716 676520
rect 606860 676468 606912 676520
rect 390200 676264 390252 676316
rect 390384 676264 390436 676316
rect 614588 676264 614640 676316
rect 616704 676264 616756 676316
rect 612472 676128 612524 676180
rect 614588 676128 614640 676180
rect 643200 675924 643252 675976
rect 650928 675924 650980 675976
rect 603548 674836 603600 674888
rect 610816 674836 610868 674888
rect 248152 674360 248204 674412
rect 287988 674360 288040 674412
rect 603456 673340 603508 673392
rect 606768 673340 606820 673392
rect 329664 673272 329716 673324
rect 360760 673272 360812 673324
rect 417524 671504 417576 671556
rect 536756 671504 536808 671556
rect 600144 671504 600196 671556
rect 612380 671504 612432 671556
rect 251648 671028 251700 671080
rect 286424 670960 286476 671012
rect 341072 670416 341124 670468
rect 352388 670416 352440 670468
rect 208132 669804 208184 669856
rect 209052 669804 209104 669856
rect 610816 669328 610868 669380
rect 617808 669328 617860 669380
rect 613392 668716 613444 668768
rect 616980 668716 617032 668768
rect 489284 668240 489336 668292
rect 516884 668240 516936 668292
rect 341506 667818 342830 667890
rect 252844 667764 252896 667816
rect 286608 667764 286660 667816
rect 286884 667764 286936 667816
rect 209328 667560 209380 667612
rect 210156 667560 210208 667612
rect 220076 667552 222120 667728
rect 615600 667628 615652 667680
rect 618912 667628 618964 667680
rect 335552 667560 335604 667612
rect 208132 667288 208184 667340
rect 210064 667288 210116 667340
rect 286884 667356 286936 667408
rect 337300 667356 337352 667408
rect 270232 667288 270284 667340
rect 290748 667288 290800 667340
rect 315496 667288 315548 667340
rect 316048 667288 316100 667340
rect 342544 667492 342596 667544
rect 341072 667433 341124 667476
rect 341072 667424 341081 667433
rect 341081 667424 341115 667433
rect 341115 667424 341124 667433
rect 338956 667356 339008 667408
rect 267840 667172 267892 667224
rect 270232 667152 270284 667204
rect 303168 667220 303220 667272
rect 337300 667220 337352 667272
rect 342544 667288 342596 667340
rect 362324 667288 362376 667340
rect 382932 667288 382984 667340
rect 360484 667220 360536 667272
rect 362416 667220 362468 667272
rect 308228 667084 308280 667136
rect 321936 667084 321988 667136
rect 340998 667088 342546 667170
rect 361128 667152 361180 667204
rect 361864 667152 361916 667204
rect 362692 667152 362744 667204
rect 363888 667152 363940 667204
rect 390108 667152 390160 667204
rect 569232 667152 569284 667204
rect 635472 667152 635524 667204
rect 643200 667152 643252 667204
rect 342912 667084 342964 667136
rect 236536 665954 242984 667020
rect 310160 667016 310212 667068
rect 361772 667084 361824 667136
rect 381092 667084 381144 667136
rect 318164 666948 318216 667000
rect 361220 667016 361272 667068
rect 297556 666880 297608 666932
rect 335644 666880 335696 666932
rect 342728 666948 342780 667000
rect 342912 666948 342964 667000
rect 375204 666948 375256 667000
rect 342820 666880 342872 666932
rect 344108 666880 344160 666932
rect 360484 666880 360536 666932
rect 361680 666880 361732 666932
rect 368856 666880 368908 666932
rect 369132 666880 369184 666932
rect 290656 666812 290708 666864
rect 390476 666812 390528 666864
rect 251556 666744 251608 666796
rect 289368 666744 289420 666796
rect 298752 666744 298804 666796
rect 373180 666744 373232 666796
rect 377136 666744 377188 666796
rect 379252 666744 379304 666796
rect 576500 666744 576552 666796
rect 250544 666676 250596 666728
rect 296176 666676 296228 666728
rect 377228 666676 377280 666728
rect 389372 666676 389424 666728
rect 612932 666676 612984 666728
rect 252752 666608 252804 666660
rect 290656 666608 290708 666660
rect 321016 666608 321068 666660
rect 365084 666608 365136 666660
rect 385324 666608 385376 666660
rect 615784 666608 615836 666660
rect 316876 666540 316928 666592
rect 637220 666540 637272 666592
rect 314116 666472 314168 666524
rect 598580 666472 598632 666524
rect 294796 666404 294848 666456
rect 370512 666404 370564 666456
rect 371156 666404 371208 666456
rect 288264 666336 288316 666388
rect 335552 666336 335604 666388
rect 335644 666336 335696 666388
rect 344108 666336 344160 666388
rect 611184 666336 611236 666388
rect 613392 666336 613444 666388
rect 290840 666268 290892 666320
rect 298752 666268 298804 666320
rect 288540 666200 288592 666252
rect 306480 666200 306532 666252
rect 252016 666132 252068 666184
rect 321292 666268 321344 666320
rect 363244 666268 363296 666320
rect 375204 666200 375256 666252
rect 605664 666200 605716 666252
rect 362508 666132 362560 666184
rect 615600 666132 615652 666184
rect 288448 666064 288500 666116
rect 594624 666064 594676 666116
rect 606860 666064 606912 666116
rect 613484 666064 613536 666116
rect 288172 665996 288224 666048
rect 598580 665996 598632 666048
rect 290748 665860 290800 665912
rect 321200 665860 321252 665912
rect 267840 665792 267892 665844
rect 320924 665792 320976 665844
rect 251464 665520 251516 665572
rect 290840 665520 290892 665572
rect 287988 665452 288040 665504
rect 390292 665452 390344 665504
rect 320740 665384 320792 665436
rect 389372 665384 389424 665436
rect 297832 665316 297884 665368
rect 298844 665316 298896 665368
rect 304916 665316 304968 665368
rect 305836 665316 305888 665368
rect 209052 665248 209104 665300
rect 320832 665316 320884 665368
rect 377136 665316 377188 665368
rect 248520 665180 248572 665232
rect 362876 665180 362928 665232
rect 378884 665180 378936 665232
rect 506304 665180 506356 665232
rect 210156 665112 210208 665164
rect 338956 665112 339008 665164
rect 362600 665112 362652 665164
rect 532340 665112 532392 665164
rect 288080 665044 288132 665096
rect 301604 665044 301656 665096
rect 304364 665044 304416 665096
rect 610264 665044 610316 665096
rect 292036 664976 292088 665028
rect 604652 664976 604704 665028
rect 289092 664908 289144 664960
rect 615968 664908 616020 664960
rect 287896 664840 287948 664892
rect 321476 664840 321528 664892
rect 319728 664772 319780 664824
rect 367108 664772 367160 664824
rect 617900 664772 617952 664824
rect 620016 664772 620068 664824
rect 608976 664500 609028 664552
rect 612196 664500 612248 664552
rect 569232 663956 569284 664008
rect 574752 663956 574804 664008
rect 675676 663956 675728 664008
rect 676044 663956 676096 664008
rect 306480 663888 306532 663940
rect 604560 663888 604612 663940
rect 300316 663820 300368 663872
rect 610080 663820 610132 663872
rect 615600 663820 615652 663872
rect 621304 663820 621356 663872
rect 676044 663820 676096 663872
rect 676688 663820 676740 663872
rect 675860 663616 675912 663668
rect 676228 663616 676280 663668
rect 675768 662936 675820 662988
rect 676596 662996 676648 663048
rect 614496 662868 614548 662920
rect 619096 662868 619148 662920
rect 252660 662732 252712 662784
rect 293324 662732 293376 662784
rect 362416 662732 362468 662784
rect 584228 662732 584280 662784
rect 604652 662732 604704 662784
rect 614496 662732 614548 662784
rect 675676 662256 675728 662308
rect 676136 662256 676188 662308
rect 671352 661916 671404 661968
rect 676320 661916 676372 661968
rect 615692 661848 615744 661900
rect 616796 661848 616848 661900
rect 604560 661712 604612 661764
rect 610172 661712 610224 661764
rect 612104 661304 612156 661356
rect 619372 661304 619424 661356
rect 251096 661100 251148 661152
rect 671352 661100 671404 661152
rect 359012 660488 359064 660540
rect 541172 660488 541224 660540
rect 675768 660284 675820 660336
rect 676320 660284 676372 660336
rect 606768 660080 606820 660132
rect 609160 660080 609212 660132
rect 613484 659468 613536 659520
rect 618268 659468 618320 659520
rect 402068 659400 402120 659452
rect 485972 659400 486024 659452
rect 614588 659400 614640 659452
rect 615692 659400 615744 659452
rect 616980 659060 617032 659112
rect 621488 659060 621540 659112
rect 610080 658924 610132 658976
rect 612288 658924 612340 658976
rect 615784 658448 615836 658500
rect 620108 658448 620160 658500
rect 615968 658380 616020 658432
rect 621028 658380 621080 658432
rect 307124 658312 307176 658364
rect 437488 658312 437540 658364
rect 468308 658312 468360 658364
rect 522496 658312 522548 658364
rect 574752 658312 574804 658364
rect 584688 658312 584740 658364
rect 675676 658108 675728 658160
rect 676044 658108 676096 658160
rect 637680 657768 637732 657820
rect 676228 657768 676280 657820
rect 675584 657360 675636 657412
rect 676228 657360 676280 657412
rect 506396 657224 506448 657276
rect 514032 657224 514084 657276
rect 610264 657224 610316 657276
rect 619004 657224 619056 657276
rect 282928 657156 282980 657208
rect 548900 657156 548952 657208
rect 594624 657156 594676 657208
rect 612196 657156 612248 657208
rect 675584 656680 675636 656732
rect 676320 656680 676372 656732
rect 605664 656204 605716 656256
rect 614404 656204 614456 656256
rect 675860 656204 675912 656256
rect 676320 656204 676372 656256
rect 248428 656136 248480 656188
rect 522588 656136 522640 656188
rect 584688 656136 584740 656188
rect 595728 656136 595780 656188
rect 247324 656068 247376 656120
rect 312644 656068 312696 656120
rect 315956 656068 316008 656120
rect 624432 656068 624484 656120
rect 675768 656000 675820 656052
rect 676136 656000 676188 656052
rect 675676 655592 675728 655644
rect 676320 655592 676372 655644
rect 610172 655048 610224 655100
rect 615508 655048 615560 655100
rect 620108 654912 620160 654964
rect 622132 654912 622184 654964
rect 621488 654708 621540 654760
rect 623144 654708 623196 654760
rect 213468 654504 213520 654556
rect 619280 654504 619332 654556
rect 675492 654232 675544 654284
rect 675952 654232 676004 654284
rect 675768 654164 675820 654216
rect 676044 654164 676096 654216
rect 258548 653960 258600 654012
rect 413108 653960 413160 654012
rect 501428 653960 501480 654012
rect 546692 653960 546744 654012
rect 618268 653960 618320 654012
rect 619464 653960 619516 654012
rect 250268 653892 250320 653944
rect 519184 653892 519236 653944
rect 553316 653892 553368 653944
rect 617900 653892 617952 653944
rect 620016 653620 620068 653672
rect 622592 653620 622644 653672
rect 251004 652940 251056 652992
rect 440708 652940 440760 652992
rect 250084 652872 250136 652924
rect 459476 652872 459528 652924
rect 517988 652872 518040 652924
rect 529212 652872 529264 652924
rect 609160 652872 609212 652924
rect 615600 652872 615652 652924
rect 368856 652804 368908 652856
rect 622960 652804 623012 652856
rect 361128 652736 361180 652788
rect 621672 652736 621724 652788
rect 616704 652328 616756 652380
rect 619188 652328 619240 652380
rect 676228 652396 676280 652448
rect 208132 652260 208184 652312
rect 209972 652260 210024 652312
rect 633264 652260 633316 652312
rect 208960 652056 209012 652108
rect 209144 652056 209196 652108
rect 619096 651920 619148 651972
rect 621120 651920 621172 651972
rect 250360 651784 250412 651836
rect 419916 651784 419968 651836
rect 615692 651784 615744 651836
rect 620844 651784 620896 651836
rect 251832 651716 251884 651768
rect 431876 651716 431928 651768
rect 595728 651716 595780 651768
rect 607872 651716 607924 651768
rect 249256 651648 249308 651700
rect 463984 651648 464036 651700
rect 561228 651648 561280 651700
rect 652676 651648 652728 651700
rect 668592 651648 668644 651700
rect 676044 651648 676096 651700
rect 675584 651580 675636 651632
rect 675860 651580 675912 651632
rect 675768 651376 675820 651428
rect 676228 651376 676280 651428
rect 615600 651036 615652 651088
rect 621396 651036 621448 651088
rect 619004 650832 619056 650884
rect 622224 650832 622276 650884
rect 495908 650764 495960 650816
rect 615600 650764 615652 650816
rect 619372 650764 619424 650816
rect 622408 650764 622460 650816
rect 390016 650696 390068 650748
rect 621856 650696 621908 650748
rect 389924 650628 389976 650680
rect 613300 650628 613352 650680
rect 613392 650628 613444 650680
rect 620936 650628 620988 650680
rect 370512 650560 370564 650612
rect 619740 650560 619792 650612
rect 615600 650492 615652 650544
rect 621948 650492 622000 650544
rect 613300 650424 613352 650476
rect 622868 650424 622920 650476
rect 612104 650356 612156 650408
rect 619004 650356 619056 650408
rect 676136 650362 676188 650414
rect 614496 650288 614548 650340
rect 622500 650288 622552 650340
rect 217056 650084 217108 650136
rect 551660 650084 551712 650136
rect 607872 649540 607924 649592
rect 619096 649540 619148 649592
rect 514032 649472 514084 649524
rect 617808 649472 617860 649524
rect 621212 649472 621264 649524
rect 623052 649404 623104 649456
rect 569232 649064 569284 649116
rect 676228 649064 676280 649116
rect 252292 648996 252344 649048
rect 675860 648996 675912 649048
rect 675492 648928 675544 648980
rect 675952 648928 676004 648980
rect 615508 648724 615560 648776
rect 619924 648724 619976 648776
rect 248060 648656 248112 648708
rect 304916 648656 304968 648708
rect 249440 648588 249492 648640
rect 316048 648588 316100 648640
rect 252568 648520 252620 648572
rect 319728 648520 319780 648572
rect 248244 648452 248296 648504
rect 321108 648452 321160 648504
rect 470148 648452 470200 648504
rect 569232 648452 569284 648504
rect 248336 648384 248388 648436
rect 324788 648384 324840 648436
rect 494804 648384 494856 648436
rect 618912 648384 618964 648436
rect 620660 648384 620712 648436
rect 628848 648384 628900 648436
rect 635472 648384 635524 648436
rect 622040 648316 622092 648368
rect 374284 647976 374336 648028
rect 624432 647976 624484 648028
rect 233616 647908 233668 647960
rect 623236 647908 623288 647960
rect 252476 647840 252528 647892
rect 671076 647840 671128 647892
rect 223680 647568 223732 647620
rect 622316 647568 622368 647620
rect 252108 647432 252160 647484
rect 320648 647432 320700 647484
rect 381092 647432 381144 647484
rect 388636 647432 388688 647484
rect 405380 647432 405432 647484
rect 426908 647432 426960 647484
rect 479716 647432 479768 647484
rect 625536 647432 625588 647484
rect 252200 647364 252252 647416
rect 321016 647364 321068 647416
rect 363888 647364 363940 647416
rect 412556 647364 412608 647416
rect 494068 647364 494120 647416
rect 645408 647364 645460 647416
rect 219264 647296 219316 647348
rect 288816 647296 288868 647348
rect 365268 647296 365320 647348
rect 383852 647296 383904 647348
rect 390384 647296 390436 647348
rect 619832 647296 619884 647348
rect 251372 647228 251424 647280
rect 544484 647228 544536 647280
rect 594716 647228 594768 647280
rect 642096 647228 642148 647280
rect 320556 647160 320608 647212
rect 503636 647160 503688 647212
rect 556444 647160 556496 647212
rect 620752 647160 620804 647212
rect 288816 647092 288868 647144
rect 407772 647092 407824 647144
rect 455796 647092 455848 647144
rect 640992 647092 641044 647144
rect 297556 647024 297608 647076
rect 308228 647024 308280 647076
rect 320464 647024 320516 647076
rect 393420 647024 393472 647076
rect 398204 647024 398256 647076
rect 671904 647024 671956 647076
rect 241344 646956 241396 647008
rect 619372 646956 619424 647008
rect 675676 646956 675728 647008
rect 676320 646956 676372 647008
rect 292772 646888 292824 646940
rect 323040 646888 323092 646940
rect 326260 646888 326312 646940
rect 635472 646888 635524 646940
rect 252384 646820 252436 646872
rect 255696 646820 255748 646872
rect 609068 646820 609120 646872
rect 631056 646820 631108 646872
rect 208408 646752 208460 646804
rect 268668 646752 268720 646804
rect 273636 646752 273688 646804
rect 297832 646752 297884 646804
rect 311908 646752 311960 646804
rect 638784 646752 638836 646804
rect 676228 646752 676280 646804
rect 676228 646480 676280 646532
rect 671076 646140 671128 646192
rect 676136 646140 676188 646192
rect 666752 645936 666804 645988
rect 676596 645936 676648 645988
rect 208316 644984 208368 645036
rect 210064 644984 210116 645036
rect 675768 644780 675820 644832
rect 676504 644780 676556 644832
rect 209420 643964 209472 644016
rect 233616 643964 233668 644016
rect 675584 643896 675636 643948
rect 676412 643896 676464 643948
rect 208040 640700 208092 640752
rect 208684 640700 208736 640752
rect 208592 640632 208644 640684
rect 209972 640632 210024 640684
rect 208224 640292 208276 640344
rect 208868 640292 208920 640344
rect 208224 639884 208276 639936
rect 208776 639884 208828 639936
rect 208040 638932 208092 638984
rect 208960 638932 209012 638984
rect 209328 638388 209380 638440
rect 223680 638388 223732 638440
rect 661968 637844 662020 637896
rect 668592 637844 668644 637896
rect 208684 636756 208736 636808
rect 208868 636756 208920 636808
rect 208776 636688 208828 636740
rect 209144 636688 209196 636740
rect 208408 636620 208460 636672
rect 208316 636552 208368 636604
rect 208684 636552 208736 636604
rect 208776 636552 208828 636604
rect 208040 636484 208092 636536
rect 208500 636484 208552 636536
rect 208960 635600 209012 635652
rect 623328 635124 623380 635176
rect 628848 635124 628900 635176
rect 208012 633070 208064 633122
rect 208230 633068 208282 633120
rect 230304 632880 230356 632932
rect 241344 632880 241396 632932
rect 621488 632404 621540 632456
rect 641912 632404 641964 632456
rect 208224 632200 208276 632252
rect 208316 632132 208368 632184
rect 208592 632132 208644 632184
rect 208500 632064 208552 632116
rect 208040 631996 208092 632048
rect 208592 631996 208644 632048
rect 208408 631928 208460 631980
rect 208776 631928 208828 631980
rect 208776 631792 208828 631844
rect 208960 631792 209012 631844
rect 675860 631724 675912 631776
rect 676320 631724 676372 631776
rect 676320 631588 676372 631640
rect 676688 631588 676740 631640
rect 676504 631452 676556 631504
rect 676688 631452 676740 631504
rect 208132 631044 208184 631096
rect 208960 631044 209012 631096
rect 208040 630772 208092 630824
rect 208684 630772 208736 630824
rect 641912 630704 641964 630756
rect 652032 630704 652084 630756
rect 208040 630024 208092 630076
rect 208316 630024 208368 630076
rect 209144 630024 209196 630076
rect 208040 629276 208092 629328
rect 208132 629072 208184 629124
rect 208776 629072 208828 629124
rect 208040 628800 208092 628852
rect 208592 628800 208644 628852
rect 675768 628732 675820 628784
rect 676320 628732 676372 628784
rect 675676 628664 675728 628716
rect 676228 628664 676280 628716
rect 208408 628528 208460 628580
rect 208684 628528 208736 628580
rect 676228 628528 676280 628580
rect 676688 628528 676740 628580
rect 645500 626284 645552 626336
rect 661968 626284 662020 626336
rect 228096 626012 228148 626064
rect 230304 626012 230356 626064
rect 208132 625740 208184 625792
rect 208132 625604 208184 625656
rect 619096 624516 619148 624568
rect 208408 624108 208460 624160
rect 208040 623904 208092 623956
rect 208224 623904 208276 623956
rect 208408 623836 208460 623888
rect 208316 623768 208368 623820
rect 208684 623768 208736 623820
rect 208040 623632 208092 623684
rect 208868 623632 208920 623684
rect 675584 622340 675636 622392
rect 676504 622340 676556 622392
rect 675308 621320 675360 621372
rect 675860 621320 675912 621372
rect 619096 621184 619148 621236
rect 675860 621184 675912 621236
rect 676228 621184 676280 621236
rect 675676 620980 675728 621032
rect 676320 620980 676372 621032
rect 675860 619484 675912 619536
rect 676320 619484 676372 619536
rect 619096 619212 619148 619264
rect 620016 619212 620068 619264
rect 619096 617376 619148 617428
rect 620016 617376 620068 617428
rect 620016 617172 620068 617224
rect 620660 617172 620712 617224
rect 643200 616968 643252 617020
rect 676320 616968 676372 617020
rect 676228 616424 676280 616476
rect 676320 616220 676372 616272
rect 675584 616084 675636 616136
rect 675492 615880 675544 615932
rect 625536 615812 625588 615864
rect 675768 615812 675820 615864
rect 676228 615812 676280 615864
rect 676320 615812 676372 615864
rect 675400 615744 675452 615796
rect 675492 615676 675544 615728
rect 676228 615676 676280 615728
rect 652032 615608 652084 615660
rect 654240 615608 654292 615660
rect 675860 614928 675912 614980
rect 676228 614928 676280 614980
rect 675308 614248 675360 614300
rect 676320 614248 676372 614300
rect 213744 614112 213796 614164
rect 228096 614112 228148 614164
rect 675400 613500 675452 613552
rect 675676 613500 675728 613552
rect 676228 613500 676280 613552
rect 619464 613160 619516 613212
rect 675584 613092 675636 613144
rect 676320 613092 676372 613144
rect 619096 613024 619148 613076
rect 619464 613024 619516 613076
rect 619096 612888 619148 612940
rect 675676 612208 675728 612260
rect 676228 612208 676280 612260
rect 675860 611936 675912 611988
rect 676320 611936 676372 611988
rect 207948 611800 208000 611852
rect 208684 611800 208736 611852
rect 208500 611732 208552 611784
rect 217056 611732 217108 611784
rect 208408 611638 208460 611690
rect 624432 611460 624484 611512
rect 676228 611460 676280 611512
rect 675492 611324 675544 611376
rect 676228 611324 676280 611376
rect 208049 611177 208101 611229
rect 208500 611204 208552 611256
rect 209512 610848 209564 610900
rect 213744 610848 213796 610900
rect 619096 610576 619148 610628
rect 619464 610576 619516 610628
rect 675308 609556 675360 609608
rect 208040 609148 208092 609200
rect 209788 609148 209840 609200
rect 675860 609080 675912 609132
rect 676320 609080 676372 609132
rect 675492 609012 675544 609064
rect 675952 609012 676004 609064
rect 675768 608944 675820 608996
rect 676320 608944 676372 608996
rect 208132 608536 208184 608588
rect 208776 608536 208828 608588
rect 208224 608196 208276 608248
rect 208500 608196 208552 608248
rect 675768 608128 675820 608180
rect 676228 608128 676280 608180
rect 675308 606564 675360 606616
rect 676320 606564 676372 606616
rect 675400 606156 675452 606208
rect 676320 606156 676372 606208
rect 233616 605884 233668 605936
rect 252384 605884 252436 605936
rect 625536 605884 625588 605936
rect 669696 605884 669748 605936
rect 675584 605816 675636 605868
rect 676320 605816 676372 605868
rect 643292 605340 643344 605392
rect 645500 605340 645552 605392
rect 675860 605340 675912 605392
rect 676504 605340 676556 605392
rect 675676 605272 675728 605324
rect 676596 605272 676648 605324
rect 675308 605204 675360 605256
rect 675860 605204 675912 605256
rect 675492 605136 675544 605188
rect 675952 605136 676004 605188
rect 675768 605068 675820 605120
rect 676228 605068 676280 605120
rect 208408 605000 208460 605052
rect 208408 604728 208460 604780
rect 208040 603232 208092 603284
rect 208592 603232 208644 603284
rect 654240 602008 654292 602060
rect 659760 602008 659812 602060
rect 208040 601396 208092 601448
rect 208316 601396 208368 601448
rect 209328 601396 209380 601448
rect 639888 601396 639940 601448
rect 643292 601396 643344 601448
rect 211536 599288 211588 599340
rect 244656 599288 244708 599340
rect 208132 598948 208184 599000
rect 208776 598948 208828 599000
rect 208040 598812 208092 598864
rect 208776 598812 208828 598864
rect 208040 597792 208092 597844
rect 208500 597792 208552 597844
rect 208684 597792 208736 597844
rect 208040 596772 208092 596824
rect 208776 596772 208828 596824
rect 208224 595072 208276 595124
rect 208592 595072 208644 595124
rect 209788 590448 209840 590500
rect 219356 590448 219408 590500
rect 659760 587660 659812 587712
rect 667488 587660 667540 587712
rect 637772 587184 637824 587236
rect 639888 587184 639940 587236
rect 208408 585484 208460 585536
rect 249072 585484 249124 585536
rect 208132 585416 208184 585468
rect 252384 585416 252436 585468
rect 208040 583852 208092 583904
rect 208776 583852 208828 583904
rect 209696 583852 209748 583904
rect 249164 583852 249216 583904
rect 676320 582220 676372 582272
rect 675768 582016 675820 582068
rect 635564 581880 635616 581932
rect 637772 581880 637824 581932
rect 208040 581744 208092 581796
rect 208500 581744 208552 581796
rect 675584 581404 675636 581456
rect 676504 581404 676556 581456
rect 624432 581336 624484 581388
rect 673376 581336 673428 581388
rect 208868 580792 208920 580844
rect 673376 580520 673428 580572
rect 676320 580588 676372 580640
rect 676320 580180 676372 580232
rect 675400 580044 675452 580096
rect 675860 580044 675912 580096
rect 676320 580044 676372 580096
rect 208316 578820 208368 578872
rect 208592 578820 208644 578872
rect 675676 578820 675728 578872
rect 676228 578820 676280 578872
rect 675584 578684 675636 578736
rect 676228 578684 676280 578736
rect 208040 578344 208092 578396
rect 208684 578344 208736 578396
rect 675400 578208 675452 578260
rect 676228 578208 676280 578260
rect 675492 578140 675544 578192
rect 675952 578140 676004 578192
rect 676136 578072 676188 578124
rect 676136 577936 676188 577988
rect 208224 577460 208276 577512
rect 208224 577120 208276 577172
rect 219356 576848 219408 576900
rect 221564 576848 221616 576900
rect 676320 576100 676372 576152
rect 676136 576032 676188 576084
rect 676136 575896 676188 575948
rect 675676 575760 675728 575812
rect 675952 575760 676004 575812
rect 675860 575692 675912 575744
rect 676228 575692 676280 575744
rect 675492 575556 675544 575608
rect 676228 575556 676280 575608
rect 676228 575420 676280 575472
rect 208040 575216 208092 575268
rect 208500 575216 208552 575268
rect 208316 575148 208368 575200
rect 208776 575148 208828 575200
rect 675860 575080 675912 575132
rect 676320 575080 676372 575132
rect 208040 574944 208092 574996
rect 208776 574944 208828 574996
rect 675308 574944 675360 574996
rect 675676 574944 675728 574996
rect 676044 574944 676096 574996
rect 676136 574944 676188 574996
rect 208684 574876 208736 574928
rect 208868 574876 208920 574928
rect 675768 574876 675820 574928
rect 675676 574808 675728 574860
rect 676044 574808 676096 574860
rect 676136 574808 676188 574860
rect 208224 574740 208276 574792
rect 208684 574740 208736 574792
rect 675952 574740 676004 574792
rect 676320 574740 676372 574792
rect 208316 574536 208368 574588
rect 208500 574536 208552 574588
rect 675308 574128 675360 574180
rect 676320 574128 676372 574180
rect 208040 573584 208092 573636
rect 208868 573584 208920 573636
rect 675492 573584 675544 573636
rect 676320 573584 676372 573636
rect 674112 572292 674164 572344
rect 676228 572292 676280 572344
rect 208224 571748 208276 571800
rect 208500 571748 208552 571800
rect 208132 571612 208184 571664
rect 208500 571612 208552 571664
rect 675860 571476 675912 571528
rect 676228 571476 676280 571528
rect 675584 571136 675636 571188
rect 676320 571136 676372 571188
rect 675584 571000 675636 571052
rect 675952 571000 676004 571052
rect 208224 570728 208276 570780
rect 208684 570728 208736 570780
rect 667488 570592 667540 570644
rect 676228 570592 676280 570644
rect 208040 569164 208092 569216
rect 208684 569164 208736 569216
rect 208868 569164 208920 569216
rect 208132 569096 208184 569148
rect 208592 569096 208644 569148
rect 208040 568756 208092 568808
rect 208776 568756 208828 568808
rect 675400 568756 675452 568808
rect 675952 568756 676004 568808
rect 619280 568416 619332 568468
rect 629768 568416 629820 568468
rect 623420 568348 623472 568400
rect 635564 568348 635616 568400
rect 675400 567804 675452 567856
rect 675676 567804 675728 567856
rect 208132 567736 208184 567788
rect 221472 567736 221524 567788
rect 675676 567668 675728 567720
rect 675952 567668 676004 567720
rect 208132 566648 208184 566700
rect 209052 566648 209104 566700
rect 629768 566648 629820 566700
rect 645500 566648 645552 566700
rect 675676 565696 675728 565748
rect 676228 565696 676280 565748
rect 221564 565560 221616 565612
rect 225888 565560 225940 565612
rect 675492 565356 675544 565408
rect 676320 565356 676372 565408
rect 675400 565016 675452 565068
rect 676320 565016 676372 565068
rect 675768 564540 675820 564592
rect 676596 564540 676648 564592
rect 675308 563792 675360 563844
rect 676688 563792 676740 563844
rect 675584 563384 675636 563436
rect 676228 563384 676280 563436
rect 645500 561888 645552 561940
rect 649824 561888 649876 561940
rect 676504 558964 676556 559016
rect 676688 558964 676740 559016
rect 664176 558896 664228 558948
rect 670800 558896 670852 558948
rect 676412 558828 676464 558880
rect 676688 558828 676740 558880
rect 208500 557808 208552 557860
rect 251188 557808 251240 557860
rect 208132 557672 208184 557724
rect 208500 557672 208552 557724
rect 208040 556924 208092 556976
rect 208960 556924 209012 556976
rect 225888 556856 225940 556908
rect 234720 556856 234772 556908
rect 208040 556720 208092 556772
rect 208040 556516 208092 556568
rect 208684 556516 208736 556568
rect 208408 556244 208460 556296
rect 244656 556244 244708 556296
rect 619096 554680 619148 554732
rect 619280 554680 619332 554732
rect 208316 554408 208368 554460
rect 208776 554408 208828 554460
rect 208224 554340 208276 554392
rect 208868 554340 208920 554392
rect 208224 553388 208276 553440
rect 208684 553388 208736 553440
rect 208132 552300 208184 552352
rect 208684 552300 208736 552352
rect 208040 550866 208092 550918
rect 208500 550866 208552 550918
rect 208040 549920 208092 549972
rect 208224 549920 208276 549972
rect 208040 549444 208092 549496
rect 208684 549444 208736 549496
rect 234720 548968 234772 549020
rect 243552 548968 243604 549020
rect 208040 548016 208092 548068
rect 208408 548016 208460 548068
rect 208776 548016 208828 548068
rect 208040 547676 208092 547728
rect 208868 547676 208920 547728
rect 620016 547404 620068 547456
rect 641084 547404 641136 547456
rect 208040 546588 208092 546640
rect 208224 546588 208276 546640
rect 209420 546588 209472 546640
rect 208224 546384 208276 546436
rect 208868 546384 208920 546436
rect 208040 546180 208092 546232
rect 208776 546180 208828 546232
rect 649824 545704 649876 545756
rect 651296 545704 651348 545756
rect 619096 545228 619148 545280
rect 619372 545228 619424 545280
rect 208040 544072 208092 544124
rect 208960 544072 209012 544124
rect 208408 543936 208460 543988
rect 208592 543936 208644 543988
rect 208040 543868 208092 543920
rect 208684 543868 208736 543920
rect 675860 543664 675912 543716
rect 676228 543664 676280 543716
rect 675768 543596 675820 543648
rect 676320 543596 676372 543648
rect 619096 543528 619148 543580
rect 619280 543528 619332 543580
rect 651296 543120 651348 543172
rect 661968 543120 662020 543172
rect 208040 541964 208092 542016
rect 208776 541964 208828 542016
rect 641084 541896 641136 541948
rect 644304 541896 644356 541948
rect 208316 541624 208368 541676
rect 208224 541556 208276 541608
rect 675400 540536 675452 540588
rect 676688 540536 676740 540588
rect 675584 540468 675636 540520
rect 676504 540468 676556 540520
rect 675676 540400 675728 540452
rect 676596 540400 676648 540452
rect 208040 540196 208092 540248
rect 208684 540196 208736 540248
rect 208500 540128 208552 540180
rect 214848 540128 214900 540180
rect 671904 539788 671956 539840
rect 676136 539652 676188 539704
rect 676320 539652 676372 539704
rect 676136 539448 676188 539500
rect 675492 539176 675544 539228
rect 676228 539176 676280 539228
rect 644304 538700 644356 538752
rect 648720 538700 648772 538752
rect 675584 537680 675636 537732
rect 676320 537680 676372 537732
rect 676228 537000 676280 537052
rect 676320 537000 676372 537052
rect 675676 536796 675728 536848
rect 676320 536796 676372 536848
rect 675676 535980 675728 536032
rect 676136 535980 676188 536032
rect 620016 535232 620068 535284
rect 676136 535232 676188 535284
rect 675400 535164 675452 535216
rect 675860 535164 675912 535216
rect 676044 535028 676096 535080
rect 676044 534892 676096 534944
rect 675676 534552 675728 534604
rect 676228 534552 676280 534604
rect 676044 534212 676096 534264
rect 676044 534076 676096 534128
rect 675400 533872 675452 533924
rect 675952 533872 676004 533924
rect 676320 533872 676372 533924
rect 675584 533192 675636 533244
rect 676136 533192 676188 533244
rect 675492 532580 675544 532632
rect 676320 532580 676372 532632
rect 620108 532512 620160 532564
rect 622500 532512 622552 532564
rect 675768 532376 675820 532428
rect 676136 532376 676188 532428
rect 631056 530812 631108 530864
rect 676136 530812 676188 530864
rect 675676 530200 675728 530252
rect 676320 530200 676372 530252
rect 635472 529724 635524 529776
rect 676136 529724 676188 529776
rect 675952 529588 676004 529640
rect 676136 529588 676188 529640
rect 208040 529180 208092 529232
rect 208592 529180 208644 529232
rect 208132 529112 208184 529164
rect 208224 529112 208276 529164
rect 208132 528908 208184 528960
rect 208224 528908 208276 528960
rect 675676 527752 675728 527804
rect 676228 527752 676280 527804
rect 208040 527004 208092 527056
rect 208224 527004 208276 527056
rect 208592 527004 208644 527056
rect 208224 526868 208276 526920
rect 208224 525984 208276 526036
rect 659760 525100 659812 525152
rect 664176 525100 664228 525152
rect 675584 524624 675636 524676
rect 676320 524624 676372 524676
rect 675860 523944 675912 523996
rect 676228 523944 676280 523996
rect 208023 523467 208075 523519
rect 208309 523461 208361 523513
rect 208040 522816 208092 522868
rect 208684 522816 208736 522868
rect 208037 522406 208089 522458
rect 209188 522411 209240 522463
rect 208408 522312 208460 522364
rect 209512 522312 209564 522364
rect 648720 521360 648772 521412
rect 658656 521360 658708 521412
rect 208224 521292 208276 521344
rect 208592 521292 208644 521344
rect 208500 520816 208552 520868
rect 208776 520816 208828 520868
rect 208224 520748 208276 520800
rect 208592 520748 208644 520800
rect 208132 520680 208184 520732
rect 208500 520680 208552 520732
rect 676320 520612 676372 520664
rect 676412 520408 676464 520460
rect 675768 520272 675820 520324
rect 676136 520272 676188 520324
rect 208040 519660 208092 519712
rect 208592 519660 208644 519712
rect 208040 519524 208092 519576
rect 208316 519524 208368 519576
rect 208776 519524 208828 519576
rect 208132 518164 208184 518216
rect 208316 517960 208368 518012
rect 208224 517892 208276 517944
rect 208592 517892 208644 517944
rect 668592 517008 668644 517060
rect 674204 517008 674256 517060
rect 208040 516804 208092 516856
rect 208776 516804 208828 516856
rect 208132 516124 208184 516176
rect 208132 515988 208184 516040
rect 208132 514628 208184 514680
rect 208500 514628 208552 514680
rect 208040 514356 208092 514408
rect 208500 514356 208552 514408
rect 214848 514288 214900 514340
rect 250820 514288 250872 514340
rect 208036 514169 208088 514221
rect 244854 514170 244906 514222
rect 650928 512588 650980 512640
rect 659760 512588 659812 512640
rect 658656 509256 658708 509308
rect 675768 509256 675820 509308
rect 619464 506196 619516 506248
rect 623328 506196 623380 506248
rect 243552 505380 243604 505432
rect 246864 505380 246916 505432
rect 675860 504836 675912 504888
rect 676228 504836 676280 504888
rect 208500 503748 208552 503800
rect 208776 503748 208828 503800
rect 675492 502660 675544 502712
rect 676136 502660 676188 502712
rect 676228 502660 676280 502712
rect 676688 502660 676740 502712
rect 666384 502320 666436 502372
rect 668592 502320 668644 502372
rect 676136 502116 676188 502168
rect 676504 502116 676556 502168
rect 675768 502048 675820 502100
rect 676320 502048 676372 502100
rect 208176 501708 208228 501760
rect 208520 501708 208572 501760
rect 208010 501640 208062 501692
rect 208776 501640 208828 501692
rect 675768 501572 675820 501624
rect 676596 501572 676648 501624
rect 675676 500416 675728 500468
rect 676136 500416 676188 500468
rect 676136 499940 676188 499992
rect 676412 499940 676464 499992
rect 208224 499736 208276 499788
rect 208776 499736 208828 499788
rect 208132 499668 208184 499720
rect 208500 499668 208552 499720
rect 662060 499124 662112 499176
rect 666384 499124 666436 499176
rect 676320 498920 676372 498972
rect 675584 498852 675636 498904
rect 676228 498852 676280 498904
rect 676320 498784 676372 498836
rect 675768 498716 675820 498768
rect 676228 498716 676280 498768
rect 208132 498512 208184 498564
rect 208408 498512 208460 498564
rect 208408 498376 208460 498428
rect 208684 498376 208736 498428
rect 676320 498376 676372 498428
rect 676136 498240 676188 498292
rect 676320 498240 676372 498292
rect 661968 497084 662020 497136
rect 669696 497084 669748 497136
rect 675768 496880 675820 496932
rect 676320 496880 676372 496932
rect 208316 496268 208368 496320
rect 208592 496268 208644 496320
rect 675676 496200 675728 496252
rect 676136 496200 676188 496252
rect 676320 496200 676372 496252
rect 208040 495928 208092 495980
rect 208500 495928 208552 495980
rect 675400 495452 675452 495504
rect 675860 495452 675912 495504
rect 675860 495316 675912 495368
rect 676044 495316 676096 495368
rect 673376 495112 673428 495164
rect 676136 495112 676188 495164
rect 645408 494432 645460 494484
rect 673376 494432 673428 494484
rect 675308 494160 675360 494212
rect 675676 494160 675728 494212
rect 676228 494160 676280 494212
rect 675676 493752 675728 493804
rect 676320 493752 676372 493804
rect 669696 493276 669748 493328
rect 675676 493276 675728 493328
rect 208132 493208 208184 493260
rect 208684 493208 208736 493260
rect 675400 493072 675452 493124
rect 676320 493072 676372 493124
rect 208040 492596 208092 492648
rect 208684 492596 208736 492648
rect 660864 492188 660916 492240
rect 675768 492188 675820 492240
rect 676136 492188 676188 492240
rect 675584 491780 675636 491832
rect 676320 491780 676372 491832
rect 645408 491576 645460 491628
rect 650928 491576 650980 491628
rect 675492 491576 675544 491628
rect 676136 491576 676188 491628
rect 208040 490556 208092 490608
rect 675860 490420 675912 490472
rect 676320 490420 676372 490472
rect 208132 490352 208184 490404
rect 208500 490352 208552 490404
rect 208224 490284 208276 490336
rect 208776 490284 208828 490336
rect 208040 489400 208092 489452
rect 675768 489400 675820 489452
rect 676320 489400 676372 489452
rect 208040 488652 208092 488704
rect 208684 488652 208736 488704
rect 208040 487156 208092 487208
rect 208960 487156 209012 487208
rect 675860 486952 675912 487004
rect 676044 486952 676096 487004
rect 675676 486068 675728 486120
rect 676320 486068 676372 486120
rect 208684 485796 208736 485848
rect 208408 485728 208460 485780
rect 675860 483960 675912 484012
rect 676320 483960 676372 484012
rect 675492 483552 675544 483604
rect 676228 483552 676280 483604
rect 675768 483416 675820 483468
rect 676228 483416 676280 483468
rect 659760 483348 659812 483400
rect 675860 483348 675912 483400
rect 641084 483212 641136 483264
rect 645408 483212 645460 483264
rect 208224 481716 208276 481768
rect 676044 481648 676096 481700
rect 676576 481648 676628 481700
rect 675492 481512 675544 481564
rect 676044 481512 676096 481564
rect 208224 481444 208276 481496
rect 221472 478928 221524 478980
rect 250820 478928 250872 478980
rect 657552 475528 657604 475580
rect 661968 475528 662020 475580
rect 671904 475392 671956 475444
rect 676228 475392 676280 475444
rect 211168 475052 211220 475104
rect 219264 475052 219316 475104
rect 207948 474616 208000 474668
rect 208408 474616 208460 474668
rect 208040 474236 208092 474288
rect 208868 474236 208920 474288
rect 638876 473828 638928 473880
rect 641084 473828 641136 473880
rect 208040 470986 208092 471038
rect 209052 470972 209104 471024
rect 208224 470904 208276 470956
rect 208776 470904 208828 470956
rect 208316 470836 208368 470888
rect 208224 470632 208276 470684
rect 208132 470360 208184 470412
rect 208500 470360 208552 470412
rect 208040 467640 208092 467692
rect 208868 467640 208920 467692
rect 208408 466348 208460 466400
rect 208040 466280 208092 466332
rect 208500 466144 208552 466196
rect 208040 466076 208092 466128
rect 208592 466076 208644 466128
rect 208040 465464 208092 465516
rect 208776 465464 208828 465516
rect 208040 464784 208092 464836
rect 209052 464784 209104 464836
rect 620200 464036 620252 464088
rect 621304 464036 621356 464088
rect 656448 462880 656500 462932
rect 671904 462880 671956 462932
rect 208040 462812 208092 462864
rect 208868 462812 208920 462864
rect 208224 461792 208276 461844
rect 208592 461792 208644 461844
rect 208132 459140 208184 459192
rect 208500 459140 208552 459192
rect 208316 459072 208368 459124
rect 208500 459004 208552 459056
rect 208776 459004 208828 459056
rect 644488 458460 644540 458512
rect 656448 458460 656500 458512
rect 208040 457440 208092 457492
rect 208408 457440 208460 457492
rect 623328 454652 623380 454704
rect 644488 454652 644540 454704
rect 208132 447512 208184 447564
rect 208868 447512 208920 447564
rect 207948 447202 208000 447254
rect 208408 447202 208460 447254
rect 208224 447104 208276 447156
rect 208224 446832 208276 446884
rect 208040 446628 208092 446680
rect 208684 446628 208736 446680
rect 627836 446288 627888 446340
rect 638876 446288 638928 446340
rect 208040 444384 208092 444436
rect 208776 444384 208828 444436
rect 645408 444112 645460 444164
rect 657552 444112 657604 444164
rect 208776 443568 208828 443620
rect 208132 441596 208184 441648
rect 208500 441596 208552 441648
rect 208224 441528 208276 441580
rect 208592 441528 208644 441580
rect 208500 441392 208552 441444
rect 208592 441392 208644 441444
rect 208040 438196 208092 438248
rect 208500 438196 208552 438248
rect 208868 438196 208920 438248
rect 208040 437380 208092 437432
rect 208684 437380 208736 437432
rect 208960 437380 209012 437432
rect 208132 437312 208184 437364
rect 208408 437312 208460 437364
rect 625628 437108 625680 437160
rect 627836 437108 627888 437160
rect 641084 436836 641136 436888
rect 645408 436836 645460 436888
rect 208040 433640 208092 433692
rect 208776 433640 208828 433692
rect 209512 433640 209564 433692
rect 208960 432008 209012 432060
rect 210156 432008 210208 432060
rect 208132 431736 208184 431788
rect 208132 431464 208184 431516
rect 208132 427384 208184 427436
rect 209972 427384 210024 427436
rect 635472 426636 635524 426688
rect 641084 426636 641136 426688
rect 620108 425276 620160 425328
rect 625628 425276 625680 425328
rect 620200 425004 620252 425056
rect 621120 425004 621172 425056
rect 620292 423168 620344 423220
rect 635472 423168 635524 423220
rect 208316 422080 208368 422132
rect 226992 422080 227044 422132
rect 208040 422012 208092 422064
rect 228096 422012 228148 422064
rect 232236 421536 232288 421588
rect 250820 421536 250872 421588
rect 619004 414600 619056 414652
rect 619188 414600 619240 414652
rect 208132 411200 208184 411252
rect 209972 411200 210024 411252
rect 208040 410520 208092 410572
rect 209512 410520 209564 410572
rect 210064 410520 210116 410572
rect 208040 409670 208092 409722
rect 208040 408276 208092 408328
rect 208316 408276 208368 408328
rect 208040 407528 208092 407580
rect 210248 407528 210300 407580
rect 208132 407188 208184 407240
rect 210156 407188 210208 407240
rect 208040 405488 208092 405540
rect 208868 405488 208920 405540
rect 248152 396580 248204 396632
rect 252200 396580 252252 396632
rect 208132 390664 208184 390716
rect 210248 390664 210300 390716
rect 208316 390392 208368 390444
rect 210064 390392 210116 390444
rect 208040 389780 208092 389832
rect 208868 389780 208920 389832
rect 208011 387271 208063 387323
rect 208221 387275 208273 387327
rect 208040 386312 208092 386364
rect 208408 386312 208460 386364
rect 228096 386244 228148 386296
rect 250084 386244 250136 386296
rect 227636 385428 227688 385480
rect 228096 385428 228148 385480
rect 208132 385088 208184 385140
rect 208592 385088 208644 385140
rect 208040 383456 208092 383508
rect 208408 383456 208460 383508
rect 208040 383048 208092 383100
rect 208592 383048 208644 383100
rect 208408 380600 208460 380652
rect 210432 380600 210484 380652
rect 208032 379854 208084 379906
rect 208236 379856 208288 379908
rect 209420 372032 209472 372084
rect 210524 372032 210576 372084
rect 210524 367680 210576 367732
rect 217056 367680 217108 367732
rect 217056 357616 217108 357668
rect 221472 357616 221524 357668
rect 221472 329260 221524 329312
rect 222392 329260 222444 329312
rect 222392 320488 222444 320540
rect 233708 320488 233760 320540
rect 209328 316068 209380 316120
rect 217056 316068 217108 316120
rect 217056 302808 217108 302860
rect 229200 302808 229252 302860
rect 233708 297436 233760 297488
rect 238032 297436 238084 297488
rect 229200 293968 229252 294020
rect 233708 293968 233760 294020
rect 238032 290976 238084 291028
rect 240240 290976 240292 291028
rect 233708 287508 233760 287560
rect 244656 287508 244708 287560
rect 621120 285400 621172 285452
rect 623052 285400 623104 285452
rect 229752 284516 229804 284568
rect 232328 284516 232380 284568
rect 232328 284040 232380 284092
rect 250176 284040 250228 284092
rect 634944 280890 636264 281126
rect 639520 280751 639572 280760
rect 639520 280717 639529 280751
rect 639529 280717 639563 280751
rect 639563 280717 639572 280751
rect 639520 280708 639572 280717
rect 248428 280504 248480 280556
rect 257444 280504 257496 280556
rect 617164 280504 617216 280556
rect 625076 280504 625128 280556
rect 250636 280436 250688 280488
rect 262228 280436 262280 280488
rect 607596 280436 607648 280488
rect 619832 280436 619884 280488
rect 251188 280368 251240 280420
rect 362876 280368 362928 280420
rect 588276 280368 588328 280420
rect 622040 280368 622092 280420
rect 250544 280300 250596 280352
rect 420284 280300 420336 280352
rect 435004 280300 435056 280352
rect 621120 280300 621172 280352
rect 642326 280712 643110 280916
rect 251372 280232 251424 280284
rect 271888 280232 271940 280284
rect 360576 280232 360628 280284
rect 549912 280232 549964 280284
rect 573924 280232 573976 280284
rect 621948 280232 622000 280284
rect 252108 280164 252160 280216
rect 675952 280164 676004 280216
rect 252384 280096 252436 280148
rect 643200 280096 643252 280148
rect 250728 280028 250780 280080
rect 310344 280028 310396 280080
rect 612472 280028 612524 280080
rect 633264 280028 633316 280080
rect 249164 279960 249216 280012
rect 511640 279960 511692 280012
rect 554880 279960 554932 280012
rect 646512 279960 646564 280012
rect 367936 279892 367988 279944
rect 624432 279892 624484 279944
rect 211536 279824 211588 279876
rect 463800 279824 463852 279876
rect 487720 279824 487772 279876
rect 637680 279824 637732 279876
rect 232512 279756 232564 279808
rect 473368 279756 473420 279808
rect 497288 279756 497340 279808
rect 625536 279756 625588 279808
rect 252752 279688 252804 279740
rect 430312 279688 430364 279740
rect 454232 279688 454284 279740
rect 675216 279688 675268 279740
rect 249440 279620 249492 279672
rect 415776 279620 415828 279672
rect 251556 279552 251608 279604
rect 387072 279552 387124 279604
rect 251464 279484 251516 279536
rect 286424 279484 286476 279536
rect 344016 279484 344068 279536
rect 620016 279484 620068 279536
rect 248244 279416 248296 279468
rect 377504 279416 377556 279468
rect 232328 279076 232380 279128
rect 248152 279076 248204 279128
rect 248520 279076 248572 279128
rect 251924 279076 251976 279128
rect 676136 279076 676188 279128
rect 252200 279008 252252 279060
rect 676300 279008 676352 279060
rect 249072 278940 249124 278992
rect 564448 278940 564500 278992
rect 569232 278940 569284 278992
rect 619648 278940 619700 278992
rect 535744 278872 535796 278924
rect 621672 278872 621724 278924
rect 251740 278804 251792 278856
rect 516608 278804 516660 278856
rect 526176 278804 526228 278856
rect 619740 278804 619792 278856
rect 250452 278736 250504 278788
rect 502492 278736 502544 278788
rect 506856 278736 506908 278788
rect 619556 278736 619608 278788
rect 249532 278668 249584 278720
rect 492504 278668 492556 278720
rect 578800 278668 578852 278720
rect 622960 278668 623012 278720
rect 250912 278600 250964 278652
rect 382288 278600 382340 278652
rect 401424 278600 401476 278652
rect 621764 278600 621816 278652
rect 248336 278532 248388 278584
rect 410992 278532 411044 278584
rect 248152 278464 248204 278516
rect 360576 278464 360628 278516
rect 249624 278396 249676 278448
rect 315128 278396 315180 278448
rect 252844 278328 252896 278380
rect 300776 278328 300828 278380
rect 251648 278260 251700 278312
rect 540528 278260 540580 278312
rect 244853 278019 244905 278071
rect 449468 278020 449520 278072
rect 281645 277909 281697 277962
rect 673318 277908 673370 277960
rect 611184 276288 611236 276340
rect 619096 276288 619148 276340
rect 609712 274112 609764 274164
rect 620752 274112 620804 274164
rect 229844 266360 229896 266412
rect 576960 266360 577012 266412
rect 339048 265272 339100 265324
rect 611736 265272 611788 265324
rect 324696 264184 324748 264236
rect 604560 264184 604612 264236
rect 610264 263164 610316 263216
rect 611184 263164 611236 263216
rect 208040 263028 208092 263080
rect 384312 263028 384364 263080
rect 391856 263028 391908 263080
rect 601984 263028 602036 263080
rect 577604 262076 577656 262128
rect 622868 262076 622920 262128
rect 565920 262008 565972 262060
rect 621856 262008 621908 262060
rect 252016 261940 252068 261992
rect 640256 261940 640308 261992
rect 583584 260852 583636 260904
rect 638876 260852 638928 260904
rect 587356 260240 587408 260292
rect 620016 260240 620068 260292
rect 652584 260240 652636 260292
rect 590484 260104 590536 260156
rect 592692 260104 592744 260156
rect 610816 260104 610868 260156
rect 625260 260104 625312 260156
rect 643384 260104 643436 260156
rect 397560 259900 397612 259952
rect 423872 259900 423924 259952
rect 424608 259900 424660 259952
rect 456992 259900 457044 259952
rect 489560 259900 489612 259952
rect 522220 259968 522272 260020
rect 554788 259968 554840 260020
rect 587356 260036 587408 260088
rect 610448 260036 610500 260088
rect 618636 260036 618688 260088
rect 610264 259960 610316 260012
rect 545588 259900 545640 259952
rect 548440 259900 548492 259952
rect 395076 259832 395128 259884
rect 397284 259832 397336 259884
rect 415408 259832 415460 259884
rect 423688 259832 423740 259884
rect 382826 259696 382878 259748
rect 384981 259716 385033 259768
rect 388377 259696 388429 259748
rect 389299 259716 389351 259768
rect 414856 259764 414908 259816
rect 418068 259764 418120 259816
rect 397836 259708 397888 259760
rect 210432 259628 210484 259680
rect 391985 259628 392037 259680
rect 247416 259560 247468 259612
rect 384496 259512 384548 259564
rect 389188 259512 389240 259564
rect 391396 259512 391448 259564
rect 395797 259504 395849 259556
rect 397560 259504 397612 259556
rect 397676 259504 397728 259556
rect 397836 259504 397888 259556
rect 418448 259552 418500 259604
rect 421894 259746 421946 259798
rect 426448 259764 426500 259816
rect 427736 259764 427788 259816
rect 429852 259764 429904 259816
rect 454416 259784 454468 259836
rect 457176 259764 457228 259816
rect 462696 259764 462748 259816
rect 480268 259764 480320 259816
rect 483472 259768 483524 259820
rect 430276 259696 430328 259748
rect 447838 259696 447890 259748
rect 449981 259696 450033 259748
rect 453377 259696 453429 259748
rect 457650 259696 457702 259748
rect 458028 259696 458080 259748
rect 458878 259696 458930 259748
rect 460086 259696 460138 259748
rect 462267 259696 462319 259748
rect 480426 259696 480478 259748
rect 482581 259696 482633 259748
rect 494712 259764 494764 259816
rect 513020 259832 513072 259884
rect 522404 259832 522456 259884
rect 522864 259832 522916 259884
rect 523232 259832 523284 259884
rect 524060 259832 524112 259884
rect 525256 259832 525308 259884
rect 527464 259832 527516 259884
rect 512836 259764 512888 259816
rect 423688 259628 423740 259680
rect 423856 259628 423908 259680
rect 428397 259628 428449 259680
rect 456256 259628 456308 259680
rect 460797 259628 460849 259680
rect 486899 259696 486951 259748
rect 495276 259696 495328 259748
rect 513020 259696 513072 259748
rect 515182 259696 515234 259748
rect 516148 259716 516200 259768
rect 518540 259764 518592 259816
rect 545312 259832 545364 259884
rect 558652 259900 558704 259952
rect 586620 259900 586672 259952
rect 611736 259968 611788 260020
rect 617256 259968 617308 260020
rect 638784 260036 638836 260088
rect 645592 260036 645644 260088
rect 643016 259968 643068 260020
rect 653228 260036 653280 260088
rect 545588 259764 545640 259816
rect 551200 259832 551252 259884
rect 553500 259764 553552 259816
rect 519506 259696 519558 259748
rect 527878 259696 527930 259748
rect 545036 259696 545088 259748
rect 547781 259696 547833 259748
rect 552099 259696 552151 259748
rect 555432 259832 555484 259884
rect 578064 259832 578116 259884
rect 580824 259832 580876 259884
rect 488856 259628 488908 259680
rect 493397 259628 493449 259680
rect 521456 259628 521508 259680
rect 525992 259628 526044 259680
rect 558652 259764 558704 259816
rect 577788 259764 577840 259816
rect 601984 259832 602036 259884
rect 613024 259900 613076 259952
rect 620660 259900 620712 259952
rect 642096 259900 642148 259952
rect 556677 259696 556729 259748
rect 565920 259696 565972 259748
rect 576960 259696 577012 259748
rect 584688 259746 584740 259798
rect 586068 259764 586120 259816
rect 604560 259764 604612 259816
rect 616336 259832 616388 259884
rect 640992 259832 641044 259884
rect 649916 259900 649968 259952
rect 586620 259696 586672 259748
rect 591197 259696 591249 259748
rect 621856 259764 621908 259816
rect 638876 259764 638928 259816
rect 648996 259832 649048 259884
rect 651296 259832 651348 259884
rect 657828 259832 657880 259884
rect 554052 259628 554104 259680
rect 554998 259628 555050 259680
rect 555828 259628 555880 259680
rect 557886 259628 557938 259680
rect 560067 259628 560119 259680
rect 560476 259628 560528 259680
rect 578226 259628 578278 259680
rect 580381 259628 580433 259680
rect 583777 259628 583829 259680
rect 593076 259628 593128 259680
rect 610632 259628 610684 259680
rect 619256 259696 619308 259748
rect 623788 259696 623840 259748
rect 421756 259512 421808 259564
rect 431204 259492 431256 259544
rect 446320 259492 446372 259544
rect 451012 259513 451064 259565
rect 454140 259512 454192 259564
rect 483463 259512 483515 259564
rect 516148 259512 516200 259564
rect 548440 259512 548492 259564
rect 580608 259522 580660 259574
rect 584504 259522 584556 259574
rect 643384 259628 643436 259680
rect 646462 259688 646514 259740
rect 651856 259696 651908 259748
rect 654477 259696 654529 259748
rect 659760 259696 659812 259748
rect 610908 259512 610960 259564
rect 615600 259512 615652 259564
rect 625674 259560 625726 259612
rect 627744 259560 627796 259612
rect 632528 259560 632580 259612
rect 649640 259628 649692 259680
rect 652798 259628 652850 259680
rect 653628 259628 653680 259680
rect 655686 259628 655738 259680
rect 657722 259628 657774 259680
rect 657828 259628 657880 259680
rect 676044 259628 676096 259680
rect 646462 259540 646514 259592
rect 658276 259560 658328 259612
rect 414856 259288 414908 259340
<< obsm1 >>
rect 519318 259446 519378 259448
<< metal2 >>
rect 250912 729016 250964 729022
rect 250912 728958 250964 728964
rect 246312 725684 246364 725690
rect 246312 725626 246364 725632
rect 208130 715785 208186 715794
rect 208130 715720 208186 715729
rect 208144 714858 208172 715720
rect 208222 715615 208278 715624
rect 208222 715550 208278 715559
rect 208130 714849 208186 714858
rect 208130 714784 208186 714793
rect 208144 714674 208172 714784
rect 208132 714668 208184 714674
rect 208132 714610 208184 714616
rect 208236 714106 208264 715550
rect 209972 714668 210024 714674
rect 209972 714610 210024 714616
rect 208144 714078 208264 714106
rect 208144 711478 208172 714078
rect 208130 711469 208186 711478
rect 208130 711404 208186 711413
rect 208144 711342 208172 711404
rect 208132 711336 208184 711342
rect 208132 711278 208184 711284
rect 208144 709143 208172 711278
rect 208130 709134 208186 709143
rect 208130 709069 208186 709078
rect 208866 709060 208922 709069
rect 208866 708995 208922 709004
rect 208130 704785 208186 704794
rect 208130 704720 208186 704729
rect 208144 701962 208172 704720
rect 208222 703008 208278 703017
rect 208222 702943 208278 702952
rect 208057 701934 208172 701962
rect 208057 640758 208085 701934
rect 208236 700302 208264 702943
rect 208222 700293 208278 700302
rect 208222 700228 208278 700237
rect 208236 699212 208264 700228
rect 208222 699203 208278 699212
rect 208222 699138 208278 699147
rect 208880 698733 208908 708995
rect 209984 707301 210012 714610
rect 209970 707292 210026 707301
rect 209970 707227 210026 707236
rect 209984 703357 210012 707227
rect 209970 703348 210026 703357
rect 209970 703283 210026 703292
rect 210432 699368 210484 699374
rect 210432 699310 210484 699316
rect 209970 699132 210026 699141
rect 209970 699067 210026 699076
rect 208866 698724 208922 698733
rect 208866 698659 208922 698668
rect 208222 695432 208278 695441
rect 208222 695367 208278 695376
rect 208130 694387 208186 694396
rect 208130 694322 208186 694331
rect 208144 694002 208172 694322
rect 208132 693996 208184 694002
rect 208132 693938 208184 693944
rect 208130 693889 208186 693898
rect 208130 693824 208186 693833
rect 208144 692574 208172 693824
rect 208132 692568 208184 692574
rect 208132 692510 208184 692516
rect 208236 691594 208264 695367
rect 208316 693996 208368 694002
rect 208316 693938 208368 693944
rect 208328 691797 208356 693938
rect 208314 691788 208370 691797
rect 208314 691723 208370 691732
rect 208222 691585 208278 691594
rect 208222 691520 208278 691529
rect 208236 691178 208264 691520
rect 208222 691169 208278 691178
rect 208222 691104 208278 691113
rect 208132 677608 208184 677614
rect 208132 677550 208184 677556
rect 208144 676226 208172 677550
rect 208880 676429 208908 698659
rect 209984 695469 210012 699067
rect 209970 695460 210026 695469
rect 209970 695395 210026 695404
rect 208960 692568 209012 692574
rect 208960 692510 209012 692516
rect 208866 676420 208922 676429
rect 208222 676385 208278 676394
rect 208866 676355 208922 676364
rect 208222 676320 208278 676329
rect 208130 676217 208186 676226
rect 208130 676152 208186 676161
rect 208144 675599 208172 676152
rect 208130 675590 208186 675599
rect 208130 675525 208186 675534
rect 208144 672250 208172 675525
rect 208236 675458 208264 676320
rect 208222 675449 208278 675458
rect 208222 675384 208278 675393
rect 208130 672241 208186 672250
rect 208130 672176 208186 672185
rect 208130 672068 208186 672077
rect 208130 672003 208186 672012
rect 208144 669862 208172 672003
rect 208132 669856 208184 669862
rect 208132 669798 208184 669804
rect 208130 669729 208186 669738
rect 208236 669715 208264 675384
rect 208314 672241 208370 672250
rect 208314 672176 208370 672185
rect 208186 669687 208264 669715
rect 208130 669664 208186 669673
rect 208144 667346 208172 669664
rect 208328 668103 208356 672176
rect 208314 668094 208370 668103
rect 208314 668029 208370 668038
rect 208328 667933 208356 668029
rect 208314 667924 208370 667933
rect 208314 667859 208370 667868
rect 208328 667738 208356 667859
rect 208236 667710 208356 667738
rect 208132 667340 208184 667346
rect 208132 667282 208184 667288
rect 208236 665396 208264 667710
rect 208222 665387 208278 665396
rect 208222 665322 208278 665331
rect 208130 663949 208186 663958
rect 208236 663935 208264 665322
rect 208186 663907 208264 663935
rect 208130 663884 208186 663893
rect 208144 660902 208172 663884
rect 208130 660893 208186 660902
rect 208130 660828 208186 660837
rect 208144 659811 208172 660828
rect 208130 659802 208186 659811
rect 208130 659737 208186 659746
rect 208144 656041 208172 659737
rect 208130 656032 208186 656041
rect 208130 655967 208186 655976
rect 208972 655594 209000 692510
rect 209326 691788 209382 691797
rect 209326 691723 209382 691732
rect 209052 669856 209104 669862
rect 209052 669798 209104 669804
rect 209064 665306 209092 669798
rect 209340 667618 209368 691723
rect 209970 691108 210026 691117
rect 209970 691043 210026 691052
rect 209984 677614 210012 691043
rect 209972 677608 210024 677614
rect 209972 677550 210024 677556
rect 209328 667612 209380 667618
rect 209328 667554 209380 667560
rect 210156 667612 210208 667618
rect 210156 667554 210208 667560
rect 210064 667340 210116 667346
rect 210064 667282 210116 667288
rect 209052 665300 209104 665306
rect 209052 665242 209104 665248
rect 208880 655566 209000 655594
rect 208130 654989 208186 654998
rect 208130 654924 208186 654933
rect 208144 652325 208172 654924
rect 208880 654397 208908 655566
rect 208866 654388 208922 654397
rect 208866 654323 208922 654332
rect 208130 652316 208186 652325
rect 208130 652251 208186 652260
rect 208130 652183 208186 652192
rect 208130 652118 208186 652127
rect 208144 651728 208172 652118
rect 208130 651719 208186 651728
rect 208130 651654 208186 651663
rect 208408 646804 208460 646810
rect 208408 646746 208460 646752
rect 208316 645036 208368 645042
rect 208316 644978 208368 644984
rect 208040 640752 208092 640758
rect 208040 640694 208092 640700
rect 208224 640344 208276 640350
rect 208224 640286 208276 640292
rect 208236 639942 208264 640286
rect 208224 639936 208276 639942
rect 208224 639878 208276 639884
rect 208328 639278 208356 644978
rect 208420 640138 208448 646746
rect 208684 640752 208736 640758
rect 208684 640694 208736 640700
rect 208592 640684 208644 640690
rect 208592 640626 208644 640632
rect 208420 640110 208540 640138
rect 208328 639250 208448 639278
rect 208144 639114 208356 639142
rect 208144 639074 208172 639114
rect 207962 639046 208172 639074
rect 208222 639020 208278 639029
rect 208040 638984 208092 638990
rect 208222 638955 208278 638964
rect 208040 638926 208092 638932
rect 208052 638666 208080 638926
rect 207962 638638 208080 638666
rect 208040 636536 208092 636542
rect 207962 636484 208040 636507
rect 207962 636479 208092 636484
rect 208040 636478 208092 636479
rect 208052 633414 208080 636478
rect 208236 633782 208264 638955
rect 208328 636610 208356 639114
rect 208420 638893 208448 639250
rect 208406 638884 208462 638893
rect 208406 638819 208462 638828
rect 208420 636678 208448 638819
rect 208408 636672 208460 636678
rect 208408 636614 208460 636620
rect 208316 636604 208368 636610
rect 208316 636546 208368 636552
rect 208512 636542 208540 640110
rect 208500 636536 208552 636542
rect 208500 636478 208552 636484
rect 208236 633754 208422 633782
rect 208052 633386 208156 633414
rect 208012 633123 208064 633128
rect 207948 633122 208064 633123
rect 207948 633071 208012 633122
rect 208012 633064 208064 633070
rect 208128 632856 208156 633386
rect 208230 633120 208282 633126
rect 208230 633062 208282 633068
rect 208052 632828 208156 632856
rect 208052 632189 208080 632828
rect 208242 632774 208270 633062
rect 207962 632161 208080 632189
rect 208052 632054 208080 632161
rect 208144 632746 208270 632774
rect 208040 632048 208092 632054
rect 208040 631990 208092 631996
rect 208144 631102 208172 632746
rect 208394 632678 208422 633754
rect 208236 632650 208422 632678
rect 208236 632258 208264 632650
rect 208224 632252 208276 632258
rect 208224 632194 208276 632200
rect 208604 632190 208632 640626
rect 208696 636814 208724 640694
rect 208880 640350 208908 654323
rect 208960 652108 209012 652114
rect 208960 652050 209012 652056
rect 208972 651677 209000 652050
rect 208958 651668 209014 651677
rect 208958 651603 209014 651612
rect 208868 640344 208920 640350
rect 208868 640286 208920 640292
rect 208776 639936 208828 639942
rect 208776 639878 208828 639884
rect 208684 636808 208736 636814
rect 208684 636750 208736 636756
rect 208788 636746 208816 639878
rect 208972 638990 209000 651603
rect 208960 638984 209012 638990
rect 208960 638926 209012 638932
rect 208868 636808 208920 636814
rect 208868 636750 208920 636756
rect 208776 636740 208828 636746
rect 208776 636682 208828 636688
rect 208684 636604 208736 636610
rect 208684 636546 208736 636552
rect 208776 636604 208828 636610
rect 208776 636546 208828 636552
rect 208316 632184 208368 632190
rect 208316 632126 208368 632132
rect 208592 632184 208644 632190
rect 208592 632126 208644 632132
rect 208132 631096 208184 631102
rect 208132 631038 208184 631044
rect 208040 630824 208092 630830
rect 207992 630779 208040 630814
rect 208040 630766 208092 630772
rect 208328 630302 208356 632126
rect 208500 632116 208552 632122
rect 208500 632058 208552 632064
rect 208408 631980 208460 631986
rect 208408 631922 208460 631928
rect 208052 630274 208356 630302
rect 208052 630232 208080 630274
rect 207960 630204 208080 630232
rect 208040 630076 208092 630082
rect 208040 630018 208092 630024
rect 208052 629503 208080 630018
rect 207962 629475 208080 629503
rect 208040 629328 208092 629334
rect 207960 629276 208040 629290
rect 207960 629270 208092 629276
rect 207960 629262 208080 629270
rect 208132 629124 208184 629130
rect 208132 629066 208184 629072
rect 208040 628852 208092 628858
rect 207962 628812 208040 628840
rect 208040 628794 208092 628800
rect 208144 628466 208172 629066
rect 207962 628438 208172 628466
rect 208038 628276 208094 628285
rect 208038 628211 208094 628220
rect 208052 627611 208080 628211
rect 207962 627583 208080 627611
rect 208144 626402 208172 628438
rect 207962 626374 208172 626402
rect 208144 625798 208172 626374
rect 208132 625792 208184 625798
rect 208132 625734 208184 625740
rect 208038 625705 208094 625714
rect 207962 625663 208038 625691
rect 208236 625701 208264 630274
rect 208316 630076 208368 630082
rect 208316 630018 208368 630024
rect 208222 625692 208278 625701
rect 208038 625640 208094 625649
rect 208132 625656 208184 625662
rect 208222 625627 208278 625636
rect 208132 625598 208184 625604
rect 208144 624366 208172 625598
rect 208328 624682 208356 630018
rect 208420 628586 208448 631922
rect 208408 628580 208460 628586
rect 208408 628522 208460 628528
rect 208328 624654 208448 624682
rect 207962 624338 208172 624366
rect 208052 624221 208080 624338
rect 207962 624193 208080 624221
rect 208052 623962 208080 624193
rect 208420 624166 208448 624654
rect 208408 624160 208460 624166
rect 208408 624102 208460 624108
rect 208512 624046 208540 632058
rect 208592 632048 208644 632054
rect 208592 631990 208644 631996
rect 208604 628858 208632 631990
rect 208696 630830 208724 636546
rect 208788 631986 208816 636546
rect 208776 631980 208828 631986
rect 208776 631922 208828 631928
rect 208776 631844 208828 631850
rect 208776 631786 208828 631792
rect 208684 630824 208736 630830
rect 208684 630766 208736 630772
rect 208788 629130 208816 631786
rect 208776 629124 208828 629130
rect 208776 629066 208828 629072
rect 208592 628852 208644 628858
rect 208592 628794 208644 628800
rect 208684 628580 208736 628586
rect 208684 628522 208736 628528
rect 208590 625692 208646 625701
rect 208590 625627 208646 625636
rect 208144 624018 208540 624046
rect 208040 623956 208092 623962
rect 208040 623898 208092 623904
rect 208038 623826 208094 623835
rect 207962 623784 208038 623812
rect 208038 623761 208094 623770
rect 208040 623684 208092 623690
rect 208040 623626 208092 623632
rect 207948 611852 208000 611858
rect 207948 611794 208000 611800
rect 207960 611649 207988 611794
rect 208052 611309 208080 623626
rect 208144 611370 208172 624018
rect 208224 623956 208276 623962
rect 208224 623898 208276 623904
rect 208236 611431 208264 623898
rect 208408 623888 208460 623894
rect 208408 623830 208460 623836
rect 208316 623820 208368 623826
rect 208316 623762 208368 623768
rect 208328 611536 208356 623762
rect 208420 611696 208448 623830
rect 208500 611784 208552 611790
rect 208500 611726 208552 611732
rect 208408 611690 208460 611696
rect 208512 611658 208540 611726
rect 208408 611632 208460 611638
rect 208498 611649 208554 611658
rect 208498 611584 208554 611593
rect 208314 611527 208370 611536
rect 208370 611485 208448 611513
rect 208314 611462 208370 611471
rect 208236 611403 208360 611431
rect 208144 611342 208299 611370
rect 208052 611281 208200 611309
rect 207985 611229 208101 611250
rect 207985 611222 208049 611229
rect 208049 611171 208101 611177
rect 208172 611012 208200 611281
rect 208051 610984 208200 611012
rect 208052 609206 208080 610984
rect 208271 610944 208299 611342
rect 208144 610916 208299 610944
rect 208040 609200 208092 609206
rect 208040 609142 208092 609148
rect 207962 609079 208080 609107
rect 208052 605822 208080 609079
rect 208144 608594 208172 610916
rect 208332 610878 208360 611403
rect 208236 610850 208360 610878
rect 208236 609226 208264 610850
rect 208236 609198 208356 609226
rect 208132 608588 208184 608594
rect 208132 608530 208184 608536
rect 208224 608248 208276 608254
rect 208224 608190 208276 608196
rect 208052 605794 208172 605822
rect 208038 605725 208094 605734
rect 207962 605683 208038 605711
rect 208038 605660 208094 605669
rect 208144 604789 208172 605794
rect 208236 604893 208264 608190
rect 208328 604920 208356 609198
rect 208420 605058 208448 611485
rect 208500 611256 208552 611262
rect 208500 611198 208552 611204
rect 208512 608254 208540 611198
rect 208500 608248 208552 608254
rect 208500 608190 208552 608196
rect 208408 605052 208460 605058
rect 208408 604994 208460 605000
rect 208222 604884 208278 604893
rect 208328 604892 208540 604920
rect 208222 604819 208278 604828
rect 207962 604761 208356 604789
rect 208215 604673 208224 604729
rect 208280 604673 208289 604729
rect 208038 603432 208094 603441
rect 207962 603390 208038 603418
rect 208038 603367 208094 603376
rect 208040 603284 208092 603290
rect 208040 603226 208092 603232
rect 208052 602830 208080 603226
rect 207962 602802 208080 602830
rect 208038 602117 208094 602126
rect 207962 602075 208038 602103
rect 208038 602052 208094 602061
rect 208236 601878 208264 604673
rect 207962 601850 208264 601878
rect 208040 601448 208092 601454
rect 207962 601408 208040 601436
rect 208040 601390 208092 601396
rect 208236 601062 208264 601850
rect 208328 601454 208356 604761
rect 208408 604780 208460 604786
rect 208408 604722 208460 604728
rect 208420 601498 208448 604722
rect 208512 602173 208540 604892
rect 208604 603290 208632 625627
rect 208696 623826 208724 628522
rect 208684 623820 208736 623826
rect 208684 623762 208736 623768
rect 208880 623690 208908 636750
rect 208972 635658 209000 638926
rect 208960 635652 209012 635658
rect 208960 635594 209012 635600
rect 208972 632229 209000 635594
rect 208958 632220 209014 632229
rect 208958 632155 209014 632164
rect 208972 631850 209000 632155
rect 208960 631844 209012 631850
rect 208960 631786 209012 631792
rect 208960 631096 209012 631102
rect 208960 631038 209012 631044
rect 208972 623797 209000 631038
rect 208958 623788 209014 623797
rect 208958 623723 209014 623732
rect 208868 623684 208920 623690
rect 208868 623626 208920 623632
rect 208684 611852 208736 611858
rect 208684 611794 208736 611800
rect 208696 609245 208724 611794
rect 208682 609236 208738 609245
rect 208682 609171 208738 609180
rect 208776 608588 208828 608594
rect 208776 608530 208828 608536
rect 208592 603284 208644 603290
rect 208644 603232 208724 603238
rect 208592 603226 208724 603232
rect 208604 603210 208724 603226
rect 208498 602164 208554 602173
rect 208498 602099 208554 602108
rect 208512 601606 208540 602099
rect 208512 601578 208632 601606
rect 208420 601470 208540 601498
rect 208316 601448 208368 601454
rect 208316 601390 208368 601396
rect 207962 601034 208264 601062
rect 208038 600225 208094 600234
rect 207962 600183 208038 600211
rect 208038 600160 208094 600169
rect 208144 599158 208172 601034
rect 208052 599130 208172 599158
rect 208052 599002 208080 599130
rect 207962 598974 208080 599002
rect 208052 598870 208080 598974
rect 208132 599000 208184 599006
rect 208132 598942 208184 598948
rect 208040 598864 208092 598870
rect 208040 598806 208092 598812
rect 207962 598263 208080 598291
rect 208052 597850 208080 598263
rect 208040 597844 208092 597850
rect 208040 597786 208092 597792
rect 208144 597118 208172 598942
rect 208512 598186 208540 601470
rect 208328 598158 208540 598186
rect 208144 597090 208264 597118
rect 207962 596938 208080 596966
rect 208052 596830 208080 596938
rect 208040 596824 208092 596830
rect 207962 596793 208040 596821
rect 208040 596766 208092 596772
rect 208038 596426 208094 596435
rect 207962 596384 208038 596412
rect 208038 596361 208094 596370
rect 208236 595214 208264 597090
rect 208144 595186 208264 595214
rect 208144 585474 208172 595186
rect 208224 595124 208276 595130
rect 208224 595066 208276 595072
rect 208132 585468 208184 585474
rect 208132 585410 208184 585416
rect 207962 584249 208172 584277
rect 208040 583904 208092 583910
rect 207962 583864 208040 583892
rect 207962 583834 207990 583864
rect 208040 583846 208092 583852
rect 208144 582730 208172 584249
rect 208052 582702 208172 582730
rect 208052 581802 208080 582702
rect 208040 581796 208092 581802
rect 208040 581738 208092 581744
rect 207962 581679 208172 581707
rect 208040 578396 208092 578402
rect 208040 578323 208092 578344
rect 207988 578271 208092 578323
rect 208144 577398 208172 581679
rect 208236 577518 208264 595066
rect 208328 584085 208356 598158
rect 208500 597844 208552 597850
rect 208500 597786 208552 597792
rect 208406 596452 208462 596461
rect 208406 596387 208462 596396
rect 208420 585542 208448 596387
rect 208512 593770 208540 597786
rect 208604 595130 208632 601578
rect 208696 597850 208724 603210
rect 208788 599006 208816 608530
rect 208776 599000 208828 599006
rect 208776 598942 208828 598948
rect 208776 598864 208828 598870
rect 208776 598806 208828 598812
rect 208684 597844 208736 597850
rect 208684 597786 208736 597792
rect 208788 596830 208816 598806
rect 208776 596824 208828 596830
rect 208776 596766 208828 596772
rect 208592 595124 208644 595130
rect 208592 595066 208644 595072
rect 208512 593742 208632 593770
rect 208408 585536 208460 585542
rect 208408 585478 208460 585484
rect 208314 584076 208370 584085
rect 208314 584011 208370 584020
rect 208328 578878 208356 584011
rect 208604 581886 208632 593742
rect 208788 583910 208816 596766
rect 208776 583904 208828 583910
rect 208776 583846 208828 583852
rect 208788 582730 208816 583846
rect 208788 582702 208908 582730
rect 208604 581858 208816 581886
rect 208500 581796 208552 581802
rect 208500 581738 208552 581744
rect 208316 578872 208368 578878
rect 208316 578814 208368 578820
rect 208224 577512 208276 577518
rect 208224 577454 208276 577460
rect 207962 577370 208172 577398
rect 208144 577262 208172 577370
rect 208144 577234 208448 577262
rect 208224 577172 208276 577178
rect 208224 577114 208276 577120
rect 208038 576032 208094 576041
rect 207962 575990 208038 576018
rect 208038 575967 208094 575976
rect 208038 575440 208094 575449
rect 207962 575398 208038 575426
rect 208038 575375 208094 575384
rect 208040 575268 208092 575274
rect 208040 575210 208092 575216
rect 208052 575002 208080 575210
rect 208040 574996 208092 575002
rect 208040 574938 208092 574944
rect 208236 574798 208264 577114
rect 208314 575372 208370 575381
rect 208314 575307 208370 575316
rect 208328 575206 208356 575307
rect 208316 575200 208368 575206
rect 208316 575142 208368 575148
rect 208224 574792 208276 574798
rect 208224 574734 208276 574740
rect 208236 574703 208264 574734
rect 207962 574675 208264 574703
rect 208328 574594 208356 575142
rect 208316 574588 208368 574594
rect 208316 574530 208368 574536
rect 208038 574504 208094 574513
rect 207962 574462 208038 574490
rect 208038 574439 208094 574448
rect 208038 574052 208094 574061
rect 207962 574010 208038 574038
rect 208420 574021 208448 577234
rect 208512 576061 208540 581738
rect 208592 578872 208644 578878
rect 208592 578814 208644 578820
rect 208498 576052 208554 576061
rect 208498 575987 208554 575996
rect 208604 575426 208632 578814
rect 208684 578396 208736 578402
rect 208684 578338 208736 578344
rect 208512 575398 208632 575426
rect 208512 575274 208540 575398
rect 208696 575358 208724 578338
rect 208604 575330 208724 575358
rect 208500 575268 208552 575274
rect 208500 575210 208552 575216
rect 208500 574588 208552 574594
rect 208500 574530 208552 574536
rect 208038 573987 208094 573996
rect 208406 574012 208462 574021
rect 208406 573947 208462 573956
rect 207962 573642 208080 573658
rect 207962 573636 208092 573642
rect 207962 573630 208040 573636
rect 208040 573578 208092 573584
rect 207962 572783 208172 572811
rect 208144 571670 208172 572783
rect 208224 571800 208276 571806
rect 208224 571742 208276 571748
rect 208132 571664 208184 571670
rect 208038 571616 208094 571625
rect 207962 571574 208038 571602
rect 208132 571606 208184 571612
rect 208038 571551 208094 571560
rect 208236 570891 208264 571742
rect 207962 570863 208356 570891
rect 208224 570780 208276 570786
rect 208224 570722 208276 570728
rect 207962 569550 208080 569578
rect 208052 569421 208080 569550
rect 207962 569393 208080 569421
rect 208052 569222 208080 569393
rect 208040 569216 208092 569222
rect 208040 569158 208092 569164
rect 208132 569148 208184 569154
rect 208132 569090 208184 569096
rect 208144 569012 208172 569090
rect 207962 568984 208172 569012
rect 208040 568808 208092 568814
rect 208040 568750 208092 568756
rect 208052 556982 208080 568750
rect 208144 567794 208172 568984
rect 208132 567788 208184 567794
rect 208132 567730 208184 567736
rect 208132 566700 208184 566706
rect 208132 566642 208184 566648
rect 208144 557730 208172 566642
rect 208132 557724 208184 557730
rect 208132 557666 208184 557672
rect 208040 556976 208092 556982
rect 208040 556918 208092 556924
rect 207962 556849 208172 556877
rect 208040 556772 208092 556778
rect 208040 556714 208092 556720
rect 208052 556686 208080 556714
rect 208038 556677 208094 556686
rect 208038 556612 208094 556621
rect 208040 556568 208092 556574
rect 208040 556510 208092 556516
rect 208052 556454 208080 556510
rect 207962 556426 208080 556454
rect 207962 554279 208080 554307
rect 208052 551018 208080 554279
rect 208144 552358 208172 556849
rect 208236 554398 208264 570722
rect 208328 554466 208356 570863
rect 208420 556302 208448 573947
rect 208512 571806 208540 574530
rect 208500 571800 208552 571806
rect 208500 571742 208552 571748
rect 208500 571664 208552 571670
rect 208500 571606 208552 571612
rect 208512 557866 208540 571606
rect 208604 569154 208632 575330
rect 208788 575206 208816 581858
rect 208880 580850 208908 582702
rect 208868 580844 208920 580850
rect 208868 580786 208920 580792
rect 208880 577421 208908 580786
rect 208866 577412 208922 577421
rect 208866 577347 208922 577356
rect 208776 575200 208828 575206
rect 208776 575142 208828 575148
rect 208880 575086 208908 577347
rect 208696 575058 208908 575086
rect 208696 574934 208724 575058
rect 208776 574996 208828 575002
rect 208776 574938 208828 574944
rect 208684 574928 208736 574934
rect 208684 574870 208736 574876
rect 208684 574792 208736 574798
rect 208684 574734 208736 574740
rect 208696 570786 208724 574734
rect 208684 570780 208736 570786
rect 208684 570722 208736 570728
rect 208684 569216 208736 569222
rect 208684 569158 208736 569164
rect 208592 569148 208644 569154
rect 208592 569090 208644 569096
rect 208500 557860 208552 557866
rect 208500 557802 208552 557808
rect 208500 557724 208552 557730
rect 208500 557666 208552 557672
rect 208408 556296 208460 556302
rect 208408 556238 208460 556244
rect 208316 554460 208368 554466
rect 208316 554402 208368 554408
rect 208224 554392 208276 554398
rect 208224 554334 208276 554340
rect 208224 553440 208276 553446
rect 208224 553382 208276 553388
rect 208132 552352 208184 552358
rect 208132 552294 208184 552300
rect 208052 550990 208168 551018
rect 208040 550923 208092 550924
rect 207948 550918 208092 550923
rect 207948 550871 208040 550918
rect 208040 550860 208092 550866
rect 208140 550792 208168 550990
rect 208052 550764 208168 550792
rect 208052 549994 208080 550764
rect 208130 550134 208186 550143
rect 208236 550120 208264 553382
rect 208512 551818 208540 557666
rect 208696 556574 208724 569158
rect 208788 568814 208816 574938
rect 208868 574928 208920 574934
rect 208868 574870 208920 574876
rect 208880 574565 208908 574870
rect 208866 574556 208922 574565
rect 208866 574491 208922 574500
rect 208880 573642 208908 574491
rect 208868 573636 208920 573642
rect 208868 573578 208920 573584
rect 208880 571573 208908 573578
rect 208866 571564 208922 571573
rect 208866 571499 208922 571508
rect 208880 569222 208908 571499
rect 208868 569216 208920 569222
rect 208868 569158 208920 569164
rect 208776 568808 208828 568814
rect 208776 568750 208828 568756
rect 209064 566706 209092 665242
rect 210076 659429 210104 667282
rect 210168 665170 210196 667554
rect 210156 665164 210208 665170
rect 210156 665106 210208 665112
rect 210062 659420 210118 659429
rect 210062 659355 210118 659364
rect 210076 658678 210104 659355
rect 209762 658661 210104 658678
rect 209762 658153 209784 658661
rect 210076 658153 210104 658661
rect 209762 658139 210104 658153
rect 209142 656020 209198 656029
rect 209142 655955 209198 655964
rect 209156 652114 209184 655955
rect 209972 652312 210024 652318
rect 209972 652254 210024 652260
rect 209144 652108 209196 652114
rect 209144 652050 209196 652056
rect 209420 644016 209472 644022
rect 209420 643958 209472 643964
rect 209328 638440 209380 638446
rect 209328 638382 209380 638388
rect 209144 636740 209196 636746
rect 209144 636682 209196 636688
rect 209156 630082 209184 636682
rect 209144 630076 209196 630082
rect 209144 630018 209196 630024
rect 209340 613053 209368 638382
rect 209326 613044 209382 613053
rect 209326 612979 209382 612988
rect 209328 601448 209380 601454
rect 209328 601390 209380 601396
rect 209052 566700 209104 566706
rect 209052 566642 209104 566648
rect 208960 556976 209012 556982
rect 208960 556918 209012 556924
rect 208684 556568 208736 556574
rect 208684 556510 208736 556516
rect 208696 553446 208724 556510
rect 208776 554460 208828 554466
rect 208776 554402 208828 554408
rect 208684 553440 208736 553446
rect 208684 553382 208736 553388
rect 208684 552352 208736 552358
rect 208684 552294 208736 552300
rect 208186 550092 208264 550120
rect 208328 551790 208540 551818
rect 208130 550069 208186 550078
rect 207962 549978 208080 549994
rect 207962 549972 208092 549978
rect 207962 549966 208040 549972
rect 208040 549914 208092 549920
rect 208052 549883 208080 549914
rect 208040 549496 208092 549502
rect 208040 549438 208092 549444
rect 208052 548618 208080 549438
rect 207962 548590 208080 548618
rect 208040 548068 208092 548074
rect 207962 548016 208040 548022
rect 207962 548010 208092 548016
rect 207962 547994 208080 548010
rect 208040 547728 208092 547734
rect 208040 547670 208092 547676
rect 208052 547303 208080 547670
rect 207962 547275 208080 547303
rect 208144 547172 208172 550069
rect 208224 549972 208276 549978
rect 208224 549914 208276 549920
rect 208052 547144 208172 547172
rect 208052 547090 208080 547144
rect 207962 547062 208080 547090
rect 208052 546821 208080 547062
rect 208038 546812 208094 546821
rect 208038 546747 208094 546756
rect 208236 546646 208264 549914
rect 208040 546640 208092 546646
rect 207962 546600 208040 546628
rect 208040 546582 208092 546588
rect 208224 546640 208276 546646
rect 208224 546582 208276 546588
rect 208038 546540 208094 546549
rect 208328 546526 208356 551790
rect 208500 550918 208552 550924
rect 208500 550860 208552 550866
rect 208408 548068 208460 548074
rect 208408 548010 208460 548016
rect 208038 546475 208094 546484
rect 208144 546498 208356 546526
rect 208052 546254 208080 546475
rect 207962 546238 208080 546254
rect 207962 546232 208092 546238
rect 207962 546226 208040 546232
rect 208040 546174 208092 546180
rect 208052 546143 208080 546174
rect 208038 545425 208094 545434
rect 207962 545383 208038 545411
rect 208038 545360 208094 545369
rect 208038 544228 208094 544237
rect 207960 544174 208038 544202
rect 208038 544163 208094 544172
rect 208040 544124 208092 544130
rect 208040 544066 208092 544072
rect 208052 543926 208080 544066
rect 208040 543920 208092 543926
rect 208040 543862 208092 543868
rect 208144 543534 208172 546498
rect 208224 546436 208276 546442
rect 208224 546378 208276 546384
rect 208236 543670 208264 546378
rect 208420 543994 208448 548010
rect 208408 543988 208460 543994
rect 208408 543930 208460 543936
rect 208236 543642 208448 543670
rect 208038 543505 208094 543514
rect 208144 543506 208356 543534
rect 207962 543463 208038 543491
rect 208038 543440 208094 543449
rect 207962 542146 208080 542174
rect 208052 542022 208080 542146
rect 208040 542021 208092 542022
rect 207962 542016 208092 542021
rect 207962 541993 208040 542016
rect 208040 541958 208092 541964
rect 208328 541682 208356 543506
rect 208316 541676 208368 541682
rect 208038 541626 208094 541635
rect 207962 541584 208038 541612
rect 208316 541618 208368 541624
rect 208038 541561 208094 541570
rect 208224 541608 208276 541614
rect 208224 541550 208276 541556
rect 208236 540406 208264 541550
rect 208144 540378 208264 540406
rect 208040 540248 208092 540254
rect 208040 540190 208092 540196
rect 208052 529549 208080 540190
rect 208038 529540 208094 529549
rect 208038 529475 208094 529484
rect 208040 529232 208092 529238
rect 208040 529174 208092 529180
rect 208052 529050 208080 529174
rect 208144 529170 208172 540378
rect 208420 540270 208448 543642
rect 208512 541653 208540 550860
rect 208696 549502 208724 552294
rect 208684 549496 208736 549502
rect 208684 549438 208736 549444
rect 208788 548074 208816 554402
rect 208868 554392 208920 554398
rect 208868 554334 208920 554340
rect 208776 548068 208828 548074
rect 208776 548010 208828 548016
rect 208880 547734 208908 554334
rect 208868 547728 208920 547734
rect 208868 547670 208920 547676
rect 208880 546442 208908 547670
rect 208868 546436 208920 546442
rect 208868 546378 208920 546384
rect 208776 546232 208828 546238
rect 208776 546174 208828 546180
rect 208788 544237 208816 546174
rect 208774 544228 208830 544237
rect 208774 544163 208830 544172
rect 208592 543988 208644 543994
rect 208592 543930 208644 543936
rect 208604 543557 208632 543930
rect 208684 543920 208736 543926
rect 208684 543862 208736 543868
rect 208590 543548 208646 543557
rect 208590 543483 208646 543492
rect 208498 541644 208554 541653
rect 208498 541579 208554 541588
rect 208236 540242 208448 540270
rect 208236 529170 208264 540242
rect 208512 540186 208540 541579
rect 208500 540180 208552 540186
rect 208500 540122 208552 540128
rect 208604 539998 208632 543483
rect 208696 540254 208724 543862
rect 208788 542022 208816 544163
rect 208972 544130 209000 556918
rect 208960 544124 209012 544130
rect 208960 544066 209012 544072
rect 208776 542016 208828 542022
rect 208776 541958 208828 541964
rect 208684 540248 208736 540254
rect 208684 540190 208736 540196
rect 208512 539970 208632 539998
rect 208512 536362 208540 539970
rect 208788 536362 208816 541958
rect 208420 536334 208540 536362
rect 208604 536334 208816 536362
rect 208132 529164 208184 529170
rect 208132 529106 208184 529112
rect 208224 529164 208276 529170
rect 208224 529106 208276 529112
rect 207962 529022 208080 529050
rect 208052 527062 208080 529022
rect 208132 528960 208184 528966
rect 208132 528902 208184 528908
rect 208224 528960 208276 528966
rect 208224 528902 208276 528908
rect 208040 527056 208092 527062
rect 208040 526998 208092 527004
rect 208038 526921 208094 526930
rect 207962 526879 208038 526907
rect 208038 526856 208094 526865
rect 208052 523778 208080 526856
rect 208144 523844 208172 528902
rect 208236 527062 208264 528902
rect 208420 528634 208448 536334
rect 208604 529238 208632 536334
rect 208682 529278 208738 529287
rect 208592 529232 208644 529238
rect 208682 529213 208738 529222
rect 208592 529174 208644 529180
rect 208328 528606 208448 528634
rect 208224 527056 208276 527062
rect 208224 526998 208276 527004
rect 208224 526920 208276 526926
rect 208224 526862 208276 526868
rect 208236 526042 208264 526862
rect 208224 526036 208276 526042
rect 208224 525978 208276 525984
rect 208236 523925 208264 525978
rect 208328 524008 208356 528606
rect 208592 527056 208644 527062
rect 208592 526998 208644 527004
rect 208328 523980 208436 524008
rect 208236 523897 208344 523925
rect 208144 523816 208252 523844
rect 208052 523750 208160 523778
rect 208023 523523 208075 523525
rect 207948 523519 208075 523523
rect 207948 523471 208023 523519
rect 208023 523461 208075 523467
rect 208035 523453 208063 523461
rect 208132 523209 208160 523750
rect 208052 523181 208160 523209
rect 208052 522874 208080 523181
rect 208224 523149 208252 523816
rect 208316 523519 208344 523897
rect 208309 523513 208361 523519
rect 208309 523455 208361 523461
rect 208145 523121 208252 523149
rect 208316 523447 208349 523455
rect 208145 522989 208173 523121
rect 208316 523082 208344 523447
rect 208144 522975 208173 522989
rect 208236 523054 208344 523082
rect 208040 522868 208092 522874
rect 208040 522810 208092 522816
rect 207962 522562 208079 522590
rect 208051 522458 208079 522562
rect 208031 522406 208037 522458
rect 208089 522406 208095 522458
rect 208144 520738 208172 522975
rect 208236 522613 208264 523054
rect 208328 522988 208356 522989
rect 208408 522988 208436 523980
rect 208328 522960 208436 522988
rect 208222 522604 208278 522613
rect 208222 522539 208278 522548
rect 208224 521344 208276 521350
rect 208224 521286 208276 521292
rect 208236 520806 208264 521286
rect 208224 520800 208276 520806
rect 208224 520742 208276 520748
rect 208132 520732 208184 520738
rect 208132 520674 208184 520680
rect 208328 520632 208356 522960
rect 208498 522604 208554 522613
rect 208498 522539 208554 522548
rect 208408 522364 208460 522370
rect 208408 522306 208460 522312
rect 207962 520604 208356 520632
rect 207962 519875 208080 519903
rect 208052 519718 208080 519875
rect 208040 519712 208092 519718
rect 207980 519598 208008 519690
rect 208040 519654 208092 519660
rect 207980 519582 208080 519598
rect 207980 519576 208092 519582
rect 207980 519570 208040 519576
rect 208040 519518 208092 519524
rect 208038 519476 208094 519485
rect 207980 519434 208038 519462
rect 207980 519210 208008 519434
rect 208038 519411 208094 519420
rect 208236 519238 208264 520604
rect 208316 519576 208368 519582
rect 208316 519518 208368 519524
rect 208144 519210 208264 519238
rect 208038 518864 208094 518873
rect 207962 518822 208038 518850
rect 208038 518799 208094 518808
rect 208144 518222 208172 519210
rect 208328 518941 208356 519518
rect 208314 518932 208370 518941
rect 208314 518867 208370 518876
rect 208132 518216 208184 518222
rect 208132 518158 208184 518164
rect 208420 518102 208448 522306
rect 208512 520874 208540 522539
rect 208604 521350 208632 526998
rect 208696 526965 208724 529213
rect 208682 526956 208738 526965
rect 208682 526891 208738 526900
rect 208684 522868 208736 522874
rect 208684 522810 208736 522816
rect 208592 521344 208644 521350
rect 208592 521286 208644 521292
rect 208500 520868 208552 520874
rect 208500 520810 208552 520816
rect 208592 520800 208644 520806
rect 208592 520742 208644 520748
rect 208500 520732 208552 520738
rect 208500 520674 208552 520680
rect 208052 518074 208448 518102
rect 208052 518011 208080 518074
rect 207962 517983 208080 518011
rect 208316 518012 208368 518018
rect 208316 517954 208368 517960
rect 208224 517944 208276 517950
rect 208224 517886 208276 517892
rect 208040 516856 208092 516862
rect 207962 516804 208040 516810
rect 208092 516804 208172 516810
rect 207962 516782 208172 516804
rect 208144 516182 208172 516782
rect 208132 516176 208184 516182
rect 208132 516118 208184 516124
rect 208038 516105 208094 516114
rect 207962 516063 208038 516091
rect 208038 516040 208094 516049
rect 208132 516040 208184 516046
rect 208132 515982 208184 515988
rect 208144 514770 208172 515982
rect 207962 514742 208172 514770
rect 208052 514621 208080 514742
rect 208132 514680 208184 514686
rect 208132 514622 208184 514628
rect 207962 514593 208080 514621
rect 208052 514414 208080 514593
rect 208040 514408 208092 514414
rect 208040 514350 208092 514356
rect 208036 514221 208088 514227
rect 207954 514175 208036 514221
rect 208036 514163 208088 514169
rect 208144 502173 208172 514622
rect 208236 502240 208264 517886
rect 208328 516085 208356 517954
rect 208314 516076 208370 516085
rect 208314 516011 208370 516020
rect 208328 502306 208356 516011
rect 208512 514686 208540 520674
rect 208604 519718 208632 520742
rect 208592 519712 208644 519718
rect 208592 519654 208644 519660
rect 208604 517950 208632 519654
rect 208696 519485 208724 522810
rect 209200 522469 209228 522471
rect 209188 522463 209240 522469
rect 209188 522405 209240 522411
rect 208776 520868 208828 520874
rect 208776 520810 208828 520816
rect 208788 519582 208816 520810
rect 208776 519576 208828 519582
rect 208776 519518 208828 519524
rect 208682 519476 208738 519485
rect 208682 519411 208738 519420
rect 208592 517944 208644 517950
rect 208592 517886 208644 517892
rect 208500 514680 208552 514686
rect 208500 514622 208552 514628
rect 208500 514408 208552 514414
rect 208500 514350 208552 514356
rect 208512 503806 208540 514350
rect 208500 503800 208552 503806
rect 208500 503742 208552 503748
rect 208328 502275 208470 502306
rect 208236 502212 208376 502240
rect 208144 502145 208284 502173
rect 207962 502049 208216 502077
rect 208094 502006 208150 502015
rect 208094 501941 208150 501950
rect 208010 501692 208062 501698
rect 207946 501640 208010 501674
rect 207946 501622 208062 501640
rect 208108 500786 208136 501941
rect 208188 501766 208216 502049
rect 208176 501760 208228 501766
rect 208176 501702 208228 501708
rect 208052 500758 208136 500786
rect 208052 499606 208080 500758
rect 208256 500704 208284 502145
rect 208144 500676 208284 500704
rect 208144 499726 208172 500676
rect 208348 500621 208376 502212
rect 208439 502094 208470 502275
rect 208236 500593 208376 500621
rect 208236 499794 208264 500593
rect 208440 500542 208468 502094
rect 208498 501877 208554 501886
rect 208696 501863 208724 519411
rect 208788 516862 208816 519518
rect 208776 516856 208828 516862
rect 208776 516798 208828 516804
rect 208776 503800 208828 503806
rect 208776 503742 208828 503748
rect 208554 501835 208724 501863
rect 208498 501812 208554 501821
rect 208520 501760 208572 501766
rect 208520 501702 208572 501708
rect 208328 500514 208468 500542
rect 208224 499788 208276 499794
rect 208224 499730 208276 499736
rect 208132 499720 208184 499726
rect 208132 499662 208184 499668
rect 208052 499578 208264 499606
rect 208038 499521 208094 499530
rect 207962 499479 208038 499507
rect 208038 499456 208094 499465
rect 208132 498564 208184 498570
rect 208132 498506 208184 498512
rect 208038 496125 208094 496134
rect 207962 496083 208038 496111
rect 208038 496060 208094 496069
rect 208040 495980 208092 495986
rect 208040 495922 208092 495928
rect 208052 495186 208080 495922
rect 207962 495158 208080 495186
rect 208144 493826 208172 498506
rect 207962 493798 208172 493826
rect 208236 493306 208264 499578
rect 208328 496326 208356 500514
rect 208532 500444 208560 501702
rect 208696 501102 208724 501835
rect 208788 501698 208816 503742
rect 208776 501692 208828 501698
rect 208776 501634 208828 501640
rect 208602 501074 208724 501102
rect 208602 501034 208630 501074
rect 208788 501034 208816 501634
rect 208602 501006 208632 501034
rect 208420 500413 208560 500444
rect 208420 498570 208448 500413
rect 208500 499720 208552 499726
rect 208500 499662 208552 499668
rect 208408 498564 208460 498570
rect 208408 498506 208460 498512
rect 208408 498428 208460 498434
rect 208408 498370 208460 498376
rect 208316 496320 208368 496326
rect 208316 496262 208368 496268
rect 208420 495141 208448 498370
rect 208512 495986 208540 499662
rect 208604 496444 208632 501006
rect 208696 501006 208816 501034
rect 208696 499493 208724 501006
rect 208776 499788 208828 499794
rect 208776 499730 208828 499736
rect 208682 499484 208738 499493
rect 208682 499419 208738 499428
rect 208696 498434 208724 499419
rect 208684 498428 208736 498434
rect 208684 498370 208736 498376
rect 208604 496416 208724 496444
rect 208592 496320 208644 496326
rect 208592 496262 208644 496268
rect 208500 495980 208552 495986
rect 208500 495922 208552 495928
rect 208406 495132 208462 495141
rect 208406 495067 208462 495076
rect 208236 493278 208448 493306
rect 208132 493260 208184 493266
rect 208038 493232 208094 493237
rect 207962 493228 208094 493232
rect 207962 493204 208038 493228
rect 208132 493202 208184 493208
rect 208038 493163 208094 493172
rect 208052 492654 208080 493163
rect 208040 492648 208092 492654
rect 208040 492590 208092 492596
rect 208038 492517 208094 492526
rect 207962 492475 208038 492503
rect 208038 492452 208094 492461
rect 208144 492290 208172 493202
rect 207962 492262 208172 492290
rect 208052 491838 208080 492262
rect 207962 491810 208080 491838
rect 208052 491460 208080 491810
rect 207962 491432 208080 491460
rect 208052 490614 208080 491432
rect 208040 490611 208092 490614
rect 207962 490608 208092 490611
rect 207962 490583 208040 490608
rect 208040 490550 208092 490556
rect 208420 490494 208448 493278
rect 208052 490466 208448 490494
rect 208052 489542 208080 490466
rect 208512 490410 208540 495922
rect 208604 493329 208632 496262
rect 208696 496093 208724 496416
rect 208682 496084 208738 496093
rect 208682 496019 208738 496028
rect 208682 495132 208738 495141
rect 208682 495067 208738 495076
rect 208590 493320 208646 493329
rect 208696 493266 208724 495067
rect 208590 493255 208646 493264
rect 208684 493260 208736 493266
rect 208684 493202 208736 493208
rect 208684 492648 208736 492654
rect 208684 492590 208736 492596
rect 208132 490404 208184 490410
rect 208132 490346 208184 490352
rect 208500 490404 208552 490410
rect 208500 490346 208552 490352
rect 208144 489678 208172 490346
rect 208224 490336 208276 490342
rect 208224 490278 208276 490284
rect 208236 489814 208264 490278
rect 208236 489786 208632 489814
rect 208144 489650 208540 489678
rect 208052 489514 208448 489542
rect 208040 489452 208092 489458
rect 207962 489400 208040 489406
rect 208092 489400 208172 489406
rect 207962 489378 208172 489400
rect 208052 489329 208080 489378
rect 208040 488704 208092 488710
rect 207962 488663 208040 488691
rect 208040 488646 208092 488652
rect 208144 487366 208172 489378
rect 207962 487338 208172 487366
rect 208144 487221 208172 487338
rect 207960 487208 208172 487221
rect 207960 487193 208040 487208
rect 208092 487193 208172 487208
rect 208040 487150 208092 487156
rect 208038 486826 208094 486835
rect 207962 486784 208038 486812
rect 208038 486761 208094 486770
rect 208420 486142 208448 489514
rect 208052 486114 208448 486142
rect 208052 479886 208080 486114
rect 208512 486006 208540 489650
rect 208144 485978 208540 486006
rect 208144 481654 208172 485978
rect 208604 485870 208632 489786
rect 208696 488710 208724 492590
rect 208788 492557 208816 499730
rect 208866 496084 208922 496093
rect 208866 496019 208922 496028
rect 208774 492548 208830 492557
rect 208774 492483 208830 492492
rect 208788 490342 208816 492483
rect 208776 490336 208828 490342
rect 208776 490278 208828 490284
rect 208684 488704 208736 488710
rect 208684 488646 208736 488652
rect 208236 485842 208632 485870
rect 208696 485854 208724 488646
rect 208880 486845 208908 496019
rect 208960 487208 209012 487214
rect 208960 487150 209012 487156
rect 208866 486836 208922 486845
rect 208866 486771 208922 486780
rect 208684 485848 208736 485854
rect 208236 481774 208264 485842
rect 208684 485790 208736 485796
rect 208408 485780 208460 485786
rect 208880 485734 208908 486771
rect 208408 485722 208460 485728
rect 208224 481768 208276 481774
rect 208224 481710 208276 481716
rect 208144 481626 208356 481654
rect 208224 481496 208276 481502
rect 208224 481438 208276 481444
rect 208052 479858 208172 479886
rect 207948 474668 208000 474674
rect 207948 474610 208000 474616
rect 207960 474449 207988 474610
rect 208040 474288 208092 474294
rect 208040 474230 208092 474236
rect 208052 474062 208080 474230
rect 207962 474034 208080 474062
rect 208052 471907 208080 474034
rect 207962 471879 208080 471907
rect 208052 471044 208080 471879
rect 208040 471038 208092 471044
rect 208040 470980 208092 470986
rect 208144 470418 208172 479858
rect 208236 470962 208264 481438
rect 208224 470956 208276 470962
rect 208224 470898 208276 470904
rect 208328 470894 208356 481626
rect 208420 477850 208448 485722
rect 208604 485706 208908 485734
rect 208420 477822 208540 477850
rect 208408 474668 208460 474674
rect 208408 474610 208460 474616
rect 208316 470888 208368 470894
rect 208316 470830 208368 470836
rect 208420 470774 208448 474610
rect 208328 470746 208448 470774
rect 208224 470684 208276 470690
rect 208224 470626 208276 470632
rect 208132 470412 208184 470418
rect 208132 470354 208184 470360
rect 207962 468483 208080 468511
rect 208052 467698 208080 468483
rect 208040 467692 208092 467698
rect 208040 467634 208092 467640
rect 208236 467578 208264 470626
rect 207962 467550 208264 467578
rect 208052 466338 208080 467550
rect 208040 466332 208092 466338
rect 208040 466274 208092 466280
rect 208328 466218 208356 470746
rect 208512 470536 208540 477822
rect 208604 474197 208632 485706
rect 208972 482266 209000 487150
rect 208880 482238 209000 482266
rect 208880 474294 208908 482238
rect 208868 474288 208920 474294
rect 208868 474230 208920 474236
rect 208590 474188 208646 474197
rect 208590 474123 208646 474132
rect 208866 474188 208922 474197
rect 208866 474123 208922 474132
rect 208776 470956 208828 470962
rect 208776 470898 208828 470904
rect 208420 470508 208540 470536
rect 208420 466406 208448 470508
rect 208500 470412 208552 470418
rect 208500 470354 208552 470360
rect 208408 466400 208460 466406
rect 208408 466342 208460 466348
rect 208512 466286 208540 470354
rect 207962 466190 208356 466218
rect 208420 466258 208540 466286
rect 208040 466128 208092 466134
rect 208040 466070 208092 466076
rect 208052 465632 208080 466070
rect 207962 465604 208080 465632
rect 208040 465516 208092 465522
rect 208040 465458 208092 465464
rect 208052 464903 208080 465458
rect 207962 464875 208080 464903
rect 208040 464836 208092 464842
rect 208040 464778 208092 464784
rect 208052 464690 208080 464778
rect 207962 464662 208080 464690
rect 208052 464246 208080 464662
rect 207962 464218 208080 464246
rect 208052 463860 208080 464218
rect 207962 463832 208080 463860
rect 208052 463022 208080 463832
rect 207962 462994 208080 463022
rect 208052 462870 208080 462994
rect 208040 462864 208092 462870
rect 208040 462806 208092 462812
rect 208224 461844 208276 461850
rect 208038 461812 208094 461821
rect 207962 461770 208038 461798
rect 208224 461786 208276 461792
rect 208038 461747 208094 461756
rect 208236 461091 208264 461786
rect 207962 461063 208264 461091
rect 208038 459780 208094 459789
rect 207960 459738 208038 459766
rect 208038 459715 208094 459724
rect 208038 459636 208094 459645
rect 207962 459594 208038 459622
rect 208038 459571 208094 459580
rect 207962 459198 208172 459212
rect 207962 459192 208184 459198
rect 207962 459184 208132 459192
rect 208132 459134 208184 459140
rect 208130 459096 208186 459105
rect 208130 459031 208186 459040
rect 208040 457492 208092 457498
rect 208040 457434 208092 457440
rect 207948 447254 208000 447260
rect 207948 447196 208000 447202
rect 207960 447049 207988 447196
rect 208052 446974 208080 457434
rect 208144 447570 208172 459031
rect 208132 447564 208184 447570
rect 208132 447506 208184 447512
rect 208236 447162 208264 461063
rect 208316 459124 208368 459130
rect 208316 459066 208368 459072
rect 208328 447484 208356 459066
rect 208420 457498 208448 466258
rect 208500 466196 208552 466202
rect 208500 466138 208552 466144
rect 208512 459198 208540 466138
rect 208592 466128 208644 466134
rect 208592 466070 208644 466076
rect 208604 461850 208632 466070
rect 208788 465522 208816 470898
rect 208880 467698 208908 474123
rect 209052 471024 209104 471030
rect 209052 470966 209104 470972
rect 209064 467941 209092 470966
rect 209050 467932 209106 467941
rect 209050 467867 209106 467876
rect 208868 467692 208920 467698
rect 208868 467634 208920 467640
rect 208776 465516 208828 465522
rect 208696 465476 208776 465504
rect 208592 461844 208644 461850
rect 208592 461786 208644 461792
rect 208590 459636 208646 459645
rect 208590 459571 208646 459580
rect 208500 459192 208552 459198
rect 208500 459134 208552 459140
rect 208604 459082 208632 459571
rect 208696 459373 208724 465476
rect 208776 465458 208828 465464
rect 208880 465334 208908 467634
rect 208788 465306 208908 465334
rect 208682 459364 208738 459373
rect 208682 459299 208738 459308
rect 208500 459056 208552 459062
rect 208604 459054 208724 459082
rect 208788 459062 208816 465306
rect 209064 464842 209092 467867
rect 209052 464836 209104 464842
rect 209052 464778 209104 464784
rect 209199 464623 209227 522405
rect 209098 464595 209227 464623
rect 208868 462864 208920 462870
rect 208868 462806 208920 462812
rect 208880 461821 208908 462806
rect 208866 461812 208922 461821
rect 208866 461747 208922 461756
rect 208880 459645 208908 461747
rect 208866 459636 208922 459645
rect 208866 459571 208922 459580
rect 208500 458998 208552 459004
rect 208408 457492 208460 457498
rect 208408 457434 208460 457440
rect 208512 451354 208540 458998
rect 208512 451326 208632 451354
rect 208328 447456 208540 447484
rect 208408 447254 208460 447260
rect 208408 447196 208460 447202
rect 208224 447156 208276 447162
rect 208224 447098 208276 447104
rect 208052 446946 208356 446974
rect 208224 446884 208276 446890
rect 208224 446826 208276 446832
rect 208040 446680 208092 446686
rect 207962 446634 208040 446662
rect 208040 446622 208092 446628
rect 208052 444507 208080 446622
rect 207962 444479 208080 444507
rect 208052 444442 208080 444479
rect 208040 444436 208092 444442
rect 208040 444378 208092 444384
rect 208132 441648 208184 441654
rect 208132 441590 208184 441596
rect 208038 441125 208094 441134
rect 207962 441083 208038 441111
rect 208038 441060 208094 441069
rect 208144 440189 208172 441590
rect 208236 441586 208264 446826
rect 208224 441580 208276 441586
rect 208224 441522 208276 441528
rect 208222 440334 208278 440343
rect 208222 440269 208278 440278
rect 207962 440161 208172 440189
rect 208038 438832 208094 438841
rect 207960 438790 208038 438818
rect 208038 438767 208094 438776
rect 208040 438248 208092 438254
rect 207962 438208 208040 438236
rect 208040 438190 208092 438196
rect 207962 437475 208080 437503
rect 208052 437438 208080 437475
rect 208040 437432 208092 437438
rect 208040 437374 208092 437380
rect 208144 437370 208172 440161
rect 208132 437364 208184 437370
rect 208132 437306 208184 437312
rect 207962 437262 208080 437290
rect 208052 437182 208080 437262
rect 208236 437182 208264 440269
rect 208052 437154 208264 437182
rect 208052 436842 208080 437154
rect 207962 436814 208080 436842
rect 208052 436460 208080 436814
rect 207962 436432 208080 436460
rect 208052 435618 208080 436432
rect 208328 435898 208356 446946
rect 208420 438837 208448 447196
rect 208512 441654 208540 447456
rect 208604 446861 208632 451326
rect 208590 446852 208646 446861
rect 208590 446787 208646 446796
rect 208500 441648 208552 441654
rect 208500 441590 208552 441596
rect 208604 441586 208632 446787
rect 208696 446686 208724 459054
rect 208776 459056 208828 459062
rect 208776 458998 208828 459004
rect 209098 457866 209126 464595
rect 209070 457810 209080 457866
rect 209136 457810 209146 457866
rect 208868 447564 208920 447570
rect 208868 447506 208920 447512
rect 208684 446680 208736 446686
rect 208684 446622 208736 446628
rect 208880 445070 208908 447506
rect 208696 445042 208908 445070
rect 208592 441580 208644 441586
rect 208592 441522 208644 441528
rect 208500 441444 208552 441450
rect 208500 441386 208552 441392
rect 208592 441444 208644 441450
rect 208592 441386 208644 441392
rect 208406 438828 208462 438837
rect 208406 438763 208462 438772
rect 208512 438254 208540 441386
rect 208604 441149 208632 441386
rect 208590 441140 208646 441149
rect 208590 441075 208646 441084
rect 208500 438248 208552 438254
rect 208500 438190 208552 438196
rect 208408 437364 208460 437370
rect 208408 437306 208460 437312
rect 207962 435590 208080 435618
rect 208052 434394 208080 435590
rect 207962 434366 208080 434394
rect 208052 434326 208080 434366
rect 208236 435870 208356 435898
rect 208052 434298 208172 434326
rect 208040 433692 208092 433698
rect 207962 433652 208040 433680
rect 208040 433634 208092 433640
rect 208144 432354 208172 434298
rect 207962 432326 208172 432354
rect 208052 432218 208080 432326
rect 207962 432190 208080 432218
rect 208052 432150 208080 432190
rect 208052 432122 208172 432150
rect 208038 431824 208094 431833
rect 207962 431782 208038 431810
rect 208144 431794 208172 432122
rect 208038 431759 208094 431768
rect 208132 431788 208184 431794
rect 208132 431730 208184 431736
rect 208236 431606 208264 435870
rect 208052 431578 208264 431606
rect 208052 422070 208080 431578
rect 208132 431516 208184 431522
rect 208132 431458 208184 431464
rect 208144 427442 208172 431458
rect 208420 428170 208448 437306
rect 208604 436094 208632 441075
rect 208696 437438 208724 445042
rect 208776 444436 208828 444442
rect 208776 444378 208828 444384
rect 208788 443626 208816 444378
rect 208776 443620 208828 443626
rect 208776 443562 208828 443568
rect 208788 440343 208816 443562
rect 208774 440334 208830 440343
rect 208774 440269 208830 440278
rect 208868 438248 208920 438254
rect 208868 438190 208920 438196
rect 208684 437432 208736 437438
rect 208684 437374 208736 437380
rect 208604 436066 208724 436094
rect 208696 431765 208724 436066
rect 208880 435898 208908 438190
rect 208960 437432 209012 437438
rect 208960 437374 209012 437380
rect 208788 435870 208908 435898
rect 208788 433698 208816 435870
rect 208776 433692 208828 433698
rect 208776 433634 208828 433640
rect 208972 432066 209000 437374
rect 208960 432060 209012 432066
rect 208960 432002 209012 432008
rect 208682 431756 208738 431765
rect 208682 431691 208738 431700
rect 208866 431756 208922 431765
rect 208866 431691 208922 431700
rect 208328 428142 208448 428170
rect 208132 427436 208184 427442
rect 208132 427378 208184 427384
rect 208328 422138 208356 428142
rect 208316 422132 208368 422138
rect 208316 422074 208368 422080
rect 208040 422064 208092 422070
rect 208040 422006 208092 422012
rect 207968 419202 208080 419230
rect 208052 412714 208080 419202
rect 208052 412686 208356 412714
rect 207968 411264 208080 411292
rect 208052 411206 208080 411264
rect 208132 411252 208184 411258
rect 208052 411200 208132 411206
rect 208052 411194 208184 411200
rect 208052 411178 208172 411194
rect 207968 410578 208080 410594
rect 207968 410572 208092 410578
rect 207968 410566 208040 410572
rect 208040 410514 208092 410520
rect 208040 409722 208092 409728
rect 208144 409710 208172 411178
rect 208092 409682 208172 409710
rect 208040 409664 208092 409670
rect 208052 409216 208080 409664
rect 207968 409188 208264 409216
rect 207968 408730 208080 408758
rect 208052 408622 208080 408730
rect 208236 408622 208264 409188
rect 208052 408594 208264 408622
rect 208040 408328 208092 408334
rect 208040 408270 208092 408276
rect 208052 408214 208080 408270
rect 207960 408186 208080 408214
rect 208144 407670 208172 408594
rect 208328 408334 208356 412686
rect 208316 408328 208368 408334
rect 208316 408270 208368 408276
rect 207968 407642 208172 407670
rect 208052 407586 208080 407642
rect 208040 407580 208092 407586
rect 208040 407522 208092 407528
rect 208132 407240 208184 407246
rect 207968 407188 208132 407194
rect 207968 407182 208184 407188
rect 207968 407166 208172 407182
rect 207968 406418 208080 406446
rect 208052 405546 208080 406418
rect 208040 405540 208092 405546
rect 208040 405482 208092 405488
rect 208144 400570 208172 407166
rect 208880 405546 208908 431691
rect 208868 405540 208920 405546
rect 208868 405482 208920 405488
rect 208052 400542 208172 400570
rect 208052 397258 208080 400542
rect 208052 397230 208264 397258
rect 207962 392834 208172 392862
rect 208144 390722 208172 392834
rect 208236 392842 208264 397230
rect 208880 393141 208908 405482
rect 208866 393132 208922 393141
rect 208866 393067 208922 393076
rect 208236 392814 208540 392842
rect 208132 390716 208184 390722
rect 207962 390679 208132 390707
rect 208132 390658 208184 390664
rect 208040 389832 208092 389838
rect 208040 389774 208092 389780
rect 208052 387564 208080 389774
rect 208144 387660 208172 390658
rect 208316 390444 208368 390450
rect 208316 390386 208368 390392
rect 208144 387632 208252 387660
rect 208052 387536 208160 387564
rect 208011 387323 208063 387329
rect 207948 387271 208011 387323
rect 208011 387265 208063 387271
rect 208132 387088 208160 387536
rect 208224 387333 208252 387632
rect 208221 387327 208273 387333
rect 208221 387269 208273 387275
rect 208052 387060 208160 387088
rect 208052 386386 208080 387060
rect 208224 386999 208252 387269
rect 208144 386971 208252 386999
rect 208144 386543 208172 386971
rect 208130 386534 208186 386543
rect 208130 386469 208186 386478
rect 207962 386370 208080 386386
rect 207962 386364 208092 386370
rect 207962 386358 208040 386364
rect 208040 386306 208092 386312
rect 208052 386275 208080 386306
rect 208144 385146 208172 386469
rect 208132 385140 208184 385146
rect 208328 385114 208356 390386
rect 208408 386364 208460 386370
rect 208408 386306 208460 386312
rect 208132 385082 208184 385088
rect 208236 385086 208356 385114
rect 208236 384432 208264 385086
rect 207962 384404 208264 384432
rect 208038 383717 208094 383726
rect 207962 383675 208038 383703
rect 208038 383652 208094 383661
rect 208040 383508 208092 383514
rect 207962 383462 208040 383490
rect 208040 383450 208092 383456
rect 208040 383100 208092 383106
rect 208040 383042 208092 383048
rect 208040 383038 208080 383042
rect 207962 383010 208080 383038
rect 208052 382660 208080 383010
rect 207962 382632 208080 382660
rect 208052 381811 208080 382632
rect 207962 381783 208080 381811
rect 208052 380606 208080 381783
rect 207962 380578 208080 380606
rect 208052 380050 208080 380578
rect 208052 380022 208154 380050
rect 208032 379912 208072 379914
rect 208032 379906 208084 379912
rect 207948 379854 208032 379903
rect 207948 379851 208084 379854
rect 208032 379848 208084 379851
rect 208126 379780 208154 380022
rect 208236 379926 208264 384404
rect 208420 383514 208448 386306
rect 208512 383757 208540 392814
rect 208880 389838 208908 393067
rect 208868 389832 208920 389838
rect 208868 389774 208920 389780
rect 208592 385140 208644 385146
rect 208592 385082 208644 385088
rect 208498 383748 208554 383757
rect 208498 383683 208554 383692
rect 208408 383508 208460 383514
rect 208408 383450 208460 383456
rect 208420 381966 208448 383450
rect 208328 381938 208448 381966
rect 208236 379914 208276 379926
rect 208236 379908 208288 379914
rect 208236 379850 208288 379856
rect 208052 379752 208154 379780
rect 208052 378566 208080 379752
rect 207962 378538 208080 378566
rect 208052 378430 208080 378538
rect 207962 378402 208080 378430
rect 208328 378012 208356 381938
rect 208512 381811 208540 383683
rect 208604 383106 208632 385082
rect 208592 383100 208644 383106
rect 208592 383042 208644 383048
rect 208420 381783 208540 381811
rect 208420 380658 208448 381783
rect 208408 380652 208460 380658
rect 208408 380594 208460 380600
rect 207962 377984 208356 378012
rect 208062 263086 208090 377984
rect 209340 316126 209368 601390
rect 209432 555661 209460 643958
rect 209984 640690 210012 652254
rect 210076 645042 210104 658139
rect 210168 655213 210196 665106
rect 210154 655204 210210 655213
rect 210154 655139 210210 655148
rect 210064 645036 210116 645042
rect 210064 644978 210116 644984
rect 209972 640684 210024 640690
rect 209972 640626 210024 640632
rect 209512 610900 209564 610906
rect 209512 610842 209564 610848
rect 209418 555652 209474 555661
rect 209418 555587 209474 555596
rect 209420 546640 209472 546646
rect 209420 546582 209472 546588
rect 209432 372090 209460 546582
rect 209524 522370 209552 610842
rect 209788 609200 209840 609206
rect 209788 609142 209840 609148
rect 209800 590506 209828 609142
rect 209788 590500 209840 590506
rect 209788 590442 209840 590448
rect 209694 584212 209750 584221
rect 209694 584147 209750 584156
rect 209708 583910 209736 584147
rect 209696 583904 209748 583910
rect 209696 583846 209748 583852
rect 209512 522364 209564 522370
rect 209512 522306 209564 522312
rect 210444 447133 210472 699310
rect 226248 692698 226776 692716
rect 226248 692383 226265 692698
rect 226757 692383 226776 692698
rect 226248 692366 226776 692383
rect 220034 667728 222160 667758
rect 220034 667552 220076 667728
rect 222120 667552 222160 667728
rect 220034 667516 222160 667552
rect 236436 667020 243140 667120
rect 236436 665954 236536 667020
rect 242984 665954 243140 667020
rect 236436 665890 243140 665954
rect 213466 654660 213522 654669
rect 213466 654595 213522 654604
rect 213480 654562 213508 654595
rect 213468 654556 213520 654562
rect 213468 654498 213520 654504
rect 217056 650136 217108 650142
rect 217056 650078 217108 650084
rect 211534 623788 211590 623797
rect 211534 623723 211590 623732
rect 211548 599346 211576 623723
rect 213744 614164 213796 614170
rect 213744 614106 213796 614112
rect 213756 610906 213784 614106
rect 217068 611790 217096 650078
rect 233616 647960 233668 647966
rect 233616 647902 233668 647908
rect 223680 647620 223732 647626
rect 223680 647562 223732 647568
rect 219264 647348 219316 647354
rect 219264 647290 219316 647296
rect 217056 611784 217108 611790
rect 217056 611726 217108 611732
rect 213744 610900 213796 610906
rect 213744 610842 213796 610848
rect 211536 599340 211588 599346
rect 211536 599282 211588 599288
rect 211534 556740 211590 556749
rect 211534 556675 211590 556684
rect 211168 475104 211220 475110
rect 211168 475046 211220 475052
rect 211180 474605 211208 475046
rect 211166 474596 211222 474605
rect 211166 474531 211222 474540
rect 210430 447124 210486 447133
rect 210430 447059 210486 447068
rect 209512 433692 209564 433698
rect 209512 433634 209564 433640
rect 209524 410578 209552 433634
rect 210156 432060 210208 432066
rect 210156 432002 210208 432008
rect 209972 427436 210024 427442
rect 209972 427378 210024 427384
rect 209984 411258 210012 427378
rect 209972 411252 210024 411258
rect 209972 411194 210024 411200
rect 209512 410572 209564 410578
rect 209512 410514 209564 410520
rect 210064 410572 210116 410578
rect 210064 410514 210116 410520
rect 210076 390450 210104 410514
rect 210168 407246 210196 432002
rect 210248 407580 210300 407586
rect 210248 407522 210300 407528
rect 210156 407240 210208 407246
rect 210156 407182 210208 407188
rect 210260 390722 210288 407522
rect 210248 390716 210300 390722
rect 210248 390658 210300 390664
rect 210064 390444 210116 390450
rect 210064 390386 210116 390392
rect 210432 380652 210484 380658
rect 210432 380594 210484 380600
rect 209420 372084 209472 372090
rect 209420 372026 209472 372032
rect 209328 316120 209380 316126
rect 209328 316062 209380 316068
rect 208040 263080 208092 263086
rect 208040 263022 208092 263028
rect 210444 259686 210472 380594
rect 210524 372084 210576 372090
rect 210524 372026 210576 372032
rect 210536 367738 210564 372026
rect 210524 367732 210576 367738
rect 210524 367674 210576 367680
rect 211548 279882 211576 556675
rect 214848 540180 214900 540186
rect 214848 540122 214900 540128
rect 214860 514346 214888 540122
rect 214848 514340 214900 514346
rect 214848 514282 214900 514288
rect 219276 475110 219304 647290
rect 223692 638446 223720 647562
rect 233628 644022 233656 647902
rect 241344 647008 241396 647014
rect 241344 646950 241396 646956
rect 233616 644016 233668 644022
rect 233616 643958 233668 643964
rect 223680 638440 223732 638446
rect 223680 638382 223732 638388
rect 241356 632938 241384 646950
rect 230304 632932 230356 632938
rect 230304 632874 230356 632880
rect 241344 632932 241396 632938
rect 241344 632874 241396 632880
rect 230316 626070 230344 632874
rect 228096 626064 228148 626070
rect 228096 626006 228148 626012
rect 230304 626064 230356 626070
rect 230304 626006 230356 626012
rect 228108 614170 228136 626006
rect 228096 614164 228148 614170
rect 228096 614106 228148 614112
rect 233616 605936 233668 605942
rect 233616 605878 233668 605884
rect 219356 590500 219408 590506
rect 219356 590442 219408 590448
rect 219368 576906 219396 590442
rect 219356 576900 219408 576906
rect 219356 576842 219408 576848
rect 221564 576900 221616 576906
rect 221564 576842 221616 576848
rect 221472 567788 221524 567794
rect 221472 567730 221524 567736
rect 221484 478986 221512 567730
rect 221576 565618 221604 576842
rect 221564 565612 221616 565618
rect 221564 565554 221616 565560
rect 225888 565612 225940 565618
rect 225888 565554 225940 565560
rect 225900 556914 225928 565554
rect 225888 556908 225940 556914
rect 225888 556850 225940 556856
rect 221472 478980 221524 478986
rect 221472 478922 221524 478928
rect 219264 475104 219316 475110
rect 219264 475046 219316 475052
rect 226992 422132 227044 422138
rect 226992 422074 227044 422080
rect 217056 367732 217108 367738
rect 217056 367674 217108 367680
rect 217068 357674 217096 367674
rect 217056 357668 217108 357674
rect 217056 357610 217108 357616
rect 221472 357668 221524 357674
rect 221472 357610 221524 357616
rect 221484 329318 221512 357610
rect 221472 329312 221524 329318
rect 221472 329254 221524 329260
rect 222392 329312 222444 329318
rect 222392 329254 222444 329260
rect 222404 320546 222432 329254
rect 222392 320540 222444 320546
rect 222392 320482 222444 320488
rect 217056 316120 217108 316126
rect 217056 316062 217108 316068
rect 217068 302866 217096 316062
rect 217056 302860 217108 302866
rect 217056 302802 217108 302808
rect 227004 280533 227032 422074
rect 228096 422064 228148 422070
rect 228096 422006 228148 422012
rect 228108 386302 228136 422006
rect 232236 421588 232288 421594
rect 232236 421530 232288 421536
rect 228096 386296 228148 386302
rect 228096 386238 228148 386244
rect 228108 385486 228136 386238
rect 227636 385480 227688 385486
rect 227636 385422 227688 385428
rect 228096 385480 228148 385486
rect 228096 385422 228148 385428
rect 227648 280646 227676 385422
rect 229200 302860 229252 302866
rect 229200 302802 229252 302808
rect 229212 294026 229240 302802
rect 229200 294020 229252 294026
rect 229200 293962 229252 293968
rect 231222 284740 231278 284749
rect 231222 284675 231278 284684
rect 229396 284574 229792 284590
rect 229396 284568 229804 284574
rect 229396 284562 229752 284568
rect 229752 284510 229804 284516
rect 232248 283797 232276 421530
rect 233628 284749 233656 605878
rect 244654 599580 244710 599589
rect 244654 599515 244710 599524
rect 244668 599346 244696 599515
rect 244656 599340 244708 599346
rect 244656 599282 244708 599288
rect 244654 557148 244710 557157
rect 244654 557083 244710 557092
rect 234720 556908 234772 556914
rect 234720 556850 234772 556856
rect 234732 549026 234760 556850
rect 244668 556302 244696 557083
rect 244656 556296 244708 556302
rect 244656 556238 244708 556244
rect 234720 549020 234772 549026
rect 234720 548962 234772 548968
rect 243552 549020 243604 549026
rect 243552 548962 243604 548968
rect 243564 505438 243592 548962
rect 244848 514170 244854 514222
rect 244906 514170 244913 514222
rect 243552 505432 243604 505438
rect 243552 505374 243604 505380
rect 233708 320540 233760 320546
rect 233708 320482 233760 320488
rect 233720 297494 233748 320482
rect 233708 297488 233760 297494
rect 233708 297430 233760 297436
rect 238032 297488 238084 297494
rect 238032 297430 238084 297436
rect 233708 294020 233760 294026
rect 233708 293962 233760 293968
rect 233720 287566 233748 293962
rect 238044 291034 238072 297430
rect 238032 291028 238084 291034
rect 238032 290970 238084 290976
rect 240240 291028 240292 291034
rect 240240 290970 240292 290976
rect 233708 287560 233760 287566
rect 233708 287502 233760 287508
rect 233614 284740 233670 284749
rect 233614 284675 233670 284684
rect 232328 284568 232380 284574
rect 232328 284510 232380 284516
rect 232340 284098 232368 284510
rect 232328 284092 232380 284098
rect 232328 284034 232380 284040
rect 232234 283788 232290 283797
rect 232234 283723 232290 283732
rect 227648 280618 228412 280646
rect 226990 280524 227046 280533
rect 230210 280524 230266 280533
rect 226990 280459 227046 280468
rect 229856 280482 230210 280510
rect 211536 279876 211588 279882
rect 211536 279818 211588 279824
rect 229856 266418 229884 280482
rect 230210 280459 230266 280468
rect 232156 280346 232552 280374
rect 232326 279980 232382 279989
rect 232326 279915 232382 279924
rect 232340 279134 232368 279915
rect 232524 279814 232552 280346
rect 240252 280125 240280 290970
rect 244656 287560 244708 287566
rect 244656 287502 244708 287508
rect 240238 280116 240294 280125
rect 240238 280051 240294 280060
rect 244668 279989 244696 287502
rect 244654 279980 244710 279989
rect 244654 279915 244710 279924
rect 232512 279808 232564 279814
rect 232512 279750 232564 279756
rect 232328 279128 232380 279134
rect 232328 279070 232380 279076
rect 244866 278071 244894 514170
rect 246324 316165 246352 725626
rect 246817 725504 246869 725510
rect 246817 725446 246869 725452
rect 246829 543064 246857 725446
rect 248980 700320 249032 700326
rect 248980 700262 249032 700268
rect 248152 674412 248204 674418
rect 248152 674354 248204 674360
rect 247324 656120 247376 656126
rect 247324 656062 247376 656068
rect 246784 542964 246793 543064
rect 246889 542964 246899 543064
rect 246864 505432 246916 505438
rect 246864 505374 246916 505380
rect 246876 500309 246904 505374
rect 246862 500300 246918 500309
rect 246862 500235 246918 500244
rect 247336 436661 247364 656062
rect 248060 648708 248112 648714
rect 248060 648650 248112 648656
rect 247414 613724 247470 613733
rect 247414 613659 247470 613668
rect 247322 436652 247378 436661
rect 247322 436587 247378 436596
rect 246310 316156 246366 316165
rect 246310 316091 246366 316100
rect 244846 278019 244853 278071
rect 244905 278019 244912 278071
rect 229844 266412 229896 266418
rect 229844 266354 229896 266360
rect 210432 259680 210484 259686
rect 210432 259622 210484 259628
rect 247428 259618 247456 613659
rect 248072 550085 248100 648650
rect 248058 550076 248114 550085
rect 248058 550011 248114 550020
rect 248164 396638 248192 674354
rect 248520 665232 248572 665238
rect 248520 665174 248572 665180
rect 248428 656188 248480 656194
rect 248428 656130 248480 656136
rect 248244 648504 248296 648510
rect 248244 648446 248296 648452
rect 248152 396632 248204 396638
rect 248152 396574 248204 396580
rect 248256 279474 248284 648446
rect 248336 648436 248388 648442
rect 248336 648378 248388 648384
rect 248244 279468 248296 279474
rect 248244 279410 248296 279416
rect 248152 279128 248204 279134
rect 248152 279070 248204 279076
rect 248164 278522 248192 279070
rect 248348 278590 248376 648378
rect 248440 280562 248468 656130
rect 248428 280556 248480 280562
rect 248428 280498 248480 280504
rect 248532 279134 248560 665174
rect 248992 493237 249020 700262
rect 250176 699436 250228 699442
rect 250176 699378 250228 699384
rect 249624 699164 249676 699170
rect 249624 699106 249676 699112
rect 249532 699096 249584 699102
rect 249532 699038 249584 699044
rect 249348 698960 249400 698966
rect 249348 698902 249400 698908
rect 249256 651700 249308 651706
rect 249256 651642 249308 651648
rect 249072 585536 249124 585542
rect 249072 585478 249124 585484
rect 248978 493228 249034 493237
rect 248978 493163 249034 493172
rect 248520 279128 248572 279134
rect 248520 279070 248572 279076
rect 249084 278998 249112 585478
rect 249164 583904 249216 583910
rect 249164 583846 249216 583852
rect 249176 280018 249204 583846
rect 249268 415445 249296 651642
rect 249254 415436 249310 415445
rect 249254 415371 249310 415380
rect 249360 358597 249388 698902
rect 249440 648640 249492 648646
rect 249440 648582 249492 648588
rect 249346 358588 249402 358597
rect 249346 358523 249402 358532
rect 249164 280012 249216 280018
rect 249164 279954 249216 279960
rect 249452 279678 249480 648582
rect 249440 279672 249492 279678
rect 249440 279614 249492 279620
rect 249072 278992 249124 278998
rect 249072 278934 249124 278940
rect 249544 278726 249572 699038
rect 249532 278720 249584 278726
rect 249532 278662 249584 278668
rect 248336 278584 248388 278590
rect 248336 278526 248388 278532
rect 248152 278516 248204 278522
rect 248152 278458 248204 278464
rect 249636 278454 249664 699106
rect 250084 652924 250136 652930
rect 250084 652866 250136 652872
rect 250096 585445 250124 652866
rect 250082 585436 250138 585445
rect 250082 585371 250138 585380
rect 250082 386876 250138 386885
rect 250082 386811 250138 386820
rect 250096 386302 250124 386811
rect 250084 386296 250136 386302
rect 250084 386238 250136 386244
rect 250188 284098 250216 699378
rect 250726 699132 250782 699141
rect 250726 699067 250782 699076
rect 250636 698892 250688 698898
rect 250636 698834 250688 698840
rect 250544 666728 250596 666734
rect 250544 666670 250596 666676
rect 250268 653944 250320 653950
rect 250268 653886 250320 653892
rect 250280 401029 250308 653886
rect 250360 651836 250412 651842
rect 250360 651778 250412 651784
rect 250266 401020 250322 401029
rect 250266 400955 250322 400964
rect 250372 365669 250400 651778
rect 250450 648404 250506 648413
rect 250450 648339 250506 648348
rect 250358 365660 250414 365669
rect 250358 365595 250414 365604
rect 250176 284092 250228 284098
rect 250176 284034 250228 284040
rect 250464 278794 250492 648339
rect 250556 280358 250584 666670
rect 250648 280494 250676 698834
rect 250636 280488 250688 280494
rect 250636 280430 250688 280436
rect 250544 280352 250596 280358
rect 250544 280294 250596 280300
rect 250740 280086 250768 699067
rect 250818 514444 250874 514453
rect 250818 514379 250874 514388
rect 250832 514346 250860 514379
rect 250820 514340 250872 514346
rect 250820 514282 250872 514288
rect 250818 479084 250874 479093
rect 250818 479019 250874 479028
rect 250832 478986 250860 479019
rect 250820 478980 250872 478986
rect 250820 478922 250872 478928
rect 250818 422508 250874 422517
rect 250818 422443 250874 422452
rect 250832 421594 250860 422443
rect 250820 421588 250872 421594
rect 250820 421530 250872 421536
rect 250728 280080 250780 280086
rect 250728 280022 250780 280028
rect 250452 278788 250504 278794
rect 250452 278730 250504 278736
rect 250924 278658 250952 728958
rect 287712 728472 287764 728478
rect 287712 728414 287764 728420
rect 257904 703720 257956 703726
rect 257904 703662 257956 703668
rect 255696 699572 255748 699578
rect 255696 699514 255748 699520
rect 251280 698756 251332 698762
rect 251280 698698 251332 698704
rect 251096 661152 251148 661158
rect 251096 661094 251148 661100
rect 251004 652992 251056 652998
rect 251004 652934 251056 652940
rect 251016 521525 251044 652934
rect 251002 521516 251058 521525
rect 251002 521451 251058 521460
rect 251108 464949 251136 661094
rect 251188 557860 251240 557866
rect 251188 557802 251240 557808
rect 251094 464940 251150 464949
rect 251094 464875 251150 464884
rect 251200 280426 251228 557802
rect 251292 393957 251320 698698
rect 251740 687672 251792 687678
rect 251740 687614 251792 687620
rect 251648 671080 251700 671086
rect 251648 671022 251700 671028
rect 251556 666796 251608 666802
rect 251556 666738 251608 666744
rect 251464 665572 251516 665578
rect 251464 665514 251516 665520
rect 251372 647280 251424 647286
rect 251372 647222 251424 647228
rect 251278 393948 251334 393957
rect 251278 393883 251334 393892
rect 251188 280420 251240 280426
rect 251188 280362 251240 280368
rect 251384 280290 251412 647222
rect 251372 280284 251424 280290
rect 251372 280226 251424 280232
rect 251476 279542 251504 665514
rect 251568 279610 251596 666738
rect 251556 279604 251608 279610
rect 251556 279546 251608 279552
rect 251464 279536 251516 279542
rect 251464 279478 251516 279484
rect 250912 278652 250964 278658
rect 250912 278594 250964 278600
rect 249624 278448 249676 278454
rect 249624 278390 249676 278396
rect 251660 278318 251688 671022
rect 251752 278862 251780 687614
rect 252844 667816 252896 667822
rect 252844 667758 252896 667764
rect 252752 666660 252804 666666
rect 252752 666602 252804 666608
rect 252016 666184 252068 666190
rect 252016 666126 252068 666132
rect 251832 651768 251884 651774
rect 251832 651710 251884 651716
rect 251844 627877 251872 651710
rect 251830 627868 251886 627877
rect 251830 627803 251886 627812
rect 252028 606661 252056 666126
rect 252660 662784 252712 662790
rect 252660 662726 252712 662732
rect 252292 649048 252344 649054
rect 252292 648990 252344 648996
rect 252108 647484 252160 647490
rect 252108 647426 252160 647432
rect 252014 606652 252070 606661
rect 252014 606587 252070 606596
rect 252014 535660 252070 535669
rect 252014 535595 252070 535604
rect 251922 337372 251978 337381
rect 251922 337307 251978 337316
rect 251936 279134 251964 337307
rect 251924 279128 251976 279134
rect 251924 279070 251976 279076
rect 251740 278856 251792 278862
rect 251740 278798 251792 278804
rect 251648 278312 251700 278318
rect 251648 278254 251700 278260
rect 252028 261998 252056 535595
rect 252120 429589 252148 647426
rect 252200 647416 252252 647422
rect 252200 647358 252252 647364
rect 252212 472021 252240 647358
rect 252304 486165 252332 648990
rect 252568 648572 252620 648578
rect 252568 648514 252620 648520
rect 252476 647892 252528 647898
rect 252476 647834 252528 647840
rect 252384 646872 252436 646878
rect 252384 646814 252436 646820
rect 252396 620805 252424 646814
rect 252382 620796 252438 620805
rect 252382 620731 252438 620740
rect 252382 606652 252438 606661
rect 252382 606587 252438 606596
rect 252396 605942 252424 606587
rect 252384 605936 252436 605942
rect 252384 605878 252436 605884
rect 252384 585468 252436 585474
rect 252384 585410 252436 585416
rect 252290 486156 252346 486165
rect 252290 486091 252346 486100
rect 252198 472012 252254 472021
rect 252198 471947 252254 471956
rect 252396 443733 252424 585410
rect 252488 507653 252516 647834
rect 252580 642293 252608 648514
rect 252566 642284 252622 642293
rect 252566 642219 252622 642228
rect 252474 507644 252530 507653
rect 252474 507579 252530 507588
rect 252382 443724 252438 443733
rect 252382 443659 252438 443668
rect 252106 429580 252162 429589
rect 252106 429515 252162 429524
rect 252200 396632 252252 396638
rect 252200 396574 252252 396580
rect 252106 351516 252162 351525
rect 252106 351451 252162 351460
rect 252120 280222 252148 351451
rect 252212 323237 252240 396574
rect 252672 344725 252700 662726
rect 252658 344716 252714 344725
rect 252658 344651 252714 344660
rect 252290 330300 252346 330309
rect 252290 330235 252346 330244
rect 252198 323228 252254 323237
rect 252198 323163 252254 323172
rect 252198 309084 252254 309093
rect 252198 309019 252254 309028
rect 252108 280216 252160 280222
rect 252108 280158 252160 280164
rect 252212 279066 252240 309019
rect 252304 280533 252332 330235
rect 252382 294940 252438 294949
rect 252382 294875 252438 294884
rect 252290 280524 252346 280533
rect 252290 280459 252346 280468
rect 252396 280154 252424 294875
rect 252384 280148 252436 280154
rect 252384 280090 252436 280096
rect 252764 279746 252792 666602
rect 252752 279740 252804 279746
rect 252752 279682 252804 279688
rect 252200 279060 252252 279066
rect 252200 279002 252252 279008
rect 252856 278386 252884 667758
rect 254406 646908 254462 646917
rect 255708 646878 255736 699514
rect 257916 646917 257944 703662
rect 287252 699504 287304 699510
rect 287252 699446 287304 699452
rect 286606 698860 286662 698869
rect 286606 698795 286662 698804
rect 279892 687672 279944 687678
rect 279892 687614 279944 687620
rect 279904 687445 279932 687614
rect 279890 687436 279946 687445
rect 279890 687371 279946 687380
rect 279982 681452 280038 681461
rect 279982 681387 280038 681396
rect 270232 667340 270284 667346
rect 270232 667282 270284 667288
rect 267840 667224 267892 667230
rect 270244 667210 270272 667282
rect 267840 667166 267892 667172
rect 270232 667204 270284 667210
rect 267852 665850 267880 667166
rect 270232 667146 270284 667152
rect 267840 665844 267892 665850
rect 267840 665786 267892 665792
rect 258548 654012 258600 654018
rect 258548 653954 258600 653960
rect 258560 646917 258588 653954
rect 279996 646917 280024 681387
rect 286422 671116 286478 671125
rect 286422 671051 286478 671060
rect 286436 671018 286464 671051
rect 286424 671012 286476 671018
rect 286424 670954 286476 670960
rect 286620 667822 286648 698795
rect 286608 667816 286660 667822
rect 286608 667758 286660 667764
rect 286884 667816 286936 667822
rect 286884 667758 286936 667764
rect 286896 667414 286924 667758
rect 286884 667408 286936 667414
rect 286884 667350 286936 667356
rect 282928 657208 282980 657214
rect 282928 657150 282980 657156
rect 282940 647030 282968 657150
rect 282940 647002 283336 647030
rect 287264 646917 287292 699446
rect 287724 692574 287752 728414
rect 335828 728336 335880 728342
rect 335828 728278 335880 728284
rect 320740 708004 320792 708010
rect 320740 707946 320792 707952
rect 314942 699948 314998 699957
rect 314942 699883 314998 699892
rect 288538 699812 288594 699821
rect 288538 699747 288594 699756
rect 288724 699776 288776 699782
rect 288262 695188 288318 695197
rect 288262 695123 288318 695132
rect 287712 692568 287764 692574
rect 287712 692510 287764 692516
rect 288170 679140 288226 679149
rect 288170 679075 288226 679084
rect 288078 676964 288134 676973
rect 288078 676899 288134 676908
rect 287986 674788 288042 674797
rect 287986 674723 288042 674732
rect 288000 674418 288028 674723
rect 287988 674412 288040 674418
rect 287988 674354 288040 674360
rect 287894 672884 287950 672893
rect 287894 672819 287950 672828
rect 287908 664898 287936 672819
rect 288000 665510 288028 674354
rect 287988 665504 288040 665510
rect 287988 665446 288040 665452
rect 288092 665102 288120 676899
rect 288184 666054 288212 679075
rect 288276 666394 288304 695123
rect 288446 693284 288502 693293
rect 288446 693219 288502 693228
rect 288264 666388 288316 666394
rect 288264 666330 288316 666336
rect 288460 666122 288488 693219
rect 288552 686221 288580 699747
rect 288724 699718 288776 699724
rect 288632 699300 288684 699306
rect 288632 699242 288684 699248
rect 288538 686212 288594 686221
rect 288538 686147 288594 686156
rect 288538 682948 288594 682957
rect 288538 682883 288594 682892
rect 288552 666258 288580 682883
rect 288644 682413 288672 699242
rect 288736 690573 288764 699718
rect 308136 699572 308188 699578
rect 308136 699514 308188 699520
rect 299856 699504 299908 699510
rect 299856 699446 299908 699452
rect 302616 699504 302668 699510
rect 302616 699446 302668 699452
rect 298382 699268 298438 699277
rect 289092 699232 289144 699238
rect 298382 699203 298438 699212
rect 289092 699174 289144 699180
rect 289104 698733 289132 699174
rect 292864 699164 292916 699170
rect 298396 699118 298424 699203
rect 299868 699118 299896 699446
rect 301144 699436 301196 699442
rect 301144 699378 301196 699384
rect 301156 699118 301184 699378
rect 301694 699268 301750 699277
rect 301694 699203 301750 699212
rect 292864 699106 292916 699112
rect 291482 698996 291538 699005
rect 292876 698982 292904 699106
rect 295544 699102 295664 699118
rect 297016 699102 297320 699118
rect 295544 699096 295676 699102
rect 295544 699090 295624 699096
rect 297016 699096 297332 699102
rect 297016 699090 297280 699096
rect 295624 699038 295676 699044
rect 298304 699090 298424 699118
rect 299776 699090 299896 699118
rect 301064 699090 301184 699118
rect 297280 699038 297332 699044
rect 292784 698954 292904 698982
rect 294980 699028 295032 699034
rect 294980 698970 295032 698976
rect 291482 698931 291538 698940
rect 290010 698860 290066 698869
rect 294992 698846 295020 698970
rect 301708 698898 301736 699203
rect 302628 699118 302656 699446
rect 303904 699436 303956 699442
rect 303904 699378 303956 699384
rect 303916 699118 303944 699378
rect 306846 699268 306902 699277
rect 306846 699203 306902 699212
rect 302536 699090 302656 699118
rect 303824 699090 303944 699118
rect 301788 699028 301840 699034
rect 305560 699028 305612 699034
rect 301788 698970 301840 698976
rect 305296 698976 305560 698982
rect 305296 698970 305612 698976
rect 301800 698898 301828 698970
rect 305296 698954 305600 698970
rect 306584 698966 306704 698982
rect 306584 698960 306716 698966
rect 306584 698954 306664 698960
rect 306664 698902 306716 698908
rect 306860 698898 306888 699203
rect 308148 699118 308176 699514
rect 309424 699368 309476 699374
rect 309424 699310 309476 699316
rect 309436 699118 309464 699310
rect 308056 699090 308176 699118
rect 309344 699090 309464 699118
rect 310802 699132 310858 699141
rect 310802 699067 310858 699076
rect 294256 698818 295020 698846
rect 301696 698892 301748 698898
rect 301696 698834 301748 698840
rect 301788 698892 301840 698898
rect 301788 698834 301840 698840
rect 306848 698892 306900 698898
rect 313656 698892 313708 698898
rect 306848 698834 306900 698840
rect 312090 698860 312146 698869
rect 290010 698795 290066 698804
rect 312090 698795 312146 698804
rect 313562 698860 313618 698869
rect 313618 698840 313656 698846
rect 314956 698846 314984 699883
rect 317704 699368 317756 699374
rect 317704 699310 317756 699316
rect 317716 699118 317744 699310
rect 317624 699090 317744 699118
rect 316336 698966 316640 698982
rect 316336 698960 316652 698966
rect 316336 698954 316600 698960
rect 316600 698902 316652 698908
rect 320648 698892 320700 698898
rect 313618 698834 313708 698840
rect 313618 698818 313696 698834
rect 314836 698818 314984 698846
rect 319082 698860 319138 698869
rect 313562 698795 313618 698804
rect 314836 698760 314864 698818
rect 320384 698840 320648 698846
rect 320384 698834 320700 698840
rect 320384 698818 320688 698834
rect 319082 698795 319138 698804
rect 314824 698754 314876 698760
rect 289090 698724 289146 698733
rect 314824 698696 314876 698702
rect 314836 698680 314864 698696
rect 289090 698659 289146 698668
rect 320646 696004 320702 696013
rect 320476 695962 320646 695990
rect 288814 691108 288870 691117
rect 288814 691043 288870 691052
rect 288722 690564 288778 690573
rect 288722 690499 288778 690508
rect 288630 682404 288686 682413
rect 288630 682339 288686 682348
rect 288644 681461 288672 682339
rect 288630 681452 288686 681461
rect 288630 681387 288686 681396
rect 288540 666252 288592 666258
rect 288540 666194 288592 666200
rect 288448 666116 288500 666122
rect 288448 666058 288500 666064
rect 288172 666048 288224 666054
rect 288172 665990 288224 665996
rect 288080 665096 288132 665102
rect 288080 665038 288132 665044
rect 287896 664892 287948 664898
rect 287896 664834 287948 664840
rect 288828 647354 288856 691043
rect 289090 668804 289146 668813
rect 289090 668739 289146 668748
rect 289104 664966 289132 668739
rect 290748 667340 290800 667346
rect 315496 667340 315548 667346
rect 290748 667282 290800 667288
rect 290838 667308 290894 667317
rect 289288 667130 289408 667158
rect 290576 667130 290696 667158
rect 289380 666802 289408 667130
rect 290668 666870 290696 667130
rect 290656 666864 290708 666870
rect 290656 666806 290708 666812
rect 289368 666796 289420 666802
rect 289366 666764 289368 666773
rect 289420 666764 289422 666773
rect 289366 666699 289422 666708
rect 289380 666673 289408 666699
rect 290668 666666 290696 666806
rect 290656 666660 290708 666666
rect 290656 666602 290708 666608
rect 290760 665918 290788 667282
rect 311354 667308 311410 667317
rect 303088 667278 303208 667294
rect 303088 667272 303220 667278
rect 303088 667266 303168 667272
rect 290838 667243 290894 667252
rect 290852 666326 290880 667243
rect 311354 667243 311410 667252
rect 311538 667308 311594 667317
rect 315496 667282 315548 667288
rect 316048 667340 316100 667346
rect 316048 667282 316100 667288
rect 311538 667243 311594 667252
rect 303168 667214 303220 667220
rect 301602 667172 301658 667181
rect 290840 666320 290892 666326
rect 290840 666262 290892 666268
rect 290748 665912 290800 665918
rect 290748 665854 290800 665860
rect 290852 665578 290880 666262
rect 290840 665572 290892 665578
rect 290840 665514 290892 665520
rect 292048 665034 292076 667158
rect 292036 665028 292088 665034
rect 292036 664970 292088 664976
rect 289092 664960 289144 664966
rect 289092 664902 289144 664908
rect 293336 662790 293364 667158
rect 294808 666462 294836 667158
rect 296096 667130 296216 667158
rect 296188 666734 296216 667130
rect 297568 666938 297596 667158
rect 297556 666932 297608 666938
rect 297556 666874 297608 666880
rect 298752 666796 298804 666802
rect 298752 666738 298804 666744
rect 296176 666728 296228 666734
rect 296176 666670 296228 666676
rect 294796 666456 294848 666462
rect 294796 666398 294848 666404
rect 298764 666326 298792 666738
rect 298752 666320 298804 666326
rect 298752 666262 298804 666268
rect 298856 665374 298884 667158
rect 297832 665368 297884 665374
rect 297832 665310 297884 665316
rect 298844 665368 298896 665374
rect 298844 665310 298896 665316
rect 293324 662784 293376 662790
rect 293324 662726 293376 662732
rect 288816 647348 288868 647354
rect 288816 647290 288868 647296
rect 288828 647150 288856 647290
rect 288816 647144 288868 647150
rect 288816 647086 288868 647092
rect 297556 647076 297608 647082
rect 297556 647018 297608 647024
rect 292772 646940 292824 646946
rect 257902 646908 257958 646917
rect 254406 646843 254462 646852
rect 255696 646872 255748 646878
rect 257902 646843 257958 646852
rect 258546 646908 258602 646917
rect 258546 646843 258602 646852
rect 259190 646908 259246 646917
rect 278510 646908 278566 646917
rect 259190 646843 259246 646852
rect 268680 646866 268984 646894
rect 273648 646866 273768 646894
rect 255696 646814 255748 646820
rect 268680 646810 268708 646866
rect 273648 646810 273676 646866
rect 278510 646843 278566 646852
rect 279982 646908 280038 646917
rect 279982 646843 280038 646852
rect 287250 646908 287306 646917
rect 287250 646843 287306 646852
rect 288078 646908 288134 646917
rect 297568 646894 297596 647018
rect 292824 646888 292904 646894
rect 292772 646882 292904 646888
rect 292784 646866 292904 646882
rect 297568 646866 297688 646894
rect 288078 646843 288134 646852
rect 297844 646810 297872 665310
rect 300328 663878 300356 667158
rect 308226 667172 308282 667181
rect 301602 667107 301658 667116
rect 304376 665102 304404 667158
rect 305848 665374 305876 667158
rect 307136 666909 307164 667158
rect 308226 667107 308228 667116
rect 308280 667107 308282 667116
rect 308594 667172 308650 667181
rect 309896 667130 310200 667158
rect 308594 667107 308650 667116
rect 308228 667078 308280 667084
rect 307122 666900 307178 666909
rect 307122 666835 307178 666844
rect 306480 666252 306532 666258
rect 306480 666194 306532 666200
rect 304916 665368 304968 665374
rect 304916 665310 304968 665316
rect 305836 665368 305888 665374
rect 305836 665310 305888 665316
rect 301604 665096 301656 665102
rect 301604 665038 301656 665044
rect 304364 665096 304416 665102
rect 304364 665038 304416 665044
rect 300316 663872 300368 663878
rect 300316 663814 300368 663820
rect 301616 646917 301644 665038
rect 304928 648714 304956 665310
rect 306492 663946 306520 666194
rect 306480 663940 306532 663946
rect 306480 663882 306532 663888
rect 307124 658364 307176 658370
rect 307124 658306 307176 658312
rect 304916 648708 304968 648714
rect 304916 648650 304968 648656
rect 307136 647030 307164 658306
rect 308240 647082 308268 667078
rect 310172 667074 310200 667130
rect 310160 667068 310212 667074
rect 310160 667010 310212 667016
rect 311552 648549 311580 667243
rect 315508 667158 315536 667282
rect 312656 656126 312684 667158
rect 314128 666530 314156 667158
rect 315416 667130 315536 667158
rect 314116 666524 314168 666530
rect 314116 666466 314168 666472
rect 312644 656120 312696 656126
rect 312644 656062 312696 656068
rect 315956 656120 316008 656126
rect 315956 656062 316008 656068
rect 311538 648540 311594 648549
rect 311538 648475 311594 648484
rect 308228 647076 308280 647082
rect 307136 647002 307256 647030
rect 308228 647018 308280 647024
rect 315968 646917 315996 656062
rect 316060 648646 316088 667282
rect 316888 666598 316916 667158
rect 318176 667006 318204 667158
rect 319648 667130 319768 667158
rect 318164 667000 318216 667006
rect 318164 666942 318216 666948
rect 316876 666592 316928 666598
rect 316876 666534 316928 666540
rect 319740 664830 319768 667130
rect 319728 664824 319780 664830
rect 319728 664766 319780 664772
rect 316048 648640 316100 648646
rect 316048 648582 316100 648588
rect 319740 648578 319768 664766
rect 319728 648572 319780 648578
rect 319728 648514 319780 648520
rect 320476 647082 320504 695962
rect 320646 695939 320702 695948
rect 320556 695832 320608 695838
rect 320556 695774 320608 695780
rect 320568 691366 320596 695774
rect 320648 695152 320700 695158
rect 320648 695094 320700 695100
rect 320660 691486 320688 695094
rect 320648 691480 320700 691486
rect 320648 691422 320700 691428
rect 320646 691380 320702 691389
rect 320568 691338 320646 691366
rect 320646 691315 320702 691324
rect 320646 686348 320702 686357
rect 320568 686306 320646 686334
rect 320568 647218 320596 686306
rect 320646 686283 320702 686292
rect 320646 684172 320702 684181
rect 320646 684107 320702 684116
rect 320660 647490 320688 684107
rect 320752 676973 320780 707946
rect 323040 701408 323092 701414
rect 323040 701350 323092 701356
rect 322578 700084 322634 700093
rect 322578 700019 322634 700028
rect 321108 699844 321160 699850
rect 321108 699786 321160 699792
rect 321014 698996 321070 699005
rect 321014 698931 321070 698940
rect 321028 694546 321056 698931
rect 321016 694540 321068 694546
rect 321016 694482 321068 694488
rect 320830 694236 320886 694245
rect 321120 694234 321148 699786
rect 321568 699436 321620 699442
rect 321568 699378 321620 699384
rect 321200 698756 321252 698762
rect 321200 698698 321252 698704
rect 321212 695838 321240 698698
rect 321580 698082 321608 699378
rect 321844 699164 321896 699170
rect 321844 699106 321896 699112
rect 321568 698076 321620 698082
rect 321568 698018 321620 698024
rect 321200 695832 321252 695838
rect 321200 695774 321252 695780
rect 321856 694614 321884 699106
rect 322028 699096 322080 699102
rect 322028 699038 322080 699044
rect 321936 694812 321988 694818
rect 321936 694754 321988 694760
rect 321844 694608 321896 694614
rect 321844 694550 321896 694556
rect 320830 694171 320886 694180
rect 321028 694206 321148 694234
rect 320738 676964 320794 676973
rect 320738 676899 320794 676908
rect 320738 673700 320794 673709
rect 320738 673635 320794 673644
rect 320752 665442 320780 673635
rect 320740 665436 320792 665442
rect 320740 665378 320792 665384
rect 320844 665374 320872 694171
rect 320922 691924 320978 691933
rect 320922 691859 320978 691868
rect 320936 665850 320964 691859
rect 321028 681053 321056 694206
rect 321108 691480 321160 691486
rect 321108 691422 321160 691428
rect 321120 684181 321148 691422
rect 321106 684172 321162 684181
rect 321106 684107 321162 684116
rect 321014 681044 321070 681053
rect 321014 680979 321070 680988
rect 321028 678778 321056 680979
rect 321028 678750 321148 678778
rect 321014 669620 321070 669629
rect 321014 669555 321070 669564
rect 321028 666666 321056 669555
rect 321016 666660 321068 666666
rect 321016 666602 321068 666608
rect 320924 665844 320976 665850
rect 320924 665786 320976 665792
rect 320832 665368 320884 665374
rect 320832 665310 320884 665316
rect 320648 647484 320700 647490
rect 320648 647426 320700 647432
rect 321028 647422 321056 666602
rect 321120 648510 321148 678750
rect 321198 677780 321254 677789
rect 321198 677715 321254 677724
rect 321212 665918 321240 677715
rect 321290 671660 321346 671669
rect 321290 671595 321346 671604
rect 321304 666326 321332 671595
rect 321948 667142 321976 694754
rect 322040 684346 322068 699038
rect 322592 695158 322620 700019
rect 322580 695152 322632 695158
rect 322580 695094 322632 695100
rect 322028 684340 322080 684346
rect 322028 684282 322080 684288
rect 321936 667136 321988 667142
rect 321936 667078 321988 667084
rect 321292 666320 321344 666326
rect 321292 666262 321344 666268
rect 321200 665912 321252 665918
rect 321200 665854 321252 665860
rect 321476 664892 321528 664898
rect 321476 664834 321528 664840
rect 321108 648504 321160 648510
rect 321108 648446 321160 648452
rect 321016 647416 321068 647422
rect 321016 647358 321068 647364
rect 320556 647212 320608 647218
rect 320556 647154 320608 647160
rect 320464 647076 320516 647082
rect 320464 647018 320516 647024
rect 321488 647030 321516 664834
rect 321488 647002 321608 647030
rect 323052 646946 323080 701350
rect 329664 699504 329716 699510
rect 329664 699446 329716 699452
rect 324788 699368 324840 699374
rect 324788 699310 324840 699316
rect 323682 698860 323738 698869
rect 323682 698795 323738 698804
rect 323696 698150 323724 698795
rect 323684 698144 323736 698150
rect 323684 698086 323736 698092
rect 324800 693186 324828 699310
rect 328560 699028 328612 699034
rect 328560 698970 328612 698976
rect 324788 693180 324840 693186
rect 324788 693122 324840 693128
rect 324800 648442 324828 693122
rect 328572 678838 328600 698970
rect 328560 678832 328612 678838
rect 328560 678774 328612 678780
rect 329676 673330 329704 699446
rect 330768 699300 330820 699306
rect 330768 699242 330820 699248
rect 330780 682170 330808 699242
rect 330768 682164 330820 682170
rect 330768 682106 330820 682112
rect 329664 673324 329716 673330
rect 329664 673266 329716 673272
rect 335552 667612 335604 667618
rect 335552 667554 335604 667560
rect 325246 667444 325302 667453
rect 325246 667379 325302 667388
rect 325260 666637 325288 667379
rect 325246 666628 325302 666637
rect 325246 666563 325302 666572
rect 335564 666394 335592 667554
rect 335644 666932 335696 666938
rect 335644 666874 335696 666880
rect 335656 666394 335684 666874
rect 335552 666388 335604 666394
rect 335552 666330 335604 666336
rect 335644 666388 335696 666394
rect 335644 666330 335696 666336
rect 324788 648436 324840 648442
rect 324788 648378 324840 648384
rect 335840 647030 335868 728278
rect 351296 705834 351324 729514
rect 351388 729486 351600 729514
rect 351388 714674 351416 729486
rect 351572 729446 351600 729486
rect 351693 729446 351721 729514
rect 351838 729446 351866 729514
rect 351572 729430 351866 729446
rect 351572 729424 351878 729430
rect 351572 729418 351826 729424
rect 351826 729366 351878 729372
rect 351838 729335 351866 729366
rect 353163 729310 353191 729514
rect 353872 729430 353900 729514
rect 355071 729484 355123 729552
rect 354608 729456 355123 729484
rect 353860 729424 353912 729430
rect 353860 729366 353912 729372
rect 353136 729294 353191 729310
rect 352388 729288 352440 729294
rect 352388 729230 352440 729236
rect 353136 729288 353203 729294
rect 353136 729236 353151 729288
rect 353136 729230 353203 729236
rect 351376 714668 351428 714674
rect 351376 714610 351428 714616
rect 351284 705828 351336 705834
rect 351284 705770 351336 705776
rect 344660 704740 344712 704746
rect 344660 704682 344712 704688
rect 341072 670468 341124 670474
rect 341072 670410 341124 670416
rect 341084 667482 341112 670410
rect 341484 670342 341808 670368
rect 341484 669822 341500 670342
rect 341796 669822 341808 670342
rect 341484 667906 341808 669822
rect 343144 670294 343468 670332
rect 343144 669782 343162 670294
rect 343450 669782 343468 670294
rect 341480 667890 342848 667906
rect 341480 667818 341506 667890
rect 342830 667818 342848 667890
rect 341480 667800 342848 667818
rect 342544 667544 342596 667550
rect 342544 667486 342596 667492
rect 341072 667476 341124 667482
rect 341072 667418 341124 667424
rect 337300 667408 337352 667414
rect 337300 667350 337352 667356
rect 338956 667408 339008 667414
rect 338956 667350 339008 667356
rect 337312 667278 337340 667350
rect 337300 667272 337352 667278
rect 337300 667214 337352 667220
rect 338968 665170 338996 667350
rect 342556 667346 342584 667486
rect 342544 667340 342596 667346
rect 342544 667282 342596 667288
rect 342740 667266 342952 667294
rect 340970 667170 342572 667204
rect 340970 667088 340998 667170
rect 342546 667088 342572 667170
rect 340970 667070 342572 667088
rect 342140 666736 342464 667070
rect 342740 667006 342768 667266
rect 342924 667142 342952 667266
rect 342912 667136 342964 667142
rect 342912 667078 342964 667084
rect 342728 667000 342780 667006
rect 342728 666942 342780 666948
rect 342912 667000 342964 667006
rect 342912 666942 342964 666948
rect 342820 666932 342872 666938
rect 342924 666886 342952 666942
rect 342872 666880 342952 666886
rect 342820 666874 342952 666880
rect 342832 666858 342952 666874
rect 343144 666736 343468 669782
rect 344108 666932 344160 666938
rect 344108 666874 344160 666880
rect 342140 666412 343468 666736
rect 344120 666394 344148 666874
rect 344108 666388 344160 666394
rect 344108 666330 344160 666336
rect 338956 665164 339008 665170
rect 338956 665106 339008 665112
rect 335840 647002 335960 647030
rect 323040 646940 323092 646946
rect 301602 646908 301658 646917
rect 301602 646843 301658 646852
rect 302430 646908 302486 646917
rect 315954 646908 316010 646917
rect 302430 646843 302486 646852
rect 311920 646866 312040 646894
rect 311920 646810 311948 646866
rect 315954 646843 316010 646852
rect 316782 646908 316838 646917
rect 323040 646882 323092 646888
rect 326260 646940 326312 646946
rect 344672 646917 344700 704682
rect 352400 670474 352428 729230
rect 353136 728750 353164 729230
rect 353124 728744 353176 728750
rect 353124 728686 353176 728692
rect 354608 703726 354636 729456
rect 355071 729455 355123 729456
rect 355932 729430 355960 729514
rect 355920 729424 355972 729430
rect 355920 729366 355972 729372
rect 356310 729310 356338 729514
rect 356762 729430 356790 729514
rect 356975 729446 357003 729514
rect 357644 729486 357718 729514
rect 358196 729486 358316 729514
rect 359649 729494 359701 729552
rect 356750 729424 356802 729430
rect 356975 729418 357028 729446
rect 356750 729366 356802 729372
rect 356762 729333 356790 729366
rect 356748 729324 356804 729333
rect 356310 729282 356384 729310
rect 356356 728886 356384 729282
rect 356748 729259 356804 729268
rect 356344 728880 356396 728886
rect 356344 728822 356396 728828
rect 357000 728682 357028 729418
rect 357644 728750 357672 729486
rect 358196 728818 358224 729486
rect 359649 729466 359788 729494
rect 358184 728812 358236 728818
rect 358184 728754 358236 728760
rect 357632 728744 357684 728750
rect 357632 728686 357684 728692
rect 356988 728676 357040 728682
rect 356988 728618 357040 728624
rect 359760 719094 359788 729466
rect 360572 729464 360622 729551
rect 360572 729436 360984 729464
rect 360956 728954 360984 729436
rect 361036 729424 361088 729430
rect 361036 729366 361088 729372
rect 361048 729333 361076 729366
rect 361034 729324 361090 729333
rect 361034 729259 361090 729268
rect 360944 728948 360996 728954
rect 360944 728890 360996 728896
rect 363992 728886 364020 729514
rect 366134 729430 366162 729514
rect 366476 729486 366577 729514
rect 378484 729486 378832 729514
rect 366122 729424 366174 729430
rect 366122 729366 366174 729372
rect 366134 729310 366162 729366
rect 366108 729282 366162 729310
rect 365634 728916 365690 728925
rect 363428 728880 363480 728886
rect 363428 728822 363480 728828
rect 363980 728880 364032 728886
rect 366108 728886 366136 729282
rect 365634 728851 365690 728860
rect 366096 728880 366148 728886
rect 363980 728822 364032 728828
rect 363440 719094 363468 728822
rect 359012 719088 359064 719094
rect 359012 719030 359064 719036
rect 359748 719088 359800 719094
rect 359748 719030 359800 719036
rect 363428 719088 363480 719094
rect 363428 719030 363480 719036
rect 354596 703720 354648 703726
rect 354596 703662 354648 703668
rect 354688 703584 354740 703590
rect 354688 703526 354740 703532
rect 352388 670468 352440 670474
rect 352388 670410 352440 670416
rect 354700 647030 354728 703526
rect 358736 699844 358788 699850
rect 358736 699786 358788 699792
rect 358748 694682 358776 699786
rect 358736 694676 358788 694682
rect 358736 694618 358788 694624
rect 356986 693556 357042 693565
rect 356986 693491 357042 693500
rect 357000 693186 357028 693491
rect 356988 693180 357040 693186
rect 356988 693122 357040 693128
rect 359024 660546 359052 719030
rect 365648 711342 365676 728851
rect 366096 728822 366148 728828
rect 366476 728818 366504 729486
rect 367658 729052 367714 729061
rect 367658 728987 367714 728996
rect 366464 728812 366516 728818
rect 366464 728754 366516 728760
rect 367672 727866 367700 728987
rect 368026 728916 368082 728925
rect 368026 728851 368082 728860
rect 368040 728614 368068 728851
rect 368028 728608 368080 728614
rect 368028 728550 368080 728556
rect 378804 727934 378832 729486
rect 378896 729446 378924 729514
rect 379034 729446 379062 729514
rect 378896 729430 379062 729446
rect 378896 729424 379074 729430
rect 378896 729418 379022 729424
rect 378896 728886 378924 729418
rect 379022 729366 379074 729372
rect 379034 729335 379062 729366
rect 380368 729362 380396 729514
rect 381074 729430 381102 729514
rect 381062 729424 381114 729430
rect 381062 729366 381114 729372
rect 380356 729356 380408 729362
rect 380356 729298 380408 729304
rect 382283 729310 382311 729514
rect 383132 729430 383160 729514
rect 383496 729446 383524 729514
rect 383120 729424 383172 729430
rect 383120 729366 383172 729372
rect 383404 729418 383524 729446
rect 383962 729430 383990 729514
rect 384048 729486 384203 729514
rect 384876 729486 384932 729514
rect 383950 729424 384002 729430
rect 378884 728880 378936 728886
rect 378884 728822 378936 728828
rect 380368 728750 380396 729298
rect 382283 729282 382328 729310
rect 380356 728744 380408 728750
rect 380356 728686 380408 728692
rect 378792 727928 378844 727934
rect 378792 727870 378844 727876
rect 367660 727860 367712 727866
rect 367660 727802 367712 727808
rect 382300 726778 382328 729282
rect 383404 728478 383432 729418
rect 383950 729366 384002 729372
rect 384048 728682 384076 729486
rect 384876 729362 384904 729486
rect 385490 729476 385548 729504
rect 386849 729494 386901 729552
rect 384864 729356 384916 729362
rect 384864 729298 384916 729304
rect 384876 728750 384904 729298
rect 385520 728818 385548 729476
rect 386624 729466 386901 729494
rect 387771 729494 387823 729554
rect 387771 729466 388124 729494
rect 385508 728812 385560 728818
rect 385508 728754 385560 728760
rect 384864 728744 384916 728750
rect 384864 728686 384916 728692
rect 384036 728676 384088 728682
rect 384036 728618 384088 728624
rect 383392 728472 383444 728478
rect 383392 728414 383444 728420
rect 382288 726772 382340 726778
rect 382288 726714 382340 726720
rect 365636 711336 365688 711342
rect 365636 711278 365688 711284
rect 383404 701414 383432 728414
rect 383392 701408 383444 701414
rect 383392 701350 383444 701356
rect 386624 700326 386652 729466
rect 386978 729426 387034 729435
rect 386978 729361 387034 729370
rect 388096 728002 388124 729466
rect 391178 729310 391206 729514
rect 393340 729430 393368 729514
rect 393616 729486 393777 729514
rect 405392 729486 405512 729514
rect 393328 729424 393380 729430
rect 393328 729366 393380 729372
rect 391132 729282 391206 729310
rect 391132 728478 391160 729282
rect 392222 729052 392278 729061
rect 392222 728987 392278 728996
rect 392236 728614 392264 728987
rect 393340 728886 393368 729366
rect 393328 728880 393380 728886
rect 393328 728822 393380 728828
rect 393616 728818 393644 729486
rect 394522 729052 394578 729061
rect 394522 728987 394578 728996
rect 393604 728812 393656 728818
rect 393604 728754 393656 728760
rect 392224 728608 392276 728614
rect 392224 728550 392276 728556
rect 391120 728472 391172 728478
rect 391120 728414 391172 728420
rect 394536 728070 394564 728987
rect 394524 728064 394576 728070
rect 394524 728006 394576 728012
rect 388084 727996 388136 728002
rect 388084 727938 388136 727944
rect 386612 700320 386664 700326
rect 386612 700262 386664 700268
rect 379066 700084 379122 700093
rect 379066 700019 379122 700028
rect 361772 699232 361824 699238
rect 361772 699174 361824 699180
rect 361680 698892 361732 698898
rect 361680 698834 361732 698840
rect 360666 684988 360722 684997
rect 360666 684923 360722 684932
rect 360680 684346 360708 684923
rect 360668 684340 360720 684346
rect 360668 684282 360720 684288
rect 359840 682164 359892 682170
rect 359840 682106 359892 682112
rect 359852 682005 359880 682106
rect 359838 681996 359894 682005
rect 359838 681931 359894 681940
rect 360758 673564 360814 673573
rect 360758 673499 360814 673508
rect 360772 673330 360800 673499
rect 360760 673324 360812 673330
rect 360760 673266 360812 673272
rect 360484 667272 360536 667278
rect 360484 667214 360536 667220
rect 360496 666938 360524 667214
rect 361128 667204 361180 667210
rect 361128 667146 361180 667152
rect 361140 667045 361168 667146
rect 361220 667068 361272 667074
rect 361126 667036 361182 667045
rect 361310 667036 361366 667045
rect 361272 667016 361310 667022
rect 361220 667010 361310 667016
rect 361232 666994 361310 667010
rect 361126 666971 361182 666980
rect 361310 666971 361366 666980
rect 360484 666932 360536 666938
rect 360484 666874 360536 666880
rect 359012 660540 359064 660546
rect 359012 660482 359064 660488
rect 361140 652794 361168 666971
rect 361692 666938 361720 698834
rect 361784 667142 361812 699174
rect 367106 698724 367162 698733
rect 367106 698659 367162 698668
rect 361864 694744 361916 694750
rect 367120 694738 367148 698659
rect 370788 694812 370840 694818
rect 370788 694754 370840 694760
rect 361864 694686 361916 694692
rect 361876 667210 361904 694686
rect 370800 694653 370828 694754
rect 376688 694750 377084 694766
rect 376676 694744 377084 694750
rect 376728 694738 377084 694744
rect 379080 694738 379108 700019
rect 385138 699948 385194 699957
rect 385138 699883 385194 699892
rect 381090 699812 381146 699821
rect 381090 699747 381146 699756
rect 384956 699776 385008 699782
rect 381104 694902 381132 699747
rect 384956 699718 385008 699724
rect 384968 695362 384996 699718
rect 384956 695356 385008 695362
rect 384956 695298 385008 695304
rect 381104 694874 381316 694902
rect 381104 694738 381132 694874
rect 376676 694686 376728 694692
rect 381288 694682 381316 694874
rect 385152 694738 385180 699883
rect 390016 698144 390068 698150
rect 390016 698086 390068 698092
rect 387164 695356 387216 695362
rect 387164 695298 387216 695304
rect 387176 694738 387204 695298
rect 372812 694676 372864 694682
rect 370786 694644 370842 694653
rect 370786 694579 370842 694588
rect 371154 694644 371210 694653
rect 381276 694676 381328 694682
rect 375018 694644 375074 694653
rect 372864 694624 373220 694630
rect 372812 694618 373220 694624
rect 372824 694602 373220 694618
rect 371154 694579 371210 694588
rect 375018 694579 375074 694588
rect 375202 694644 375258 694653
rect 381276 694618 381328 694624
rect 388832 694614 389228 694630
rect 375202 694579 375258 694588
rect 388820 694608 389228 694614
rect 375216 694546 375244 694579
rect 388872 694602 389228 694608
rect 388820 694550 388872 694556
rect 375204 694540 375256 694546
rect 365082 694508 365138 694517
rect 375204 694482 375256 694488
rect 383114 694508 383170 694517
rect 365082 694443 365138 694452
rect 383114 694443 383170 694452
rect 390028 690922 390056 698086
rect 390028 690894 390424 690922
rect 362874 690564 362930 690573
rect 362874 690499 362930 690508
rect 362414 687572 362470 687581
rect 362414 687507 362470 687516
rect 362322 675604 362378 675613
rect 362322 675539 362378 675548
rect 362336 667346 362364 675539
rect 362324 667340 362376 667346
rect 362324 667282 362376 667288
rect 362428 667278 362456 687507
rect 362506 684988 362562 684997
rect 362506 684923 362562 684932
rect 362416 667272 362468 667278
rect 362416 667214 362468 667220
rect 361864 667204 361916 667210
rect 361864 667146 361916 667152
rect 361772 667136 361824 667142
rect 361772 667078 361824 667084
rect 361680 666932 361732 666938
rect 361680 666874 361732 666880
rect 362428 662790 362456 667214
rect 362520 666190 362548 684923
rect 362598 679004 362654 679013
rect 362598 678939 362654 678948
rect 362612 678838 362640 678939
rect 362600 678832 362652 678838
rect 362600 678774 362652 678780
rect 362508 666184 362560 666190
rect 362508 666126 362560 666132
rect 362612 665170 362640 678774
rect 362690 673564 362746 673573
rect 362690 673499 362746 673508
rect 362704 667210 362732 673499
rect 362692 667204 362744 667210
rect 362692 667146 362744 667152
rect 362888 665238 362916 690499
rect 390290 689204 390346 689213
rect 390290 689139 390346 689148
rect 390304 683194 390332 689139
rect 390396 687173 390424 690894
rect 390382 687164 390438 687173
rect 390382 687099 390438 687108
rect 389936 683166 390332 683194
rect 382932 667340 382984 667346
rect 382984 667288 383340 667294
rect 382932 667282 383340 667288
rect 382944 667266 383340 667282
rect 363888 667204 363940 667210
rect 363256 666326 363284 667158
rect 381090 667172 381146 667181
rect 363888 667146 363940 667152
rect 363244 666320 363296 666326
rect 363244 666262 363296 666268
rect 362876 665232 362928 665238
rect 362876 665174 362928 665180
rect 362600 665164 362652 665170
rect 362600 665106 362652 665112
rect 362416 662784 362468 662790
rect 362416 662726 362468 662732
rect 361128 652788 361180 652794
rect 361128 652730 361180 652736
rect 363900 647422 363928 667146
rect 365096 666666 365124 667158
rect 365084 666660 365136 666666
rect 365084 666602 365136 666608
rect 365266 664996 365322 665005
rect 365266 664931 365322 664940
rect 363888 647416 363940 647422
rect 363888 647358 363940 647364
rect 365280 647354 365308 664931
rect 367120 664830 367148 667158
rect 369144 666938 369172 667158
rect 368856 666932 368908 666938
rect 368856 666874 368908 666880
rect 369132 666932 369184 666938
rect 369132 666874 369184 666880
rect 367108 664824 367160 664830
rect 367108 664766 367160 664772
rect 368868 652862 368896 666874
rect 371168 666462 371196 667158
rect 373192 666802 373220 667158
rect 375216 667006 375244 667158
rect 375204 667000 375256 667006
rect 375204 666942 375256 666948
rect 373180 666796 373232 666802
rect 373180 666738 373232 666744
rect 370512 666456 370564 666462
rect 370512 666398 370564 666404
rect 371156 666456 371208 666462
rect 371156 666398 371208 666404
rect 368856 652856 368908 652862
rect 368856 652798 368908 652804
rect 370524 650618 370552 666398
rect 375216 666258 375244 666942
rect 377136 666796 377188 666802
rect 377136 666738 377188 666744
rect 375204 666252 375256 666258
rect 375204 666194 375256 666200
rect 377148 665374 377176 666738
rect 377240 666734 377268 667158
rect 379264 666802 379292 667158
rect 381090 667107 381092 667116
rect 381144 667107 381146 667116
rect 381274 667172 381330 667181
rect 381274 667107 381330 667116
rect 381092 667078 381144 667084
rect 379252 666796 379304 666802
rect 379252 666738 379304 666744
rect 377228 666728 377280 666734
rect 377228 666670 377280 666676
rect 377136 665368 377188 665374
rect 377136 665310 377188 665316
rect 378884 665232 378936 665238
rect 378884 665174 378936 665180
rect 370512 650612 370564 650618
rect 370512 650554 370564 650560
rect 374284 648028 374336 648034
rect 374284 647970 374336 647976
rect 365268 647348 365320 647354
rect 365268 647290 365320 647296
rect 374296 647030 374324 647970
rect 378896 647030 378924 665174
rect 381104 647490 381132 667078
rect 385336 666666 385364 667158
rect 389384 666734 389412 667158
rect 389372 666728 389424 666734
rect 389372 666670 389424 666676
rect 385324 666660 385376 666666
rect 385324 666602 385376 666608
rect 385336 666501 385364 666602
rect 385322 666492 385378 666501
rect 385322 666427 385378 666436
rect 389384 665442 389412 666670
rect 389372 665436 389424 665442
rect 389372 665378 389424 665384
rect 389936 650686 389964 683166
rect 390290 680228 390346 680237
rect 390290 680163 390346 680172
rect 390200 676656 390252 676662
rect 390200 676598 390252 676604
rect 390212 676406 390240 676598
rect 390028 676378 390240 676406
rect 390028 650754 390056 676378
rect 390200 676316 390252 676322
rect 390200 676258 390252 676264
rect 390212 676134 390240 676258
rect 390120 676106 390240 676134
rect 390120 667210 390148 676106
rect 390304 675466 390332 680163
rect 390396 676322 390424 687099
rect 390658 677780 390714 677789
rect 390658 677715 390714 677724
rect 390672 676662 390700 677715
rect 390660 676656 390712 676662
rect 390660 676598 390712 676604
rect 390384 676316 390436 676322
rect 390384 676258 390436 676264
rect 390212 675438 390332 675466
rect 390212 667317 390240 675438
rect 390290 674244 390346 674253
rect 390290 674179 390346 674188
rect 390198 667308 390254 667317
rect 390198 667243 390254 667252
rect 390108 667204 390160 667210
rect 390108 667146 390160 667152
rect 390304 665510 390332 674179
rect 390474 671524 390530 671533
rect 390474 671459 390530 671468
rect 390382 668940 390438 668949
rect 390382 668875 390438 668884
rect 390396 666909 390424 668875
rect 390382 666900 390438 666909
rect 390488 666870 390516 671459
rect 390382 666835 390438 666844
rect 390476 666864 390528 666870
rect 390292 665504 390344 665510
rect 390292 665446 390344 665452
rect 390016 650748 390068 650754
rect 390016 650690 390068 650696
rect 389924 650680 389976 650686
rect 389924 650622 389976 650628
rect 381092 647484 381144 647490
rect 381092 647426 381144 647432
rect 388636 647484 388688 647490
rect 388636 647426 388688 647432
rect 383852 647348 383904 647354
rect 383852 647290 383904 647296
rect 383864 647030 383892 647290
rect 388648 647030 388676 647426
rect 390396 647354 390424 666835
rect 390476 666806 390528 666812
rect 402068 659452 402120 659458
rect 402068 659394 402120 659400
rect 390384 647348 390436 647354
rect 390384 647290 390436 647296
rect 393420 647076 393472 647082
rect 354700 647002 355096 647030
rect 374296 647002 374416 647030
rect 378896 647002 379200 647030
rect 383864 647002 383984 647030
rect 388648 647002 388768 647030
rect 393420 647018 393472 647024
rect 398204 647076 398256 647082
rect 398204 647018 398256 647024
rect 344658 646908 344714 646917
rect 326312 646888 326392 646894
rect 326260 646882 326392 646888
rect 326272 646866 326392 646882
rect 316782 646843 316838 646852
rect 344658 646843 344714 646852
rect 345486 646908 345542 646917
rect 393432 646894 393460 647018
rect 398216 646894 398244 647018
rect 402080 646917 402108 659394
rect 405392 647490 405420 729486
rect 405884 729484 405930 729546
rect 406026 729484 406078 729552
rect 407351 729494 407403 729552
rect 405760 729456 406432 729484
rect 405760 728886 405788 729456
rect 406026 729454 406078 729456
rect 406392 729430 406432 729456
rect 407048 729466 407403 729494
rect 406392 729424 406444 729430
rect 406392 729366 406444 729372
rect 405748 728880 405800 728886
rect 405748 728822 405800 728828
rect 407048 728750 407076 729466
rect 408060 729430 408088 729514
rect 408048 729424 408100 729430
rect 408048 729366 408100 729372
rect 409283 729310 409311 729514
rect 410130 729430 410158 729514
rect 410510 729486 410756 729514
rect 410118 729424 410170 729430
rect 410118 729366 410170 729372
rect 410130 729333 410158 729366
rect 409256 729282 409311 729310
rect 410116 729324 410172 729333
rect 407036 728744 407088 728750
rect 407036 728686 407088 728692
rect 409256 728138 409284 729282
rect 410116 729259 410172 729268
rect 410728 728478 410756 729486
rect 410962 729333 410990 729514
rect 410948 729324 411004 729333
rect 410948 729259 411004 729268
rect 411188 728682 411216 729514
rect 411904 729446 411932 729514
rect 411904 729418 411952 729446
rect 411924 728750 411952 729418
rect 412476 728818 412504 729514
rect 413849 729484 413901 729552
rect 414771 729494 414823 729552
rect 413120 729456 413901 729484
rect 412464 728812 412516 728818
rect 412464 728754 412516 728760
rect 411912 728744 411964 728750
rect 411912 728686 411964 728692
rect 411176 728676 411228 728682
rect 411176 728618 411228 728624
rect 410716 728472 410768 728478
rect 410716 728414 410768 728420
rect 409244 728132 409296 728138
rect 409244 728074 409296 728080
rect 413120 654018 413148 729456
rect 413849 729455 413901 729456
rect 414684 729466 414823 729494
rect 414304 729424 414356 729430
rect 414304 729366 414356 729372
rect 414316 729333 414344 729366
rect 414302 729324 414358 729333
rect 414302 729259 414358 729268
rect 414684 728206 414712 729466
rect 418180 728478 418208 729514
rect 420296 729486 420362 729514
rect 420190 729460 420246 729469
rect 420296 729430 420324 729486
rect 420190 729395 420246 729404
rect 420284 729424 420336 729430
rect 419914 729324 419970 729333
rect 419914 729259 419970 729268
rect 417524 728472 417576 728478
rect 417524 728414 417576 728420
rect 418168 728472 418220 728478
rect 418168 728414 418220 728420
rect 414672 728200 414724 728206
rect 414672 728142 414724 728148
rect 417536 671562 417564 728414
rect 417524 671556 417576 671562
rect 417524 671498 417576 671504
rect 413108 654012 413160 654018
rect 413108 653954 413160 653960
rect 419928 651842 419956 729259
rect 420204 728614 420232 729395
rect 420284 729366 420336 729372
rect 420296 728886 420324 729366
rect 420284 728880 420336 728886
rect 420284 728822 420336 728828
rect 420756 728818 420784 729514
rect 432684 729294 432712 729514
rect 433084 729446 433112 729514
rect 433238 729446 433266 729514
rect 433084 729430 433266 729446
rect 433084 729424 433278 729430
rect 433084 729418 433226 729424
rect 431876 729288 431928 729294
rect 431876 729230 431928 729236
rect 432672 729288 432724 729294
rect 432672 729230 432724 729236
rect 420744 728812 420796 728818
rect 420744 728754 420796 728760
rect 420192 728608 420244 728614
rect 420192 728550 420244 728556
rect 419916 651836 419968 651842
rect 419916 651778 419968 651784
rect 431888 651774 431916 729230
rect 433084 728886 433112 729418
rect 433226 729366 433278 729372
rect 433238 729335 433266 729366
rect 434563 729362 434591 729514
rect 435274 729430 435302 729514
rect 436471 729494 436523 729552
rect 436396 729466 436523 729494
rect 435262 729424 435314 729430
rect 435262 729366 435314 729372
rect 434551 729356 434603 729362
rect 434551 729298 434603 729304
rect 433072 728880 433124 728886
rect 433072 728822 433124 728828
rect 434556 728750 434584 729298
rect 434544 728744 434596 728750
rect 434544 728686 434596 728692
rect 436396 728274 436424 729466
rect 437332 729430 437360 729514
rect 437500 729486 437620 729514
rect 437320 729424 437372 729430
rect 437320 729366 437372 729372
rect 437500 728478 437528 729486
rect 437592 729446 437620 729486
rect 437710 729446 437738 729514
rect 437592 729418 437738 729446
rect 438162 729430 438190 729514
rect 438374 729446 438402 729514
rect 438150 729424 438202 729430
rect 438150 729366 438202 729372
rect 438328 729418 438402 729446
rect 439110 729446 439138 729514
rect 439616 729486 439718 729514
rect 439110 729418 439184 729446
rect 438162 729333 438190 729366
rect 438148 729324 438204 729333
rect 438148 729259 438204 729268
rect 438328 728682 438356 729418
rect 439156 729362 439184 729418
rect 439144 729356 439196 729362
rect 439144 729298 439196 729304
rect 439156 728750 439184 729298
rect 439616 728818 439644 729486
rect 440720 729446 440932 729474
rect 441061 729446 441089 729514
rect 439604 728812 439656 728818
rect 439604 728754 439656 728760
rect 439144 728744 439196 728750
rect 439144 728686 439196 728692
rect 438316 728676 438368 728682
rect 438316 728618 438368 728624
rect 437488 728472 437540 728478
rect 437488 728414 437540 728420
rect 436384 728268 436436 728274
rect 436384 728210 436436 728216
rect 437500 658370 437528 728414
rect 437488 658364 437540 658370
rect 437488 658306 437540 658312
rect 440720 652998 440748 729446
rect 440904 729418 441089 729446
rect 441260 729424 441312 729430
rect 441983 729412 442011 729514
rect 441983 729384 442036 729412
rect 441260 729366 441312 729372
rect 441272 729333 441300 729366
rect 441258 729324 441314 729333
rect 441258 729259 441314 729268
rect 442008 728342 442036 729384
rect 445366 729310 445394 729514
rect 447528 729430 447556 729514
rect 447943 729484 447983 729540
rect 447804 729457 447983 729484
rect 459488 729486 459912 729514
rect 447804 729456 447970 729457
rect 447516 729424 447568 729430
rect 447516 729366 447568 729372
rect 445320 729282 445394 729310
rect 445320 728478 445348 729282
rect 447528 728886 447556 729366
rect 447698 729324 447754 729333
rect 447698 729259 447754 729268
rect 447516 728880 447568 728886
rect 447516 728822 447568 728828
rect 447712 728614 447740 729259
rect 447804 728818 447832 729456
rect 448066 729052 448122 729061
rect 448066 728987 448122 728996
rect 447792 728812 447844 728818
rect 447792 728754 447844 728760
rect 447700 728608 447752 728614
rect 447700 728550 447752 728556
rect 445308 728472 445360 728478
rect 445308 728414 445360 728420
rect 441996 728336 442048 728342
rect 441996 728278 442048 728284
rect 448080 724602 448108 728987
rect 448068 724596 448120 724602
rect 448068 724538 448120 724544
rect 450736 693180 450788 693186
rect 450736 693122 450788 693128
rect 440708 652992 440760 652998
rect 440708 652934 440760 652940
rect 431876 651768 431928 651774
rect 431876 651710 431928 651716
rect 405380 647484 405432 647490
rect 405380 647426 405432 647432
rect 426908 647484 426960 647490
rect 426908 647426 426960 647432
rect 412556 647416 412608 647422
rect 412556 647358 412608 647364
rect 407772 647144 407824 647150
rect 407772 647086 407824 647092
rect 407784 647030 407812 647086
rect 412568 647030 412596 647358
rect 417338 647316 417394 647325
rect 417338 647251 417394 647260
rect 417352 647030 417380 647251
rect 426920 647030 426948 647426
rect 446226 647180 446282 647189
rect 446226 647115 446282 647124
rect 446240 647030 446268 647115
rect 450748 647030 450776 693122
rect 459488 652930 459516 729486
rect 460293 729446 460321 729514
rect 460438 729446 460466 729514
rect 460293 729430 460466 729446
rect 461763 729446 461791 729514
rect 460293 729424 460478 729430
rect 460293 729418 460426 729424
rect 460293 729310 460321 729418
rect 461763 729418 461816 729446
rect 462478 729430 462506 729514
rect 460426 729366 460478 729372
rect 460438 729335 460466 729366
rect 460293 729282 460344 729310
rect 460316 728886 460344 729282
rect 460304 728880 460356 728886
rect 460304 728822 460356 728828
rect 461788 728750 461816 729418
rect 462466 729424 462518 729430
rect 462466 729366 462518 729372
rect 463674 729276 463702 729514
rect 464532 729430 464560 729514
rect 464520 729424 464572 729430
rect 464520 729366 464572 729372
rect 463628 729248 463702 729276
rect 463628 729022 463656 729248
rect 463616 729016 463668 729022
rect 463616 728958 463668 728964
rect 464916 728886 464944 729514
rect 465376 729430 465404 729514
rect 465364 729424 465416 729430
rect 465364 729366 465416 729372
rect 465560 729090 465588 729514
rect 465548 729084 465600 729090
rect 465548 729026 465600 729032
rect 463984 728880 464036 728886
rect 463984 728822 464036 728828
rect 464904 728880 464956 728886
rect 464904 728822 464956 728828
rect 461776 728744 461828 728750
rect 461776 728686 461828 728692
rect 460580 694676 460632 694682
rect 460580 694618 460632 694624
rect 459476 652924 459528 652930
rect 459476 652866 459528 652872
rect 455796 647144 455848 647150
rect 455796 647086 455848 647092
rect 455808 647030 455836 647086
rect 460592 647030 460620 694618
rect 463996 651706 464024 728822
rect 465560 728682 465588 729026
rect 466296 728750 466324 729514
rect 466894 729446 466922 729514
rect 466894 729418 466968 729446
rect 466940 728818 466968 729418
rect 468274 729276 468302 729514
rect 469171 729484 469223 729552
rect 472567 729484 472619 729552
rect 468872 729456 469223 729484
rect 472276 729456 472619 729484
rect 468584 729424 468636 729430
rect 468584 729366 468636 729372
rect 468596 729333 468624 729366
rect 468582 729324 468638 729333
rect 468274 729248 468348 729276
rect 468582 729259 468638 729268
rect 466928 728812 466980 728818
rect 466928 728754 466980 728760
rect 466284 728744 466336 728750
rect 466284 728686 466336 728692
rect 465548 728676 465600 728682
rect 465548 728618 465600 728624
rect 468320 728546 468348 729248
rect 468308 728540 468360 728546
rect 468308 728482 468360 728488
rect 464536 724596 464588 724602
rect 464536 724538 464588 724544
rect 464548 715762 464576 724538
rect 468872 722358 468900 729456
rect 472276 728886 472304 729456
rect 474734 729446 474762 729514
rect 475149 729486 475248 729514
rect 474734 729430 474788 729446
rect 474734 729424 474800 729430
rect 474734 729418 474748 729424
rect 474748 729366 474800 729372
rect 474760 728886 474788 729366
rect 474930 729324 474986 729333
rect 474930 729259 474986 729268
rect 474944 729022 474972 729259
rect 474932 729016 474984 729022
rect 474932 728958 474984 728964
rect 472264 728880 472316 728886
rect 472264 728822 472316 728828
rect 474748 728880 474800 728886
rect 474748 728822 474800 728828
rect 474944 728614 474972 728958
rect 475220 728818 475248 729486
rect 486536 729486 486912 729514
rect 487293 729486 487466 729514
rect 476402 729052 476458 729061
rect 476402 728987 476458 728996
rect 475208 728812 475260 728818
rect 475208 728754 475260 728760
rect 474932 728608 474984 728614
rect 474932 728550 474984 728556
rect 476416 728342 476444 728987
rect 476404 728336 476456 728342
rect 476404 728278 476456 728284
rect 468308 722352 468360 722358
rect 468308 722294 468360 722300
rect 468860 722352 468912 722358
rect 468860 722294 468912 722300
rect 464536 715756 464588 715762
rect 464536 715698 464588 715704
rect 468320 658370 468348 722294
rect 486536 718890 486564 729486
rect 487364 729430 487392 729486
rect 487352 729424 487404 729430
rect 487352 729366 487404 729372
rect 487364 728886 487392 729366
rect 488763 729362 488791 729514
rect 489474 729430 489502 729514
rect 490671 729484 490723 729552
rect 490671 729456 491072 729484
rect 489462 729424 489514 729430
rect 489462 729366 489514 729372
rect 488751 729356 488803 729362
rect 488744 729304 488751 729344
rect 488744 729298 488803 729304
rect 487352 728880 487404 728886
rect 487352 728822 487404 728828
rect 488744 728750 488772 729298
rect 488732 728744 488784 728750
rect 488732 728686 488784 728692
rect 491044 726846 491072 729456
rect 491532 729430 491560 729514
rect 491520 729424 491572 729430
rect 491520 729366 491572 729372
rect 491918 729310 491946 729514
rect 492362 729430 492390 729514
rect 492575 729486 492728 729514
rect 493304 729486 493464 729514
rect 492350 729424 492402 729430
rect 492350 729366 492402 729372
rect 491918 729282 491992 729310
rect 491964 728478 491992 729282
rect 492700 729090 492728 729486
rect 493436 729362 493464 729486
rect 493424 729356 493476 729362
rect 493424 729298 493476 729304
rect 492688 729084 492740 729090
rect 492688 729026 492740 729032
rect 492700 728614 492728 729026
rect 493436 728750 493464 729298
rect 493896 728818 493924 729514
rect 495249 729484 495301 729552
rect 496171 729484 496223 729552
rect 494816 729456 495301 729484
rect 495920 729456 496223 729484
rect 493884 728812 493936 728818
rect 493884 728754 493936 728760
rect 493424 728744 493476 728750
rect 493424 728686 493476 728692
rect 492688 728608 492740 728614
rect 492688 728550 492740 728556
rect 491952 728472 492004 728478
rect 491952 728414 492004 728420
rect 491032 726840 491084 726846
rect 491032 726782 491084 726788
rect 485972 718884 486024 718890
rect 485972 718826 486024 718832
rect 486524 718884 486576 718890
rect 486524 718826 486576 718832
rect 468768 715756 468820 715762
rect 468768 715698 468820 715704
rect 468780 711342 468808 715698
rect 468768 711336 468820 711342
rect 468768 711278 468820 711284
rect 478704 711336 478756 711342
rect 478704 711278 478756 711284
rect 474288 698824 474340 698830
rect 474288 698766 474340 698772
rect 468308 658364 468360 658370
rect 468308 658306 468360 658312
rect 463984 651700 464036 651706
rect 463984 651642 464036 651648
rect 470148 648504 470200 648510
rect 470148 648446 470200 648452
rect 470160 647030 470188 648446
rect 407784 647002 407904 647030
rect 412568 647002 412688 647030
rect 417352 647002 417472 647030
rect 426920 647002 427040 647030
rect 446240 647002 446360 647030
rect 450748 647002 451144 647030
rect 455808 647002 455928 647030
rect 460592 647002 460712 647030
rect 470160 647002 470280 647030
rect 474300 646917 474328 698766
rect 478716 696994 478744 711278
rect 478704 696988 478756 696994
rect 478704 696930 478756 696936
rect 485984 659458 486012 718826
rect 489744 696988 489796 696994
rect 489744 696930 489796 696936
rect 489756 687066 489784 696930
rect 489744 687060 489796 687066
rect 489744 687002 489796 687008
rect 489284 668292 489336 668298
rect 489284 668234 489336 668240
rect 485972 659452 486024 659458
rect 485972 659394 486024 659400
rect 479716 647484 479768 647490
rect 479716 647426 479768 647432
rect 479728 647030 479756 647426
rect 489296 647030 489324 668234
rect 494816 648442 494844 729456
rect 495448 729424 495500 729430
rect 495448 729366 495500 729372
rect 495460 729333 495488 729366
rect 495446 729324 495502 729333
rect 495446 729259 495502 729268
rect 495920 650822 495948 729456
rect 499579 729446 499607 729514
rect 501610 729460 501666 729469
rect 499579 729418 499628 729446
rect 499600 728478 499628 729418
rect 501734 729430 501762 729514
rect 502149 729486 502204 729514
rect 501722 729424 501774 729430
rect 501610 729395 501666 729404
rect 501426 729052 501482 729061
rect 500416 729016 500468 729022
rect 501426 728987 501482 728996
rect 500416 728958 500468 728964
rect 500428 728682 500456 728958
rect 500416 728676 500468 728682
rect 500416 728618 500468 728624
rect 499588 728472 499640 728478
rect 499588 728414 499640 728420
rect 499600 726914 499628 728414
rect 499588 726908 499640 726914
rect 499588 726850 499640 726856
rect 496368 687060 496420 687066
rect 496368 687002 496420 687008
rect 496380 682170 496408 687002
rect 496368 682164 496420 682170
rect 496368 682106 496420 682112
rect 501440 654018 501468 728987
rect 501624 728682 501652 729395
rect 501716 729372 501722 729412
rect 501716 729366 501774 729372
rect 501716 728886 501744 729366
rect 501704 728880 501756 728886
rect 501704 728822 501756 728828
rect 502176 728818 502204 729486
rect 513584 729486 514112 729514
rect 502164 728812 502216 728818
rect 502164 728754 502216 728760
rect 501612 728676 501664 728682
rect 501612 728618 501664 728624
rect 512468 705828 512520 705834
rect 512468 705770 512520 705776
rect 508144 698076 508196 698082
rect 508144 698018 508196 698024
rect 506304 689848 506356 689854
rect 506304 689790 506356 689796
rect 506316 665238 506344 689790
rect 506396 682164 506448 682170
rect 506396 682106 506448 682112
rect 506304 665232 506356 665238
rect 506304 665174 506356 665180
rect 506408 657282 506436 682106
rect 506396 657276 506448 657282
rect 506396 657218 506448 657224
rect 501428 654012 501480 654018
rect 501428 653954 501480 653960
rect 495908 650816 495960 650822
rect 495908 650758 495960 650764
rect 494804 648436 494856 648442
rect 494804 648378 494856 648384
rect 494068 647416 494120 647422
rect 494068 647358 494120 647364
rect 494080 647030 494108 647358
rect 503636 647212 503688 647218
rect 503636 647154 503688 647160
rect 503648 647030 503676 647154
rect 508156 647030 508184 698018
rect 479728 647002 479848 647030
rect 489296 647002 489416 647030
rect 494080 647002 494200 647030
rect 503648 647002 503768 647030
rect 508156 647002 508552 647030
rect 512480 646917 512508 705770
rect 513584 703590 513612 729486
rect 514504 729446 514532 729514
rect 514638 729446 514666 729514
rect 514504 729430 514666 729446
rect 514504 729424 514678 729430
rect 514504 729418 514626 729424
rect 514504 728886 514532 729418
rect 514626 729366 514678 729372
rect 514638 729335 514666 729366
rect 515976 729362 516004 729514
rect 516674 729430 516702 729514
rect 516662 729424 516714 729430
rect 516662 729366 516714 729372
rect 515964 729356 516016 729362
rect 515964 729298 516016 729304
rect 514492 728880 514544 728886
rect 514492 728822 514544 728828
rect 515976 728750 516004 729298
rect 517883 729294 517911 729514
rect 518736 729430 518764 729514
rect 519110 729486 519224 729514
rect 518724 729424 518776 729430
rect 518724 729366 518776 729372
rect 519196 729294 519224 729486
rect 519564 729430 519592 729514
rect 519656 729486 519803 729514
rect 519552 729424 519604 729430
rect 519552 729366 519604 729372
rect 516884 729288 516936 729294
rect 516884 729230 516936 729236
rect 517871 729288 517923 729294
rect 517871 729230 517923 729236
rect 519184 729288 519236 729294
rect 519184 729230 519236 729236
rect 515964 728744 516016 728750
rect 515964 728686 516016 728692
rect 513572 703584 513624 703590
rect 513572 703526 513624 703532
rect 516896 668298 516924 729230
rect 516884 668292 516936 668298
rect 516884 668234 516936 668240
rect 514032 657276 514084 657282
rect 514032 657218 514084 657224
rect 514044 649530 514072 657218
rect 519196 653950 519224 729230
rect 519656 728614 519684 729486
rect 520504 729446 520532 729514
rect 521078 729484 521130 729552
rect 521078 729456 521432 729484
rect 520484 729418 520532 729446
rect 520484 729362 520512 729418
rect 520472 729356 520524 729362
rect 520472 729298 520524 729304
rect 520484 728750 520512 729298
rect 521404 728886 521432 729456
rect 522462 729208 522490 729514
rect 522680 729424 522732 729430
rect 522680 729366 522732 729372
rect 522588 729356 522640 729362
rect 522692 729333 522720 729366
rect 523382 729362 523410 729514
rect 526779 729362 526807 729514
rect 528948 729430 528976 729514
rect 529316 729486 529377 729514
rect 528936 729424 528988 729430
rect 528936 729366 528988 729372
rect 523370 729356 523422 729362
rect 522588 729298 522640 729304
rect 522678 729324 522734 729333
rect 522462 729180 522536 729208
rect 522508 729022 522536 729180
rect 522496 729016 522548 729022
rect 522496 728958 522548 728964
rect 521392 728880 521444 728886
rect 521392 728822 521444 728828
rect 520472 728744 520524 728750
rect 520472 728686 520524 728692
rect 519644 728608 519696 728614
rect 519644 728550 519696 728556
rect 522496 658364 522548 658370
rect 522496 658306 522548 658312
rect 519184 653944 519236 653950
rect 519184 653886 519236 653892
rect 517988 652924 518040 652930
rect 517988 652866 518040 652872
rect 514032 649524 514084 649530
rect 514032 649466 514084 649472
rect 518000 647030 518028 652866
rect 522508 647030 522536 658306
rect 522600 656194 522628 729298
rect 523370 729298 523422 729304
rect 526767 729356 526819 729362
rect 526767 729298 526819 729304
rect 522678 729259 522734 729268
rect 528948 728818 528976 729366
rect 529118 729324 529174 729333
rect 529118 729259 529174 729268
rect 529132 729090 529160 729259
rect 529120 729084 529172 729090
rect 529120 729026 529172 729032
rect 529210 729052 529266 729061
rect 528936 728812 528988 728818
rect 528936 728754 528988 728760
rect 529132 728682 529160 729026
rect 529210 728987 529266 728996
rect 529120 728676 529172 728682
rect 529120 728618 529172 728624
rect 522588 656188 522640 656194
rect 522588 656130 522640 656136
rect 529224 652930 529252 728987
rect 529316 728886 529344 729486
rect 529304 728880 529356 728886
rect 529304 728822 529356 728828
rect 541276 704746 541304 729514
rect 541684 729494 541730 729546
rect 541826 729494 541878 729552
rect 541368 729466 541948 729494
rect 541368 728818 541396 729466
rect 541920 729430 541948 729466
rect 541908 729424 541960 729430
rect 541908 729366 541960 729372
rect 543163 729362 543191 729514
rect 543874 729430 543902 729514
rect 545071 729484 545123 729552
rect 544496 729456 545123 729484
rect 543862 729424 543914 729430
rect 543862 729366 543914 729372
rect 543151 729356 543203 729362
rect 543116 729304 543151 729310
rect 543116 729298 543203 729304
rect 543116 729282 543191 729298
rect 541356 728812 541408 728818
rect 541356 728754 541408 728760
rect 543116 728750 543144 729282
rect 543104 728744 543156 728750
rect 543104 728686 543156 728692
rect 541264 704740 541316 704746
rect 541264 704682 541316 704688
rect 536756 671556 536808 671562
rect 536756 671498 536808 671504
rect 532340 665164 532392 665170
rect 532340 665106 532392 665112
rect 529212 652924 529264 652930
rect 529212 652866 529264 652872
rect 532352 647030 532380 665106
rect 518000 647002 518120 647030
rect 522508 647002 522904 647030
rect 532352 647002 532656 647030
rect 536768 646917 536796 671498
rect 541172 660540 541224 660546
rect 541172 660482 541224 660488
rect 541184 646917 541212 660482
rect 544496 647286 544524 729456
rect 545922 729430 545950 729514
rect 545910 729424 545962 729430
rect 545910 729366 545962 729372
rect 546310 729310 546338 729514
rect 546750 729430 546778 729514
rect 546738 729424 546790 729430
rect 546738 729366 546790 729372
rect 546750 729333 546778 729366
rect 546736 729324 546792 729333
rect 546310 729282 546364 729310
rect 546336 728478 546364 729282
rect 546736 729259 546792 729268
rect 546980 728750 547008 729514
rect 547716 729362 547744 729514
rect 548290 729446 548318 729514
rect 549649 729474 549700 729552
rect 550571 729484 550623 729552
rect 548268 729418 548318 729446
rect 548912 729446 549700 729474
rect 550476 729456 550623 729484
rect 547704 729356 547756 729362
rect 547704 729298 547756 729304
rect 547716 728818 547744 729298
rect 548268 728886 548296 729418
rect 548256 728880 548308 728886
rect 548256 728822 548308 728828
rect 547704 728812 547756 728818
rect 547704 728754 547756 728760
rect 546968 728744 547020 728750
rect 546968 728686 547020 728692
rect 546980 728614 547008 728686
rect 546968 728608 547020 728614
rect 546968 728550 547020 728556
rect 546324 728472 546376 728478
rect 546324 728414 546376 728420
rect 548912 657214 548940 729446
rect 550476 728614 550504 729456
rect 553040 729424 553092 729430
rect 553040 729366 553092 729372
rect 553052 729333 553080 729366
rect 553038 729324 553094 729333
rect 553038 729259 553094 729268
rect 553972 729158 554000 729514
rect 556134 729430 556162 729514
rect 556122 729424 556174 729430
rect 556174 729372 556208 729412
rect 556122 729366 556208 729372
rect 554694 729188 554750 729197
rect 553316 729152 553368 729158
rect 553316 729094 553368 729100
rect 553960 729152 554012 729158
rect 554694 729123 554750 729132
rect 553960 729094 554012 729100
rect 550464 728608 550516 728614
rect 550464 728550 550516 728556
rect 553328 728478 553356 729094
rect 554708 729090 554736 729123
rect 554696 729084 554748 729090
rect 554696 729026 554748 729032
rect 555524 729084 555576 729090
rect 555524 729026 555576 729032
rect 555536 728886 555564 729026
rect 555524 728880 555576 728886
rect 555524 728822 555576 728828
rect 556180 728682 556208 729366
rect 556258 729188 556314 729197
rect 556258 729123 556314 729132
rect 556272 728886 556300 729123
rect 556548 729090 556576 729514
rect 568484 729486 568536 729514
rect 568893 729486 568996 729514
rect 556536 729084 556588 729090
rect 556536 729026 556588 729032
rect 557088 729084 557140 729090
rect 557088 729026 557140 729032
rect 556260 728880 556312 728886
rect 556260 728822 556312 728828
rect 556168 728676 556220 728682
rect 556168 728618 556220 728624
rect 553316 728472 553368 728478
rect 553316 728414 553368 728420
rect 548900 657208 548952 657214
rect 548900 657150 548952 657156
rect 546692 654012 546744 654018
rect 546692 653954 546744 653960
rect 544484 647280 544536 647286
rect 544484 647222 544536 647228
rect 546704 647030 546732 653954
rect 553328 653950 553356 728414
rect 557100 695430 557128 729026
rect 568508 728886 568536 729486
rect 568968 729446 568996 729486
rect 569038 729446 569066 729514
rect 568968 729418 569066 729446
rect 570348 729430 570376 729514
rect 570336 729424 570388 729430
rect 568968 729362 568996 729418
rect 570336 729366 570388 729372
rect 568956 729356 569008 729362
rect 568956 729298 569008 729304
rect 568864 728948 568916 728954
rect 568864 728890 568916 728896
rect 568496 728880 568548 728886
rect 568496 728822 568548 728828
rect 568876 725758 568904 728890
rect 568968 728682 568996 729298
rect 570348 728818 570376 729366
rect 571074 729362 571102 729514
rect 572280 729362 572308 729514
rect 573132 729446 573160 729514
rect 573200 729486 573412 729514
rect 573200 729446 573228 729486
rect 573132 729418 573228 729446
rect 573384 729446 573412 729486
rect 573522 729446 573550 729514
rect 573384 729430 573550 729446
rect 573962 729430 573990 729514
rect 574175 729486 574240 729514
rect 574904 729498 575068 729514
rect 574904 729492 575080 729498
rect 574904 729486 575028 729492
rect 573384 729424 573562 729430
rect 573384 729418 573510 729424
rect 573132 729362 573160 729418
rect 573510 729366 573562 729372
rect 573950 729424 574002 729430
rect 573950 729366 574002 729372
rect 571062 729356 571114 729362
rect 571062 729298 571114 729304
rect 572268 729356 572320 729362
rect 572268 729298 572320 729304
rect 573120 729356 573172 729362
rect 573120 729298 573172 729304
rect 570336 728812 570388 728818
rect 570336 728754 570388 728760
rect 574212 728682 574240 729486
rect 574948 728750 574976 729486
rect 575478 729474 575530 729552
rect 576849 729484 576901 729552
rect 575478 729446 575896 729474
rect 575028 729434 575080 729440
rect 574936 728744 574988 728750
rect 574936 728686 574988 728692
rect 568956 728676 569008 728682
rect 568956 728618 569008 728624
rect 574200 728676 574252 728682
rect 574200 728618 574252 728624
rect 575868 728478 575896 729446
rect 576512 729456 576901 729484
rect 577771 729474 577823 729552
rect 576512 728954 576540 729456
rect 577432 729446 577823 729474
rect 577052 729424 577104 729430
rect 577052 729366 577104 729372
rect 577064 729333 577092 729366
rect 577050 729324 577106 729333
rect 577050 729259 577106 729268
rect 576500 728948 576552 728954
rect 576500 728890 576552 728896
rect 575856 728472 575908 728478
rect 575856 728414 575908 728420
rect 569876 726772 569928 726778
rect 569876 726714 569928 726720
rect 568864 725752 568916 725758
rect 568864 725694 568916 725700
rect 557088 695424 557140 695430
rect 557088 695366 557140 695372
rect 569232 667204 569284 667210
rect 569232 667146 569284 667152
rect 569244 664014 569272 667146
rect 569232 664008 569284 664014
rect 569232 663950 569284 663956
rect 553316 653944 553368 653950
rect 553316 653886 553368 653892
rect 561228 651700 561280 651706
rect 561228 651642 561280 651648
rect 551660 650136 551712 650142
rect 551660 650078 551712 650084
rect 551672 647030 551700 650078
rect 556444 647212 556496 647218
rect 556444 647154 556496 647160
rect 556456 647030 556484 647154
rect 561240 647030 561268 651642
rect 569232 649116 569284 649122
rect 569232 649058 569284 649064
rect 569244 648510 569272 649058
rect 569232 648504 569284 648510
rect 569232 648446 569284 648452
rect 546704 647002 547008 647030
rect 551672 647002 551792 647030
rect 556456 647002 556576 647030
rect 561240 647002 561360 647030
rect 569888 646917 569916 726714
rect 575396 719088 575448 719094
rect 575396 719030 575448 719036
rect 574752 664008 574804 664014
rect 574752 663950 574804 663956
rect 574764 658370 574792 663950
rect 574752 658364 574804 658370
rect 574752 658306 574804 658312
rect 575408 647030 575436 719030
rect 576512 666802 576540 728890
rect 577432 728886 577460 729446
rect 577420 728880 577472 728886
rect 577420 728822 577472 728828
rect 577616 728818 577644 729446
rect 581179 729430 581207 729514
rect 583320 729430 583348 729514
rect 581167 729424 581219 729430
rect 581167 729366 581219 729372
rect 583308 729424 583360 729430
rect 583308 729366 583360 729372
rect 578430 729052 578486 729061
rect 578430 728987 578486 728996
rect 577604 728812 577656 728818
rect 577604 728754 577656 728760
rect 578444 725690 578472 728987
rect 583320 728886 583348 729366
rect 583749 729310 583777 729514
rect 595280 729486 595400 729514
rect 594164 729424 594216 729430
rect 594164 729366 594216 729372
rect 583688 729282 583777 729310
rect 583582 728916 583638 728925
rect 583308 728880 583360 728886
rect 583582 728851 583638 728860
rect 583308 728822 583360 728828
rect 583596 728818 583624 728851
rect 583584 728812 583636 728818
rect 583584 728754 583636 728760
rect 583688 728478 583716 729282
rect 594176 728886 594204 729366
rect 594164 728880 594216 728886
rect 594164 728822 594216 728828
rect 583676 728472 583728 728478
rect 583676 728414 583728 728420
rect 584688 728200 584740 728206
rect 584688 728142 584740 728148
rect 584700 726778 584728 728142
rect 589104 728064 589156 728070
rect 589104 728006 589156 728012
rect 585608 727860 585660 727866
rect 585608 727802 585660 727808
rect 584688 726772 584740 726778
rect 584688 726714 584740 726720
rect 583584 725752 583636 725758
rect 583584 725694 583636 725700
rect 578432 725684 578484 725690
rect 578432 725626 578484 725632
rect 583596 724194 583624 725694
rect 583584 724188 583636 724194
rect 583584 724130 583636 724136
rect 585620 723514 585648 727802
rect 588000 724188 588052 724194
rect 588000 724130 588052 724136
rect 585608 723508 585660 723514
rect 585608 723450 585660 723456
rect 588012 711342 588040 724130
rect 589116 722290 589144 728006
rect 593520 727928 593572 727934
rect 593520 727870 593572 727876
rect 593532 722698 593560 727870
rect 594624 726908 594676 726914
rect 594624 726850 594676 726856
rect 594636 723514 594664 726850
rect 594624 723508 594676 723514
rect 594624 723450 594676 723456
rect 593520 722692 593572 722698
rect 593520 722634 593572 722640
rect 594716 722692 594768 722698
rect 594716 722634 594768 722640
rect 589104 722284 589156 722290
rect 589104 722226 589156 722232
rect 594624 722284 594676 722290
rect 594624 722226 594676 722232
rect 588000 711336 588052 711342
rect 588000 711278 588052 711284
rect 594636 710322 594664 722226
rect 594728 712634 594756 722634
rect 594716 712628 594768 712634
rect 594716 712570 594768 712576
rect 594624 710316 594676 710322
rect 594624 710258 594676 710264
rect 595280 708010 595308 729486
rect 595372 729446 595400 729486
rect 595484 729446 595512 729514
rect 595372 729418 595512 729446
rect 595893 729446 595921 729514
rect 596038 729446 596066 729514
rect 595893 729430 596066 729446
rect 597363 729430 597391 729514
rect 595881 729424 596066 729430
rect 595933 729418 596066 729424
rect 597351 729424 597403 729430
rect 595881 729366 595933 729372
rect 597350 729372 597351 729412
rect 597350 729366 597403 729372
rect 597350 729276 597378 729366
rect 598074 729362 598102 729514
rect 598062 729356 598114 729362
rect 598062 729298 598114 729304
rect 599282 729294 599310 729514
rect 600132 729362 600160 729514
rect 600524 729362 600552 729514
rect 600120 729356 600172 729362
rect 600120 729298 600172 729304
rect 600512 729356 600564 729362
rect 600962 729333 600990 729514
rect 600512 729298 600564 729304
rect 600948 729324 601004 729333
rect 597304 729248 597378 729276
rect 598580 729288 598632 729294
rect 597304 728750 597332 729248
rect 598580 729230 598632 729236
rect 599270 729288 599322 729294
rect 599270 729230 599322 729236
rect 597292 728744 597344 728750
rect 597292 728686 597344 728692
rect 597936 728404 597988 728410
rect 597936 728346 597988 728352
rect 596832 726840 596884 726846
rect 596832 726782 596884 726788
rect 595728 726772 595780 726778
rect 595728 726714 595780 726720
rect 595740 720658 595768 726714
rect 596844 721474 596872 726782
rect 596832 721468 596884 721474
rect 596832 721410 596884 721416
rect 595728 720652 595780 720658
rect 595728 720594 595780 720600
rect 596832 720652 596884 720658
rect 596832 720594 596884 720600
rect 596844 714538 596872 720594
rect 597948 719094 597976 728346
rect 597936 719088 597988 719094
rect 597936 719030 597988 719036
rect 596832 714532 596884 714538
rect 596832 714474 596884 714480
rect 597936 714532 597988 714538
rect 597936 714474 597988 714480
rect 595268 708004 595320 708010
rect 595268 707946 595320 707952
rect 597948 700462 597976 714474
rect 598028 710316 598080 710322
rect 598028 710258 598080 710264
rect 598040 702502 598068 710258
rect 598028 702496 598080 702502
rect 598028 702438 598080 702444
rect 597936 700456 597988 700462
rect 597936 700398 597988 700404
rect 596832 698960 596884 698966
rect 596832 698902 596884 698908
rect 576960 698756 577012 698762
rect 576960 698698 577012 698704
rect 576972 689242 577000 698698
rect 576960 689236 577012 689242
rect 576960 689178 577012 689184
rect 590208 689236 590260 689242
rect 590208 689178 590260 689184
rect 590220 681558 590248 689178
rect 596844 684550 596872 698902
rect 596832 684544 596884 684550
rect 596832 684486 596884 684492
rect 590208 681552 590260 681558
rect 590208 681494 590260 681500
rect 576500 666796 576552 666802
rect 576500 666738 576552 666744
rect 598592 666530 598620 729230
rect 600524 728818 600552 729298
rect 600948 729259 600950 729268
rect 601002 729259 601004 729268
rect 600950 729230 601002 729236
rect 600962 729199 600990 729230
rect 600512 728812 600564 728818
rect 600512 728754 600564 728760
rect 601168 728682 601196 729514
rect 601904 729430 601932 729514
rect 601892 729424 601944 729430
rect 601892 729366 601944 729372
rect 601904 728750 601932 729366
rect 602502 729276 602530 729514
rect 603861 729362 603889 729514
rect 604783 729430 604811 729514
rect 604771 729424 604823 729430
rect 604771 729366 604823 729372
rect 603849 729356 603901 729362
rect 604783 729333 604811 729366
rect 608179 729362 608207 729514
rect 610334 729486 610488 729514
rect 610460 729430 610488 729486
rect 610448 729424 610500 729430
rect 610448 729366 610500 729372
rect 608167 729356 608219 729362
rect 603849 729298 603901 729304
rect 604769 729324 604825 729333
rect 602502 729248 602576 729276
rect 604769 729259 604825 729268
rect 608165 729324 608167 729333
rect 608219 729324 608221 729333
rect 608165 729259 608221 729268
rect 602548 729090 602576 729248
rect 602536 729084 602588 729090
rect 602536 729026 602588 729032
rect 610460 728818 610488 729366
rect 610749 729310 610777 729514
rect 610736 729282 610777 729310
rect 611458 729324 611514 729333
rect 610736 729090 610764 729282
rect 611458 729259 611514 729268
rect 610724 729084 610776 729090
rect 610724 729026 610776 729032
rect 611472 728886 611500 729259
rect 619556 729016 619608 729022
rect 619556 728958 619608 728964
rect 611460 728880 611512 728886
rect 611460 728822 611512 728828
rect 610448 728812 610500 728818
rect 610448 728754 610500 728760
rect 601892 728744 601944 728750
rect 601892 728686 601944 728692
rect 601156 728676 601208 728682
rect 601156 728618 601208 728624
rect 610080 728336 610132 728342
rect 610080 728278 610132 728284
rect 600144 728268 600196 728274
rect 600144 728210 600196 728216
rect 599040 723440 599092 723446
rect 599040 723382 599092 723388
rect 599052 713518 599080 723382
rect 600156 713586 600184 728210
rect 600236 728132 600288 728138
rect 600236 728074 600288 728080
rect 600248 722154 600276 728074
rect 600328 727996 600380 728002
rect 600328 727938 600380 727944
rect 600236 722148 600288 722154
rect 600236 722090 600288 722096
rect 600340 721338 600368 727938
rect 607320 723508 607372 723514
rect 607320 723450 607372 723456
rect 602352 722148 602404 722154
rect 602352 722090 602404 722096
rect 600328 721332 600380 721338
rect 600328 721274 600380 721280
rect 600144 713580 600196 713586
rect 600144 713522 600196 713528
rect 599040 713512 599092 713518
rect 599040 713454 599092 713460
rect 602364 712770 602392 722090
rect 603732 721468 603784 721474
rect 603732 721410 603784 721416
rect 603744 716850 603772 721410
rect 604560 721332 604612 721338
rect 604560 721274 604612 721280
rect 603732 716844 603784 716850
rect 603732 716786 603784 716792
rect 602352 712764 602404 712770
rect 602352 712706 602404 712712
rect 600144 712628 600196 712634
rect 600144 712570 600196 712576
rect 600156 708350 600184 712570
rect 600144 708344 600196 708350
rect 600144 708286 600196 708292
rect 602352 708344 602404 708350
rect 602352 708286 602404 708292
rect 600144 700456 600196 700462
rect 600144 700398 600196 700404
rect 600156 683122 600184 700398
rect 602364 684822 602392 708286
rect 604572 699850 604600 721274
rect 607332 720114 607360 723450
rect 610092 720182 610120 728278
rect 610080 720176 610132 720182
rect 610080 720118 610132 720124
rect 616704 720176 616756 720182
rect 616704 720118 616756 720124
rect 607320 720108 607372 720114
rect 607320 720050 607372 720056
rect 613484 720108 613536 720114
rect 613484 720050 613536 720056
rect 605848 719088 605900 719094
rect 605848 719030 605900 719036
rect 605860 717938 605888 719030
rect 605848 717932 605900 717938
rect 605848 717874 605900 717880
rect 613392 717932 613444 717938
rect 613392 717874 613444 717880
rect 608976 716844 609028 716850
rect 608976 716786 609028 716792
rect 604836 713580 604888 713586
rect 604836 713522 604888 713528
rect 604652 712764 604704 712770
rect 604652 712706 604704 712712
rect 604664 706378 604692 712706
rect 604744 711336 604796 711342
rect 604744 711278 604796 711284
rect 604756 707330 604784 711278
rect 604744 707324 604796 707330
rect 604744 707266 604796 707272
rect 604652 706372 604704 706378
rect 604652 706314 604704 706320
rect 604848 700530 604876 713522
rect 606768 713512 606820 713518
rect 606768 713454 606820 713460
rect 605848 707324 605900 707330
rect 605848 707266 605900 707272
rect 605664 702496 605716 702502
rect 605664 702438 605716 702444
rect 604836 700524 604888 700530
rect 604836 700466 604888 700472
rect 605676 700394 605704 702438
rect 605860 701074 605888 707266
rect 606780 707058 606808 713454
rect 608988 708350 609016 716786
rect 608976 708344 609028 708350
rect 608976 708286 609028 708292
rect 611184 708344 611236 708350
rect 611184 708286 611236 708292
rect 606768 707052 606820 707058
rect 606768 706994 606820 707000
rect 608056 707052 608108 707058
rect 608056 706994 608108 707000
rect 607872 706372 607924 706378
rect 607872 706314 607924 706320
rect 605848 701068 605900 701074
rect 605848 701010 605900 701016
rect 605664 700388 605716 700394
rect 605664 700330 605716 700336
rect 604560 699844 604612 699850
rect 604560 699786 604612 699792
rect 605664 699844 605716 699850
rect 605664 699786 605716 699792
rect 602352 684816 602404 684822
rect 602352 684758 602404 684764
rect 603548 684544 603600 684550
rect 603548 684486 603600 684492
rect 600144 683116 600196 683122
rect 600144 683058 600196 683064
rect 603456 683116 603508 683122
rect 603456 683058 603508 683064
rect 600144 681552 600196 681558
rect 600144 681494 600196 681500
rect 600156 671562 600184 681494
rect 603468 673398 603496 683058
rect 603560 674894 603588 684486
rect 605676 676526 605704 699786
rect 607884 676662 607912 706314
rect 607964 701068 608016 701074
rect 607964 701010 608016 701016
rect 607976 681490 608004 701010
rect 608068 692098 608096 706994
rect 610080 700524 610132 700530
rect 610080 700466 610132 700472
rect 608056 692092 608108 692098
rect 608056 692034 608108 692040
rect 607964 681484 608016 681490
rect 607964 681426 608016 681432
rect 610092 681014 610120 700466
rect 611196 690670 611224 708286
rect 611276 700388 611328 700394
rect 611276 700330 611328 700336
rect 611184 690664 611236 690670
rect 611184 690606 611236 690612
rect 611184 684816 611236 684822
rect 611184 684758 611236 684764
rect 610080 681008 610132 681014
rect 610080 680950 610132 680956
rect 607872 676656 607924 676662
rect 607872 676598 607924 676604
rect 608976 676656 609028 676662
rect 608976 676598 609028 676604
rect 605664 676520 605716 676526
rect 605664 676462 605716 676468
rect 606860 676520 606912 676526
rect 606860 676462 606912 676468
rect 603548 674888 603600 674894
rect 603548 674830 603600 674836
rect 603456 673392 603508 673398
rect 603456 673334 603508 673340
rect 606768 673392 606820 673398
rect 606768 673334 606820 673340
rect 600144 671556 600196 671562
rect 600144 671498 600196 671504
rect 598580 666524 598632 666530
rect 598580 666466 598632 666472
rect 605664 666252 605716 666258
rect 605664 666194 605716 666200
rect 594624 666116 594676 666122
rect 594624 666058 594676 666064
rect 584228 662784 584280 662790
rect 584228 662726 584280 662732
rect 575408 647002 575712 647030
rect 584240 646917 584268 662726
rect 584688 658364 584740 658370
rect 584688 658306 584740 658312
rect 584700 656194 584728 658306
rect 594636 657214 594664 666058
rect 598580 666048 598632 666054
rect 598580 665990 598632 665996
rect 594624 657208 594676 657214
rect 594624 657150 594676 657156
rect 584688 656188 584740 656194
rect 584688 656130 584740 656136
rect 595728 656188 595780 656194
rect 595728 656130 595780 656136
rect 595740 651774 595768 656130
rect 595728 651768 595780 651774
rect 595728 651710 595780 651716
rect 594716 647280 594768 647286
rect 594716 647222 594768 647228
rect 594728 647030 594756 647222
rect 594728 647002 594848 647030
rect 598592 646917 598620 665990
rect 604652 665028 604704 665034
rect 604652 664970 604704 664976
rect 604560 663940 604612 663946
rect 604560 663882 604612 663888
rect 604572 661770 604600 663882
rect 604664 662790 604692 664970
rect 604652 662784 604704 662790
rect 604652 662726 604704 662732
rect 604560 661764 604612 661770
rect 604560 661706 604612 661712
rect 605676 656262 605704 666194
rect 606780 660138 606808 673334
rect 606872 666122 606900 676462
rect 606860 666116 606912 666122
rect 606860 666058 606912 666064
rect 608988 664558 609016 676598
rect 610816 674888 610868 674894
rect 610816 674830 610868 674836
rect 610828 669386 610856 674830
rect 610816 669380 610868 669386
rect 610816 669322 610868 669328
rect 611196 666394 611224 684758
rect 611288 681150 611316 700330
rect 613404 699918 613432 717874
rect 613496 713586 613524 720050
rect 613484 713580 613536 713586
rect 613484 713522 613536 713528
rect 614588 713580 614640 713586
rect 614588 713522 614640 713528
rect 614600 700054 614628 713522
rect 614588 700048 614640 700054
rect 614588 699990 614640 699996
rect 615600 700048 615652 700054
rect 615600 699990 615652 699996
rect 613392 699912 613444 699918
rect 613392 699854 613444 699860
rect 614496 699912 614548 699918
rect 614496 699854 614548 699860
rect 611460 692092 611512 692098
rect 611460 692034 611512 692040
rect 611276 681144 611328 681150
rect 611276 681086 611328 681092
rect 611472 681082 611500 692034
rect 612288 690664 612340 690670
rect 612288 690606 612340 690612
rect 611460 681076 611512 681082
rect 611460 681018 611512 681024
rect 612300 671050 612328 690606
rect 614508 684618 614536 699854
rect 614496 684612 614548 684618
rect 614496 684554 614548 684560
rect 612564 681484 612616 681490
rect 612564 681426 612616 681432
rect 612472 681144 612524 681150
rect 612472 681086 612524 681092
rect 612484 676186 612512 681086
rect 612576 677818 612604 681426
rect 614588 681076 614640 681082
rect 614588 681018 614640 681024
rect 613392 681008 613444 681014
rect 613392 680950 613444 680956
rect 612564 677812 612616 677818
rect 612564 677754 612616 677760
rect 612472 676180 612524 676186
rect 612472 676122 612524 676128
rect 612380 671556 612432 671562
rect 612380 671498 612432 671504
rect 612116 671022 612328 671050
rect 611184 666388 611236 666394
rect 611184 666330 611236 666336
rect 610264 665096 610316 665102
rect 610264 665038 610316 665044
rect 608976 664552 609028 664558
rect 608976 664494 609028 664500
rect 610080 663872 610132 663878
rect 610080 663814 610132 663820
rect 606768 660132 606820 660138
rect 606768 660074 606820 660080
rect 609160 660132 609212 660138
rect 609160 660074 609212 660080
rect 605664 656256 605716 656262
rect 605664 656198 605716 656204
rect 609172 652930 609200 660074
rect 610092 658982 610120 663814
rect 610172 661764 610224 661770
rect 610172 661706 610224 661712
rect 610080 658976 610132 658982
rect 610080 658918 610132 658924
rect 610184 655106 610212 661706
rect 610276 657282 610304 665038
rect 612116 661362 612144 671022
rect 612196 664552 612248 664558
rect 612196 664494 612248 664500
rect 612104 661356 612156 661362
rect 612104 661298 612156 661304
rect 612208 659406 612236 664494
rect 612116 659378 612236 659406
rect 610264 657276 610316 657282
rect 610264 657218 610316 657224
rect 610172 655100 610224 655106
rect 610172 655042 610224 655048
rect 609160 652924 609212 652930
rect 609160 652866 609212 652872
rect 607872 651768 607924 651774
rect 607872 651710 607924 651716
rect 607884 649598 607912 651710
rect 612116 650414 612144 659378
rect 612288 658976 612340 658982
rect 612288 658918 612340 658924
rect 612196 657208 612248 657214
rect 612196 657150 612248 657156
rect 612208 651541 612236 657150
rect 612194 651532 612250 651541
rect 612194 651467 612250 651476
rect 612300 650861 612328 658918
rect 612392 651677 612420 671498
rect 613404 668774 613432 680950
rect 614496 677812 614548 677818
rect 614496 677754 614548 677760
rect 613392 668768 613444 668774
rect 613392 668710 613444 668716
rect 612932 666728 612984 666734
rect 612932 666670 612984 666676
rect 612378 651668 612434 651677
rect 612378 651603 612434 651612
rect 612286 650852 612342 650861
rect 612286 650787 612342 650796
rect 612104 650408 612156 650414
rect 612104 650350 612156 650356
rect 607872 649592 607924 649598
rect 607872 649534 607924 649540
rect 612944 646917 612972 666670
rect 613392 666388 613444 666394
rect 613392 666330 613444 666336
rect 613404 650686 613432 666330
rect 613484 666116 613536 666122
rect 613484 666058 613536 666064
rect 613496 659526 613524 666058
rect 614508 662926 614536 677754
rect 614600 676322 614628 681018
rect 614588 676316 614640 676322
rect 614588 676258 614640 676264
rect 614588 676180 614640 676186
rect 614588 676122 614640 676128
rect 614496 662920 614548 662926
rect 614496 662862 614548 662868
rect 614496 662784 614548 662790
rect 614496 662726 614548 662732
rect 613484 659520 613536 659526
rect 613484 659462 613536 659468
rect 614404 656256 614456 656262
rect 614404 656198 614456 656204
rect 614416 651949 614444 656198
rect 614402 651940 614458 651949
rect 614402 651875 614458 651884
rect 613300 650680 613352 650686
rect 613300 650622 613352 650628
rect 613392 650680 613444 650686
rect 613392 650622 613444 650628
rect 613312 650482 613340 650622
rect 613300 650476 613352 650482
rect 613300 650418 613352 650424
rect 614508 650346 614536 662726
rect 614600 659458 614628 676122
rect 615612 667686 615640 699990
rect 615692 684612 615744 684618
rect 615692 684554 615744 684560
rect 615600 667680 615652 667686
rect 615600 667622 615652 667628
rect 615600 666184 615652 666190
rect 615600 666126 615652 666132
rect 615612 663878 615640 666126
rect 615600 663872 615652 663878
rect 615600 663814 615652 663820
rect 615704 661906 615732 684554
rect 616716 684142 616744 720118
rect 616704 684136 616756 684142
rect 616704 684078 616756 684084
rect 617900 684136 617952 684142
rect 617900 684078 617952 684084
rect 616704 676316 616756 676322
rect 616704 676258 616756 676264
rect 615784 666660 615836 666666
rect 615784 666602 615836 666608
rect 615692 661900 615744 661906
rect 615692 661842 615744 661848
rect 614588 659452 614640 659458
rect 614588 659394 614640 659400
rect 615692 659452 615744 659458
rect 615692 659394 615744 659400
rect 615508 655100 615560 655106
rect 615508 655042 615560 655048
rect 614496 650340 614548 650346
rect 614496 650282 614548 650288
rect 615520 648782 615548 655042
rect 615600 652924 615652 652930
rect 615600 652866 615652 652872
rect 615612 651094 615640 652866
rect 615704 651842 615732 659394
rect 615796 658506 615824 666602
rect 615968 664960 616020 664966
rect 615968 664902 616020 664908
rect 615784 658500 615836 658506
rect 615784 658442 615836 658448
rect 615980 658438 616008 664902
rect 615968 658432 616020 658438
rect 615968 658374 616020 658380
rect 616716 652386 616744 676258
rect 617808 669380 617860 669386
rect 617808 669322 617860 669328
rect 616980 668768 617032 668774
rect 616980 668710 617032 668716
rect 616796 661900 616848 661906
rect 616796 661842 616848 661848
rect 616704 652380 616756 652386
rect 616704 652322 616756 652328
rect 615692 651836 615744 651842
rect 616808 651813 616836 661842
rect 616992 659118 617020 668710
rect 616980 659112 617032 659118
rect 616980 659054 617032 659060
rect 615692 651778 615744 651784
rect 616794 651804 616850 651813
rect 616794 651739 616850 651748
rect 615600 651088 615652 651094
rect 615600 651030 615652 651036
rect 615600 650816 615652 650822
rect 615600 650758 615652 650764
rect 615612 650550 615640 650758
rect 615600 650544 615652 650550
rect 615600 650486 615652 650492
rect 617820 649530 617848 669322
rect 617912 664830 617940 684078
rect 618912 667680 618964 667686
rect 618912 667622 618964 667628
rect 617900 664824 617952 664830
rect 617900 664766 617952 664772
rect 618268 659520 618320 659526
rect 618268 659462 618320 659468
rect 618280 654018 618308 659462
rect 618268 654012 618320 654018
rect 618268 653954 618320 653960
rect 617900 653944 617952 653950
rect 617900 653886 617952 653892
rect 617808 649524 617860 649530
rect 617808 649466 617860 649472
rect 615508 648776 615560 648782
rect 615508 648718 615560 648724
rect 617912 646917 617940 653886
rect 618924 648442 618952 667622
rect 619096 662920 619148 662926
rect 619096 662862 619148 662868
rect 619004 657276 619056 657282
rect 619004 657218 619056 657224
rect 619016 650890 619044 657218
rect 619108 651978 619136 662862
rect 619372 661356 619424 661362
rect 619372 661298 619424 661304
rect 619280 654556 619332 654562
rect 619280 654498 619332 654504
rect 619188 652380 619240 652386
rect 619188 652322 619240 652328
rect 619096 651972 619148 651978
rect 619096 651914 619148 651920
rect 619004 650884 619056 650890
rect 619004 650826 619056 650832
rect 619004 650408 619056 650414
rect 619004 650350 619056 650356
rect 618912 648436 618964 648442
rect 618912 648378 618964 648384
rect 402066 646908 402122 646917
rect 393432 646866 393552 646894
rect 398216 646866 398336 646894
rect 345486 646843 345542 646852
rect 402066 646843 402122 646852
rect 403078 646908 403134 646917
rect 403078 646843 403134 646852
rect 474286 646908 474342 646917
rect 474286 646843 474342 646852
rect 475022 646908 475078 646917
rect 475022 646843 475078 646852
rect 512466 646908 512522 646917
rect 512466 646843 512522 646852
rect 513294 646908 513350 646917
rect 513294 646843 513350 646852
rect 536754 646908 536810 646917
rect 536754 646843 536810 646852
rect 537398 646908 537454 646917
rect 537398 646843 537454 646852
rect 541170 646908 541226 646917
rect 541170 646843 541226 646852
rect 542182 646908 542238 646917
rect 542182 646843 542238 646852
rect 569874 646908 569930 646917
rect 569874 646843 569930 646852
rect 570886 646908 570942 646917
rect 570886 646843 570942 646852
rect 584226 646908 584282 646917
rect 584226 646843 584282 646852
rect 585238 646908 585294 646917
rect 585238 646843 585294 646852
rect 598578 646908 598634 646917
rect 598578 646843 598634 646852
rect 599590 646908 599646 646917
rect 612930 646908 612986 646917
rect 609080 646878 609200 646894
rect 599590 646843 599646 646852
rect 609068 646872 609200 646878
rect 609120 646866 609200 646872
rect 612930 646843 612986 646852
rect 613942 646908 613998 646917
rect 613942 646843 613998 646852
rect 617898 646908 617954 646917
rect 617898 646843 617954 646852
rect 618726 646908 618782 646917
rect 618726 646843 618782 646852
rect 609068 646814 609120 646820
rect 268668 646804 268720 646810
rect 268668 646746 268720 646752
rect 273636 646804 273688 646810
rect 273636 646746 273688 646752
rect 297832 646804 297884 646810
rect 297832 646746 297884 646752
rect 311908 646804 311960 646810
rect 311908 646746 311960 646752
rect 619016 414658 619044 650350
rect 619096 649592 619148 649598
rect 619096 649534 619148 649540
rect 619108 624574 619136 649534
rect 619096 624568 619148 624574
rect 619096 624510 619148 624516
rect 619094 624468 619150 624477
rect 619094 624403 619150 624412
rect 619108 621349 619136 624403
rect 619094 621340 619150 621349
rect 619094 621275 619150 621284
rect 619096 621236 619148 621242
rect 619096 621178 619148 621184
rect 619108 619270 619136 621178
rect 619096 619264 619148 619270
rect 619096 619206 619148 619212
rect 619096 617428 619148 617434
rect 619096 617370 619148 617376
rect 619108 613082 619136 617370
rect 619096 613076 619148 613082
rect 619096 613018 619148 613024
rect 619096 612940 619148 612946
rect 619096 612882 619148 612888
rect 619108 611829 619136 612882
rect 619094 611820 619150 611829
rect 619094 611755 619150 611764
rect 619094 611684 619150 611693
rect 619094 611619 619150 611628
rect 619108 610741 619136 611619
rect 619094 610732 619150 610741
rect 619094 610667 619150 610676
rect 619096 610628 619148 610634
rect 619096 610570 619148 610576
rect 619108 554738 619136 610570
rect 619096 554732 619148 554738
rect 619096 554674 619148 554680
rect 619094 551300 619150 551309
rect 619094 551235 619150 551244
rect 619108 545286 619136 551235
rect 619096 545280 619148 545286
rect 619096 545222 619148 545228
rect 619096 543580 619148 543586
rect 619096 543522 619148 543528
rect 619108 519893 619136 543522
rect 619200 526965 619228 652322
rect 619292 583541 619320 654498
rect 619384 650822 619412 661298
rect 619464 654012 619516 654018
rect 619464 653954 619516 653960
rect 619372 650816 619424 650822
rect 619372 650758 619424 650764
rect 619372 647008 619424 647014
rect 619372 646950 619424 646956
rect 619384 605550 619412 646950
rect 619476 613218 619504 653954
rect 619464 613212 619516 613218
rect 619464 613154 619516 613160
rect 619464 613076 619516 613082
rect 619464 613018 619516 613024
rect 619476 610634 619504 613018
rect 619464 610628 619516 610634
rect 619464 610570 619516 610576
rect 619384 605522 619504 605550
rect 619370 605428 619426 605437
rect 619370 605363 619426 605372
rect 619384 603941 619412 605363
rect 619476 604213 619504 605522
rect 619462 604204 619518 604213
rect 619462 604139 619518 604148
rect 619370 603932 619426 603941
rect 619370 603867 619426 603876
rect 619370 583804 619426 583813
rect 619370 583739 619426 583748
rect 619278 583532 619334 583541
rect 619278 583467 619334 583476
rect 619278 575372 619334 575381
rect 619278 575307 619334 575316
rect 619292 568474 619320 575307
rect 619384 571981 619412 583739
rect 619370 571972 619426 571981
rect 619370 571907 619426 571916
rect 619280 568468 619332 568474
rect 619280 568410 619332 568416
rect 619280 554732 619332 554738
rect 619280 554674 619332 554680
rect 619292 543586 619320 554674
rect 619372 545280 619424 545286
rect 619372 545222 619424 545228
rect 619280 543580 619332 543586
rect 619280 543522 619332 543528
rect 619278 542052 619334 542061
rect 619384 542038 619412 545222
rect 619334 542010 619412 542038
rect 619278 541987 619334 541996
rect 619186 526956 619242 526965
rect 619186 526891 619242 526900
rect 619094 519884 619150 519893
rect 619094 519819 619150 519828
rect 619464 506248 619516 506254
rect 619464 506190 619516 506196
rect 619476 504933 619504 506190
rect 619462 504924 619518 504933
rect 619462 504859 619518 504868
rect 619094 490236 619150 490245
rect 619094 490171 619150 490180
rect 619004 414652 619056 414658
rect 619004 414594 619056 414600
rect 257444 280556 257496 280562
rect 617164 280556 617216 280562
rect 257496 280504 257760 280510
rect 257444 280498 257760 280504
rect 257456 280482 257760 280498
rect 262240 280494 262544 280510
rect 607608 280494 607728 280510
rect 617216 280504 617296 280510
rect 617164 280498 617296 280504
rect 262228 280488 262544 280494
rect 262280 280482 262544 280488
rect 607596 280488 607728 280494
rect 262228 280430 262280 280436
rect 607648 280482 607728 280488
rect 617176 280482 617296 280498
rect 607596 280430 607648 280436
rect 362876 280420 362928 280426
rect 271900 280346 272112 280374
rect 271900 280290 271928 280346
rect 271888 280284 271940 280290
rect 271888 280226 271940 280232
rect 276868 279717 276896 280374
rect 276854 279708 276910 279717
rect 276854 279643 276910 279652
rect 252844 278380 252896 278386
rect 252844 278322 252896 278328
rect 281658 277962 281686 280378
rect 286436 279542 286464 280374
rect 286424 279536 286476 279542
rect 286424 279478 286476 279484
rect 300788 278386 300816 280374
rect 310356 280086 310384 280374
rect 310344 280080 310396 280086
rect 310344 280022 310396 280028
rect 315140 278454 315168 280374
rect 315128 278448 315180 278454
rect 315128 278390 315180 278396
rect 300776 278380 300828 278386
rect 300776 278322 300828 278328
rect 281639 277909 281645 277962
rect 281697 277909 281703 277962
rect 324708 264242 324736 280374
rect 339060 265330 339088 280374
rect 344028 279542 344056 280374
rect 588276 280420 588328 280426
rect 362928 280368 363192 280374
rect 362876 280362 363192 280368
rect 362888 280346 363192 280362
rect 360576 280284 360628 280290
rect 360576 280226 360628 280232
rect 344016 279536 344068 279542
rect 344016 279478 344068 279484
rect 360588 278522 360616 280226
rect 367948 279950 367976 280374
rect 367936 279944 367988 279950
rect 367936 279886 367988 279892
rect 377516 279474 377544 280374
rect 377504 279468 377556 279474
rect 377504 279410 377556 279416
rect 382300 278658 382328 280374
rect 387084 279610 387112 280374
rect 387072 279604 387124 279610
rect 387072 279546 387124 279552
rect 382288 278652 382340 278658
rect 382288 278594 382340 278600
rect 360576 278516 360628 278522
rect 360576 278458 360628 278464
rect 339048 265324 339100 265330
rect 339048 265266 339100 265272
rect 324696 264236 324748 264242
rect 324696 264178 324748 264184
rect 391868 263086 391896 280374
rect 396652 279853 396680 280374
rect 396638 279844 396694 279853
rect 396638 279779 396694 279788
rect 401436 278658 401464 280374
rect 401424 278652 401476 278658
rect 401424 278594 401476 278600
rect 411004 278590 411032 280374
rect 415788 279678 415816 280374
rect 420296 280358 420600 280374
rect 420284 280352 420600 280358
rect 420336 280346 420600 280352
rect 420284 280294 420336 280300
rect 430324 279746 430352 280374
rect 435016 280358 435136 280374
rect 435004 280352 435136 280358
rect 435056 280346 435136 280352
rect 435004 280294 435056 280300
rect 430312 279740 430364 279746
rect 430312 279682 430364 279688
rect 415776 279672 415828 279678
rect 415776 279614 415828 279620
rect 410992 278584 411044 278590
rect 410992 278526 411044 278532
rect 449479 278072 449508 280379
rect 454244 279746 454272 280374
rect 463812 279882 463840 280374
rect 463800 279876 463852 279882
rect 463800 279818 463852 279824
rect 473380 279814 473408 280374
rect 473368 279808 473420 279814
rect 473368 279750 473420 279756
rect 454232 279740 454284 279746
rect 454232 279682 454284 279688
rect 478164 279037 478192 280374
rect 487732 279882 487760 280374
rect 487720 279876 487772 279882
rect 487720 279818 487772 279824
rect 478150 279028 478206 279037
rect 478150 278963 478206 278972
rect 492516 278726 492544 280374
rect 497300 279814 497328 280374
rect 497288 279808 497340 279814
rect 497288 279750 497340 279756
rect 502504 278794 502532 280374
rect 506868 278794 506896 280374
rect 511652 280018 511680 280374
rect 511640 280012 511692 280018
rect 511640 279954 511692 279960
rect 516620 278862 516648 280374
rect 526188 278862 526216 280374
rect 535756 278930 535784 280374
rect 535744 278924 535796 278930
rect 535744 278866 535796 278872
rect 516608 278856 516660 278862
rect 516608 278798 516660 278804
rect 526176 278856 526228 278862
rect 526176 278798 526228 278804
rect 502492 278788 502544 278794
rect 502492 278730 502544 278736
rect 506856 278788 506908 278794
rect 506856 278730 506908 278736
rect 492504 278720 492556 278726
rect 492504 278662 492556 278668
rect 540540 278318 540568 280374
rect 549924 280346 550136 280374
rect 549924 280290 549952 280346
rect 549912 280284 549964 280290
rect 549912 280226 549964 280232
rect 554892 280018 554920 280374
rect 554880 280012 554932 280018
rect 554880 279954 554932 279960
rect 564460 278998 564488 280374
rect 569244 278998 569272 280374
rect 573936 280346 574056 280374
rect 573936 280290 573964 280346
rect 573924 280284 573976 280290
rect 573924 280226 573976 280232
rect 564448 278992 564500 278998
rect 564448 278934 564500 278940
rect 569232 278992 569284 278998
rect 569232 278934 569284 278940
rect 578812 278726 578840 280374
rect 578800 278720 578852 278726
rect 578800 278662 578852 278668
rect 540528 278312 540580 278318
rect 540528 278254 540580 278260
rect 449461 278020 449468 278072
rect 449520 278020 449526 278072
rect 576960 266412 577012 266418
rect 576960 266354 577012 266360
rect 384312 263080 384364 263086
rect 384312 263022 384364 263028
rect 391856 263080 391908 263086
rect 391856 263022 391908 263028
rect 252016 261992 252068 261998
rect 252016 261934 252068 261940
rect 382826 259748 382878 259754
rect 384324 259745 384352 263022
rect 565920 262060 565972 262066
rect 565920 262002 565972 262008
rect 522220 260020 522272 260026
rect 522220 259962 522272 259968
rect 554788 260020 554840 260026
rect 554788 259962 554840 259968
rect 397560 259952 397612 259958
rect 397560 259894 397612 259900
rect 423872 259952 423924 259958
rect 423872 259894 423924 259900
rect 424608 259952 424660 259958
rect 424608 259894 424660 259900
rect 456992 259952 457044 259958
rect 456992 259894 457044 259900
rect 489560 259952 489612 259958
rect 489560 259894 489612 259900
rect 395076 259884 395128 259890
rect 395076 259826 395128 259832
rect 397284 259884 397336 259890
rect 397284 259826 397336 259832
rect 384981 259768 385033 259774
rect 382826 259690 382878 259696
rect 384310 259736 384366 259745
rect 247416 259612 247468 259618
rect 247416 259554 247468 259560
rect 382838 259470 382866 259690
rect 384310 259671 384366 259680
rect 384494 259736 384550 259745
rect 389299 259768 389351 259774
rect 388377 259748 388429 259754
rect 384981 259710 385033 259716
rect 388375 259716 388377 259725
rect 388429 259716 388431 259725
rect 384494 259671 384550 259680
rect 384508 259570 384536 259671
rect 384496 259564 384548 259570
rect 384496 259506 384548 259512
rect 384993 259490 385021 259710
rect 395088 259725 395116 259826
rect 389299 259710 389351 259716
rect 392196 259716 392252 259725
rect 388375 259651 388431 259660
rect 388389 259470 388417 259651
rect 389311 259586 389339 259710
rect 391985 259680 392037 259686
rect 392196 259651 392252 259660
rect 392636 259716 392692 259725
rect 392636 259651 392692 259660
rect 393026 259716 393082 259725
rect 393026 259651 393082 259660
rect 393875 259716 393931 259725
rect 393875 259651 393931 259660
rect 395074 259716 395130 259725
rect 395074 259651 395130 259660
rect 391985 259622 392037 259628
rect 389200 259570 389339 259586
rect 389188 259564 389339 259570
rect 389240 259558 389339 259564
rect 389188 259506 389240 259512
rect 389311 259470 389339 259558
rect 391270 259570 391436 259586
rect 391270 259564 391448 259570
rect 391270 259558 391396 259564
rect 391270 259490 391298 259558
rect 391396 259506 391448 259512
rect 391997 259470 392025 259622
rect 392210 259470 392238 259651
rect 392650 259470 392678 259651
rect 393040 259470 393068 259651
rect 393889 259470 393917 259651
rect 395088 259470 395116 259651
rect 397296 259576 397324 259826
rect 395797 259556 395849 259562
rect 395797 259498 395849 259504
rect 397134 259548 397324 259576
rect 397572 259562 397600 259894
rect 415408 259884 415460 259890
rect 415408 259826 415460 259832
rect 423688 259884 423740 259890
rect 423688 259826 423740 259832
rect 414856 259816 414908 259822
rect 397836 259760 397888 259766
rect 414856 259758 414908 259764
rect 414868 259725 414896 259758
rect 415420 259725 415448 259826
rect 418068 259816 418120 259822
rect 418068 259758 418120 259764
rect 421894 259798 421946 259804
rect 397836 259702 397888 259708
rect 414854 259716 414910 259725
rect 397848 259562 397876 259702
rect 415420 259716 415480 259725
rect 415420 259674 415424 259716
rect 414854 259651 414910 259660
rect 415424 259651 415480 259660
rect 417579 259716 417635 259725
rect 417579 259651 417635 259660
rect 397560 259556 397612 259562
rect 395809 259482 395837 259498
rect 397134 259470 397162 259548
rect 397279 259470 397307 259548
rect 397560 259498 397612 259504
rect 397676 259556 397728 259562
rect 397676 259498 397728 259504
rect 397836 259556 397888 259562
rect 397836 259498 397888 259504
rect 397688 259470 397716 259498
rect 414868 259346 414896 259651
rect 415438 259470 415466 259651
rect 417593 259470 417621 259651
rect 418080 259637 418108 259758
rect 421894 259740 421946 259746
rect 420972 259716 421028 259725
rect 420972 259651 421028 259660
rect 418080 259609 418500 259637
rect 418448 259604 418500 259609
rect 418448 259546 418500 259552
rect 420986 259470 421014 259651
rect 421906 259586 421934 259740
rect 423700 259686 423728 259826
rect 423884 259686 423912 259894
rect 423688 259680 423740 259686
rect 423688 259622 423740 259628
rect 423856 259680 423912 259686
rect 423908 259640 423912 259680
rect 423856 259622 423908 259628
rect 421768 259570 421934 259586
rect 421756 259564 421934 259570
rect 421808 259538 421934 259564
rect 421756 259506 421808 259512
rect 421906 259470 421934 259538
rect 423868 259470 423896 259622
rect 424620 259566 424648 259894
rect 454416 259836 454468 259842
rect 426448 259816 426500 259822
rect 426448 259758 426500 259764
rect 427736 259816 427788 259822
rect 427736 259758 427788 259764
rect 429852 259816 429904 259822
rect 454416 259778 454468 259784
rect 429852 259758 429904 259764
rect 426460 259725 426488 259758
rect 424790 259716 424846 259725
rect 424790 259651 424846 259660
rect 425248 259716 425304 259725
rect 425248 259651 425304 259660
rect 425618 259716 425674 259725
rect 425618 259651 425674 259660
rect 426446 259716 426502 259725
rect 426446 259651 426502 259660
rect 424597 259538 424648 259566
rect 424597 259470 424625 259538
rect 424804 259470 424832 259651
rect 425262 259470 425290 259651
rect 425632 259470 425660 259651
rect 426460 259566 426488 259651
rect 427748 259566 427776 259758
rect 429864 259702 429892 259758
rect 430276 259748 430328 259754
rect 428397 259680 428449 259686
rect 429864 259674 429907 259702
rect 447838 259748 447890 259754
rect 430276 259690 430328 259696
rect 446318 259716 446374 259725
rect 428397 259622 428449 259628
rect 426460 259538 426517 259566
rect 426489 259470 426517 259538
rect 427702 259538 427776 259566
rect 427702 259470 427730 259538
rect 428409 259470 428437 259622
rect 429879 259566 429907 259674
rect 429734 259538 429907 259566
rect 429734 259470 429762 259538
rect 429879 259470 429907 259538
rect 430288 259566 430316 259690
rect 447838 259690 447890 259696
rect 449981 259748 450033 259754
rect 453377 259748 453429 259754
rect 449981 259690 450033 259696
rect 451010 259716 451066 259725
rect 446318 259651 446374 259660
rect 430288 259550 431244 259566
rect 446332 259550 446360 259651
rect 430288 259544 431256 259550
rect 430288 259538 431204 259544
rect 430288 259470 430316 259538
rect 431204 259486 431256 259492
rect 446320 259544 446372 259550
rect 446320 259486 446372 259492
rect 447850 259470 447878 259690
rect 449993 259470 450021 259690
rect 453377 259690 453429 259696
rect 451010 259651 451066 259660
rect 451024 259571 451052 259651
rect 451012 259565 451064 259571
rect 451012 259507 451064 259513
rect 453389 259470 453417 259690
rect 454152 259660 454339 259688
rect 454152 259570 454180 259660
rect 454311 259626 454339 259660
rect 454428 259649 454456 259778
rect 456256 259680 456308 259686
rect 454414 259640 454470 259649
rect 454311 259598 454414 259626
rect 454140 259564 454192 259570
rect 454140 259506 454192 259512
rect 454311 259490 454339 259598
rect 456256 259622 456308 259628
rect 454414 259575 454470 259584
rect 456268 259470 456296 259622
rect 457004 259470 457032 259894
rect 457176 259816 457228 259822
rect 457176 259758 457228 259764
rect 462696 259816 462748 259822
rect 462696 259758 462748 259764
rect 480268 259816 480320 259822
rect 480268 259758 480320 259764
rect 483472 259820 483524 259826
rect 483472 259762 483524 259768
rect 457188 259566 457216 259758
rect 457650 259748 457702 259754
rect 457650 259690 457702 259696
rect 458028 259748 458080 259754
rect 458028 259690 458080 259696
rect 458878 259748 458930 259754
rect 458878 259690 458930 259696
rect 460086 259748 460138 259754
rect 460086 259690 460138 259696
rect 462267 259748 462319 259754
rect 462267 259690 462319 259696
rect 457188 259538 457238 259566
rect 457210 259470 457238 259538
rect 457662 259470 457690 259690
rect 458040 259470 458068 259690
rect 458890 259470 458918 259690
rect 460098 259470 460126 259690
rect 460797 259680 460849 259686
rect 460797 259622 460849 259628
rect 460809 259470 460837 259622
rect 462279 259566 462307 259690
rect 462708 259566 462736 259758
rect 480280 259725 480308 259758
rect 480426 259748 480478 259754
rect 480266 259716 480322 259725
rect 482581 259748 482633 259754
rect 480426 259690 480478 259696
rect 482579 259716 482581 259725
rect 482633 259716 482635 259725
rect 480266 259651 480322 259660
rect 462134 259538 462307 259566
rect 462134 259470 462162 259538
rect 462279 259470 462307 259538
rect 462688 259538 462736 259566
rect 462688 259470 462716 259538
rect 480438 259470 480466 259690
rect 482579 259651 482635 259660
rect 482593 259470 482621 259651
rect 483476 259570 483513 259762
rect 486899 259748 486951 259754
rect 485970 259716 486026 259725
rect 486899 259690 486951 259696
rect 485970 259651 486026 259660
rect 483463 259564 483515 259570
rect 483463 259506 483515 259512
rect 485984 259470 486012 259651
rect 486911 259470 486939 259690
rect 488856 259680 488908 259686
rect 488856 259622 488908 259628
rect 488868 259470 488896 259622
rect 489572 259566 489600 259894
rect 513020 259884 513072 259890
rect 513020 259826 513072 259832
rect 494712 259816 494764 259822
rect 494712 259758 494764 259764
rect 512836 259816 512888 259822
rect 512836 259758 512888 259764
rect 494724 259725 494752 259758
rect 495276 259748 495328 259754
rect 489788 259716 489844 259725
rect 489788 259651 489844 259660
rect 490248 259716 490304 259725
rect 490248 259651 490304 259660
rect 490616 259716 490672 259725
rect 490616 259651 490672 259660
rect 491475 259716 491531 259725
rect 491475 259651 491531 259660
rect 492684 259716 492740 259725
rect 494710 259716 494766 259725
rect 492684 259651 492740 259660
rect 493397 259680 493449 259686
rect 489572 259538 489625 259566
rect 489597 259470 489625 259538
rect 489802 259470 489830 259651
rect 490262 259470 490290 259651
rect 490630 259470 490658 259651
rect 491489 259470 491517 259651
rect 492698 259470 492726 259651
rect 512848 259725 512876 259758
rect 513032 259754 513060 259826
rect 518540 259816 518592 259822
rect 516148 259768 516200 259774
rect 513020 259748 513072 259754
rect 495276 259690 495328 259696
rect 512834 259716 512890 259725
rect 494710 259651 494766 259660
rect 493397 259622 493449 259628
rect 493409 259470 493437 259622
rect 494724 259566 494752 259651
rect 494724 259538 494907 259566
rect 494724 259470 494752 259538
rect 494879 259470 494907 259538
rect 495288 259470 495316 259690
rect 513020 259690 513072 259696
rect 515182 259748 515234 259754
rect 515182 259690 515234 259696
rect 516146 259736 516148 259745
rect 518540 259758 518592 259764
rect 516200 259736 516202 259745
rect 518552 259725 518580 259758
rect 519506 259748 519558 259754
rect 512834 259651 512890 259660
rect 513032 259470 513060 259690
rect 515194 259470 515222 259690
rect 516146 259671 516202 259680
rect 518538 259716 518594 259725
rect 516160 259570 516188 259671
rect 519506 259690 519558 259696
rect 518538 259651 518594 259660
rect 516148 259564 516200 259570
rect 518552 259566 518580 259651
rect 518552 259538 518617 259566
rect 516148 259506 516200 259512
rect 518589 259470 518617 259538
rect 519518 259470 519546 259690
rect 521456 259680 521508 259686
rect 521456 259622 521508 259628
rect 521468 259470 521496 259622
rect 522232 259566 522260 259962
rect 545588 259952 545640 259958
rect 545588 259894 545640 259900
rect 548440 259952 548492 259958
rect 548440 259894 548492 259900
rect 522404 259884 522456 259890
rect 522404 259826 522456 259832
rect 522864 259884 522916 259890
rect 522864 259826 522916 259832
rect 523232 259884 523284 259890
rect 523232 259826 523284 259832
rect 524060 259884 524112 259890
rect 524060 259826 524112 259832
rect 525256 259884 525308 259890
rect 525256 259826 525308 259832
rect 527464 259884 527516 259890
rect 527464 259826 527516 259832
rect 545312 259884 545364 259890
rect 545312 259826 545364 259832
rect 522416 259725 522444 259826
rect 522402 259716 522458 259725
rect 522402 259651 522458 259660
rect 522197 259538 522260 259566
rect 522197 259470 522225 259538
rect 522416 259470 522444 259651
rect 522876 259566 522904 259826
rect 522862 259538 522904 259566
rect 522862 259470 522890 259538
rect 523244 259470 523272 259826
rect 524072 259566 524100 259826
rect 525268 259702 525296 259826
rect 525268 259674 525326 259702
rect 524072 259538 524117 259566
rect 524089 259470 524117 259538
rect 525298 259470 525326 259674
rect 525992 259680 526044 259686
rect 525992 259622 526044 259628
rect 526004 259470 526032 259622
rect 527476 259566 527504 259826
rect 527878 259748 527930 259754
rect 527878 259690 527930 259696
rect 545036 259748 545088 259754
rect 545324 259702 545352 259826
rect 545600 259822 545628 259894
rect 545588 259816 545640 259822
rect 545588 259758 545640 259764
rect 545036 259690 545088 259696
rect 527338 259538 527504 259566
rect 527338 259470 527366 259538
rect 527476 259470 527504 259538
rect 527890 259470 527918 259690
rect 545048 259653 545076 259690
rect 545223 259674 545352 259702
rect 545600 259702 545628 259758
rect 547781 259748 547833 259754
rect 545600 259674 545674 259702
rect 547781 259690 547833 259696
rect 545034 259644 545090 259653
rect 545034 259579 545090 259588
rect 545223 259470 545251 259674
rect 545646 259470 545674 259674
rect 547793 259470 547821 259690
rect 548452 259570 548480 259894
rect 551200 259884 551252 259890
rect 551200 259826 551252 259832
rect 551212 259725 551240 259826
rect 553500 259816 553552 259822
rect 553482 259764 553500 259804
rect 553482 259758 553552 259764
rect 551175 259716 551240 259725
rect 551231 259674 551240 259716
rect 552099 259748 552151 259754
rect 552099 259690 552151 259696
rect 551175 259651 551231 259660
rect 548440 259564 548492 259570
rect 548440 259506 548492 259512
rect 551189 259470 551217 259651
rect 552111 259470 552139 259690
rect 553482 259470 553510 259758
rect 554052 259680 554104 259686
rect 554052 259622 554104 259628
rect 554064 259470 554092 259622
rect 554800 259470 554828 259962
rect 558652 259952 558704 259958
rect 558652 259894 558704 259900
rect 555432 259884 555484 259890
rect 555432 259826 555484 259832
rect 554996 259716 555052 259725
rect 555444 259702 555472 259826
rect 558664 259822 558692 259894
rect 558652 259816 558704 259822
rect 558652 259758 558704 259764
rect 556677 259748 556729 259754
rect 555444 259674 555490 259702
rect 556677 259690 556729 259696
rect 554996 259651 554998 259660
rect 555050 259651 555052 259660
rect 554998 259622 555050 259628
rect 555010 259470 555038 259622
rect 555462 259470 555490 259674
rect 555828 259680 555880 259686
rect 555828 259622 555880 259628
rect 555840 259470 555868 259622
rect 556689 259470 556717 259690
rect 557886 259680 557938 259686
rect 557886 259622 557938 259628
rect 557898 259470 557926 259622
rect 558664 259566 558692 259758
rect 565932 259754 565960 262002
rect 576972 259754 577000 266354
rect 577604 262128 577656 262134
rect 577604 262070 577656 262076
rect 565920 259748 565972 259754
rect 565920 259690 565972 259696
rect 576960 259748 577012 259754
rect 576960 259690 577012 259696
rect 560067 259680 560119 259686
rect 560067 259622 560119 259628
rect 560476 259680 560528 259686
rect 560476 259622 560528 259628
rect 560079 259566 560107 259622
rect 558618 259538 558692 259566
rect 559934 259538 560107 259566
rect 558618 259470 558646 259538
rect 559934 259470 559962 259538
rect 560079 259470 560107 259538
rect 560488 259470 560516 259622
rect 577616 259513 577644 262070
rect 583596 260910 583624 280374
rect 588328 280368 588408 280374
rect 588276 280362 588408 280368
rect 588288 280346 588408 280362
rect 612484 280086 612512 280374
rect 612472 280080 612524 280086
rect 612472 280022 612524 280028
rect 619108 276346 619136 490171
rect 619188 414652 619240 414658
rect 619188 414594 619240 414600
rect 619200 406469 619228 414594
rect 619186 406460 619242 406469
rect 619186 406395 619242 406404
rect 619568 278794 619596 728958
rect 622696 728886 622724 729514
rect 623064 729486 623121 729514
rect 623064 729446 623092 729486
rect 623238 729446 623266 729514
rect 623064 729430 623266 729446
rect 624432 729482 624484 729488
rect 624551 729484 624579 729515
rect 624536 729470 624579 729484
rect 624484 729456 624579 729470
rect 624484 729442 624564 729456
rect 623064 729424 623278 729430
rect 624432 729424 624484 729430
rect 623064 729418 623226 729424
rect 622684 728880 622736 728886
rect 622684 728822 622736 728828
rect 623064 728818 623092 729418
rect 623226 729366 623278 729372
rect 623238 729335 623266 729366
rect 623052 728812 623104 728818
rect 623052 728754 623104 728760
rect 624536 728750 624564 729442
rect 625274 729430 625302 729514
rect 626483 729430 626511 729514
rect 627342 729430 627370 729514
rect 627710 729430 627738 729514
rect 628170 729430 628198 729514
rect 628375 729446 628403 729514
rect 629104 729492 629440 729514
rect 629104 729486 629216 729492
rect 625262 729424 625314 729430
rect 625262 729366 625314 729372
rect 626471 729424 626523 729430
rect 626471 729366 626523 729372
rect 627330 729424 627382 729430
rect 627330 729366 627382 729372
rect 627698 729424 627750 729430
rect 627698 729366 627750 729372
rect 628158 729424 628210 729430
rect 628375 729418 628428 729446
rect 629268 729486 629440 729492
rect 629216 729434 629268 729440
rect 628158 729366 628210 729372
rect 628400 728750 628428 729418
rect 629228 729403 629256 729434
rect 624524 728744 624576 728750
rect 624524 728686 624576 728692
rect 628388 728744 628440 728750
rect 628388 728686 628440 728692
rect 621764 728608 621816 728614
rect 621764 728550 621816 728556
rect 619648 695356 619700 695362
rect 619648 695298 619700 695304
rect 619660 278998 619688 695298
rect 620016 664824 620068 664830
rect 620016 664766 620068 664772
rect 620028 653678 620056 664766
rect 621304 663872 621356 663878
rect 621304 663814 621356 663820
rect 620108 658500 620160 658506
rect 620108 658442 620160 658448
rect 620120 654970 620148 658442
rect 621028 658432 621080 658438
rect 621028 658374 621080 658380
rect 620108 654964 620160 654970
rect 620108 654906 620160 654912
rect 620016 653672 620068 653678
rect 620016 653614 620068 653620
rect 620844 651836 620896 651842
rect 620844 651778 620896 651784
rect 619740 650612 619792 650618
rect 619740 650554 619792 650560
rect 619648 278992 619700 278998
rect 619648 278934 619700 278940
rect 619752 278862 619780 650554
rect 619924 648776 619976 648782
rect 619924 648718 619976 648724
rect 619832 647348 619884 647354
rect 619832 647290 619884 647296
rect 619844 280494 619872 647290
rect 619936 292501 619964 648718
rect 620660 648436 620712 648442
rect 620660 648378 620712 648384
rect 620014 636708 620070 636717
rect 620014 636643 620070 636652
rect 620028 632093 620056 636643
rect 620014 632084 620070 632093
rect 620014 632019 620070 632028
rect 620016 619264 620068 619270
rect 620016 619206 620068 619212
rect 620028 617434 620056 619206
rect 620016 617428 620068 617434
rect 620016 617370 620068 617376
rect 620672 617230 620700 648378
rect 620752 647212 620804 647218
rect 620752 647154 620804 647160
rect 620016 617224 620068 617230
rect 620016 617166 620068 617172
rect 620660 617224 620712 617230
rect 620660 617166 620712 617172
rect 620028 597141 620056 617166
rect 620014 597132 620070 597141
rect 620014 597067 620070 597076
rect 620014 547628 620070 547637
rect 620014 547563 620070 547572
rect 620028 547462 620056 547563
rect 620016 547456 620068 547462
rect 620016 547398 620068 547404
rect 620016 535284 620068 535290
rect 620016 535226 620068 535232
rect 619922 292492 619978 292501
rect 619922 292427 619978 292436
rect 619832 280488 619884 280494
rect 619832 280430 619884 280436
rect 620028 279542 620056 535226
rect 620108 532564 620160 532570
rect 620108 532506 620160 532512
rect 620120 469573 620148 532506
rect 620106 469564 620162 469573
rect 620106 469499 620162 469508
rect 620200 464088 620252 464094
rect 620200 464030 620252 464036
rect 620212 441285 620240 464030
rect 620198 441276 620254 441285
rect 620198 441211 620254 441220
rect 620108 425328 620160 425334
rect 620108 425270 620160 425276
rect 620120 313717 620148 425270
rect 620200 425056 620252 425062
rect 620200 424998 620252 425004
rect 620212 420069 620240 424998
rect 620292 423220 620344 423226
rect 620292 423162 620344 423168
rect 620198 420060 620254 420069
rect 620198 419995 620254 420004
rect 620304 416026 620332 423162
rect 620212 415998 620332 416026
rect 620212 370293 620240 415998
rect 620198 370284 620254 370293
rect 620198 370219 620254 370228
rect 620106 313708 620162 313717
rect 620106 313643 620162 313652
rect 620016 279536 620068 279542
rect 620016 279478 620068 279484
rect 619740 278856 619792 278862
rect 619740 278798 619792 278804
rect 619556 278788 619608 278794
rect 619556 278730 619608 278736
rect 611184 276340 611236 276346
rect 611184 276282 611236 276288
rect 619096 276340 619148 276346
rect 619096 276282 619148 276288
rect 609712 274164 609764 274170
rect 609712 274106 609764 274112
rect 604560 264236 604612 264242
rect 604560 264178 604612 264184
rect 601984 263080 602036 263086
rect 601984 263022 602036 263028
rect 583584 260904 583636 260910
rect 583584 260846 583636 260852
rect 587356 260292 587408 260298
rect 587356 260234 587408 260240
rect 587368 260094 587396 260234
rect 590484 260156 590536 260162
rect 590484 260098 590536 260104
rect 592692 260156 592744 260162
rect 592692 260098 592744 260104
rect 587356 260088 587408 260094
rect 587356 260030 587408 260036
rect 586620 259952 586672 259958
rect 586620 259894 586672 259900
rect 578064 259884 578116 259890
rect 578064 259826 578116 259832
rect 580824 259884 580876 259890
rect 580824 259826 580876 259832
rect 577788 259816 577840 259822
rect 577840 259764 577851 259804
rect 577788 259758 577851 259764
rect 577602 259504 577658 259513
rect 577823 259470 577851 259758
rect 578076 259725 578104 259826
rect 580836 259725 580864 259826
rect 586068 259816 586120 259822
rect 584688 259798 584740 259804
rect 586068 259758 586120 259764
rect 584688 259740 584740 259746
rect 578062 259716 578118 259725
rect 580822 259716 580878 259725
rect 578062 259651 578118 259660
rect 578226 259680 578278 259686
rect 578226 259622 578278 259628
rect 580381 259680 580433 259686
rect 580822 259651 580878 259660
rect 583775 259716 583831 259725
rect 583775 259651 583777 259660
rect 580381 259622 580433 259628
rect 583829 259651 583831 259660
rect 584502 259716 584558 259725
rect 584502 259651 584558 259660
rect 583777 259622 583829 259628
rect 578238 259470 578266 259622
rect 580393 259566 580421 259622
rect 580608 259580 580648 259581
rect 580608 259574 580660 259580
rect 580393 259538 580608 259566
rect 580393 259470 580421 259538
rect 580608 259516 580660 259522
rect 583789 259470 583817 259622
rect 584516 259580 584544 259651
rect 584504 259574 584556 259580
rect 584504 259516 584556 259522
rect 584700 259470 584728 259740
rect 586080 259470 586108 259758
rect 586632 259754 586660 259894
rect 586620 259748 586672 259754
rect 586620 259690 586672 259696
rect 586632 259566 586660 259690
rect 587368 259566 587396 260030
rect 590496 259725 590524 260098
rect 591197 259748 591249 259754
rect 587584 259716 587640 259725
rect 587584 259651 587640 259660
rect 588044 259716 588100 259725
rect 588044 259651 588100 259660
rect 588426 259716 588482 259725
rect 588426 259651 588482 259660
rect 590482 259716 590538 259725
rect 591197 259690 591249 259696
rect 590482 259651 590538 259660
rect 586632 259538 586696 259566
rect 587368 259538 587425 259566
rect 586668 259470 586696 259538
rect 587397 259470 587425 259538
rect 587598 259470 587626 259651
rect 588058 259470 588086 259651
rect 588440 259470 588468 259651
rect 590496 259470 590524 259651
rect 591209 259470 591237 259690
rect 592704 259566 592732 260098
rect 601996 259890 602024 263022
rect 601984 259884 602036 259890
rect 601984 259826 602036 259832
rect 604572 259822 604600 264178
rect 609724 259997 609752 274106
rect 611196 263222 611224 276282
rect 620764 274170 620792 647154
rect 620856 334933 620884 651778
rect 620936 650680 620988 650686
rect 620936 650622 620988 650628
rect 620948 342005 620976 650622
rect 621040 384437 621068 658374
rect 621120 651972 621172 651978
rect 621120 651914 621172 651920
rect 621132 425062 621160 651914
rect 621212 649524 621264 649530
rect 621212 649466 621264 649472
rect 621224 427141 621252 649466
rect 621316 464094 621344 663814
rect 621488 659112 621540 659118
rect 621488 659054 621540 659060
rect 621500 654766 621528 659054
rect 621488 654760 621540 654766
rect 621488 654702 621540 654708
rect 621672 652788 621724 652794
rect 621672 652730 621724 652736
rect 621396 651088 621448 651094
rect 621396 651030 621448 651036
rect 621408 497861 621436 651030
rect 621488 632456 621540 632462
rect 621488 632398 621540 632404
rect 621500 632229 621528 632398
rect 621486 632220 621542 632229
rect 621486 632155 621542 632164
rect 621394 497852 621450 497861
rect 621394 497787 621450 497796
rect 621304 464088 621356 464094
rect 621304 464030 621356 464036
rect 621210 427132 621266 427141
rect 621210 427067 621266 427076
rect 621120 425056 621172 425062
rect 621120 424998 621172 425004
rect 621026 384428 621082 384437
rect 621026 384363 621082 384372
rect 620934 341996 620990 342005
rect 620934 341931 620990 341940
rect 620842 334924 620898 334933
rect 620842 334859 620898 334868
rect 621120 285452 621172 285458
rect 621120 285394 621172 285400
rect 621132 280358 621160 285394
rect 621120 280352 621172 280358
rect 621120 280294 621172 280300
rect 621684 278930 621712 652730
rect 621672 278924 621724 278930
rect 621672 278866 621724 278872
rect 621776 278658 621804 728550
rect 629412 728546 629440 729486
rect 631049 729464 631101 729552
rect 631049 729436 631188 729464
rect 631049 729435 631101 729436
rect 631160 728954 631188 729436
rect 631240 729424 631292 729430
rect 631240 729366 631292 729372
rect 631252 729333 631280 729366
rect 631988 729333 632016 729514
rect 635392 729430 635420 729514
rect 637534 729446 637562 729514
rect 637508 729430 637562 729446
rect 635380 729424 635432 729430
rect 635380 729366 635432 729372
rect 637496 729424 637562 729430
rect 637548 729418 637562 729424
rect 649885 729373 649916 729521
rect 637496 729366 637548 729372
rect 631238 729324 631294 729333
rect 631238 729259 631294 729268
rect 631974 729324 632030 729333
rect 631974 729259 632030 729268
rect 631148 728948 631200 728954
rect 631148 728890 631200 728896
rect 631988 728886 632016 729259
rect 637218 729052 637274 729061
rect 637218 728987 637274 728996
rect 631976 728880 632028 728886
rect 631976 728822 632028 728828
rect 629400 728540 629452 728546
rect 629400 728482 629452 728488
rect 625076 694540 625128 694546
rect 625076 694482 625128 694488
rect 624432 694268 624484 694274
rect 624432 694210 624484 694216
rect 624444 656126 624472 694210
rect 624432 656120 624484 656126
rect 624432 656062 624484 656068
rect 622132 654964 622184 654970
rect 622132 654906 622184 654912
rect 621856 650748 621908 650754
rect 621856 650690 621908 650696
rect 621764 278652 621816 278658
rect 621764 278594 621816 278600
rect 620752 274164 620804 274170
rect 620752 274106 620804 274112
rect 611736 265324 611788 265330
rect 611736 265266 611788 265272
rect 610264 263216 610316 263222
rect 610264 263158 610316 263164
rect 611184 263216 611236 263222
rect 611184 263158 611236 263164
rect 610276 260018 610304 263158
rect 610816 260156 610868 260162
rect 610816 260098 610868 260104
rect 610448 260088 610500 260094
rect 610448 260030 610500 260036
rect 610264 260012 610316 260018
rect 609710 259988 609766 259997
rect 610264 259954 610316 259960
rect 609710 259923 609766 259932
rect 604560 259816 604612 259822
rect 610460 259804 610488 260030
rect 604560 259758 604612 259764
rect 610423 259776 610488 259804
rect 610630 259852 610686 259861
rect 610630 259787 610686 259796
rect 593076 259680 593128 259686
rect 593076 259622 593128 259628
rect 592534 259538 592732 259566
rect 592534 259470 592562 259538
rect 592679 259470 592707 259538
rect 593088 259470 593116 259622
rect 610423 259470 610451 259776
rect 610644 259686 610672 259787
rect 610632 259680 610684 259686
rect 610632 259622 610684 259628
rect 610828 259566 610856 260098
rect 611748 260026 611776 265266
rect 621868 262066 621896 650690
rect 621948 650544 622000 650550
rect 621948 650486 622000 650492
rect 621960 280290 621988 650486
rect 622040 648368 622092 648374
rect 622040 648310 622092 648316
rect 622052 280426 622080 648310
rect 622144 320789 622172 654906
rect 623144 654760 623196 654766
rect 623144 654702 623196 654708
rect 622592 653672 622644 653678
rect 622592 653614 622644 653620
rect 622224 650884 622276 650890
rect 622224 650826 622276 650832
rect 622236 349077 622264 650826
rect 622408 650816 622460 650822
rect 622408 650758 622460 650764
rect 622316 647620 622368 647626
rect 622316 647562 622368 647568
rect 622328 412997 622356 647562
rect 622420 462501 622448 650758
rect 622500 650340 622552 650346
rect 622500 650282 622552 650288
rect 622512 532570 622540 650282
rect 622604 561781 622632 653614
rect 622960 652856 623012 652862
rect 622960 652798 623012 652804
rect 622868 650476 622920 650482
rect 622868 650418 622920 650424
rect 622590 561772 622646 561781
rect 622590 561707 622646 561716
rect 622500 532564 622552 532570
rect 622500 532506 622552 532512
rect 622406 462492 622462 462501
rect 622406 462427 622462 462436
rect 622314 412988 622370 412997
rect 622314 412923 622370 412932
rect 622222 349068 622278 349077
rect 622222 349003 622278 349012
rect 622130 320780 622186 320789
rect 622130 320715 622186 320724
rect 622040 280420 622092 280426
rect 622040 280362 622092 280368
rect 621948 280284 622000 280290
rect 621948 280226 622000 280232
rect 622880 262134 622908 650418
rect 622972 278726 623000 652798
rect 623052 649456 623104 649462
rect 623052 649398 623104 649404
rect 623064 285458 623092 649398
rect 623156 398853 623184 654702
rect 624432 648028 624484 648034
rect 624432 647970 624484 647976
rect 623236 647960 623288 647966
rect 623236 647902 623288 647908
rect 623248 434213 623276 647902
rect 623328 635176 623380 635182
rect 623328 635118 623380 635124
rect 623340 506254 623368 635118
rect 624444 611518 624472 647970
rect 624432 611512 624484 611518
rect 624432 611454 624484 611460
rect 624432 581388 624484 581394
rect 624432 581330 624484 581336
rect 623418 568844 623474 568853
rect 623418 568779 623474 568788
rect 623432 568406 623460 568779
rect 623420 568400 623472 568406
rect 623420 568342 623472 568348
rect 623328 506248 623380 506254
rect 623328 506190 623380 506196
rect 623326 455420 623382 455429
rect 623326 455355 623382 455364
rect 623340 454710 623368 455355
rect 623328 454704 623380 454710
rect 623328 454646 623380 454652
rect 623234 434204 623290 434213
rect 623234 434139 623290 434148
rect 623142 398844 623198 398853
rect 623142 398779 623198 398788
rect 623052 285452 623104 285458
rect 623052 285394 623104 285400
rect 624444 279950 624472 581330
rect 625088 280562 625116 694482
rect 635472 667204 635524 667210
rect 635472 667146 635524 667152
rect 633264 652312 633316 652318
rect 633264 652254 633316 652260
rect 628848 648436 628900 648442
rect 628848 648378 628900 648384
rect 625536 647484 625588 647490
rect 625536 647426 625588 647432
rect 625548 615870 625576 647426
rect 627742 647316 627798 647325
rect 627742 647251 627798 647260
rect 625536 615864 625588 615870
rect 625536 615806 625588 615812
rect 625536 605936 625588 605942
rect 625536 605878 625588 605884
rect 625076 280556 625128 280562
rect 625076 280498 625128 280504
rect 624432 279944 624484 279950
rect 624432 279886 624484 279892
rect 625548 279814 625576 605878
rect 625628 437160 625680 437166
rect 625628 437102 625680 437108
rect 625640 425334 625668 437102
rect 625628 425328 625680 425334
rect 625628 425270 625680 425276
rect 625536 279808 625588 279814
rect 625536 279750 625588 279756
rect 622960 278720 623012 278726
rect 622960 278662 623012 278668
rect 622868 262128 622920 262134
rect 622868 262070 622920 262076
rect 621856 262060 621908 262066
rect 621856 262002 621908 262008
rect 620016 260292 620068 260298
rect 620016 260234 620068 260240
rect 618636 260088 618688 260094
rect 618636 260030 618688 260036
rect 611736 260020 611788 260026
rect 611736 259962 611788 259968
rect 617256 260020 617308 260026
rect 617256 259962 617308 259968
rect 613024 259952 613076 259958
rect 613024 259894 613076 259900
rect 610892 259566 610960 259570
rect 613036 259566 613064 259894
rect 616336 259884 616388 259890
rect 616336 259826 616388 259832
rect 616348 259736 616376 259826
rect 617268 259736 617296 259962
rect 615598 259716 615654 259725
rect 616348 259708 616417 259736
rect 617268 259708 617339 259736
rect 615598 259651 615654 259660
rect 615612 259570 615640 259651
rect 610828 259564 610960 259566
rect 610828 259538 610908 259564
rect 610828 259470 610856 259538
rect 610908 259506 610960 259512
rect 612993 259538 613064 259566
rect 615600 259564 615652 259570
rect 612993 259470 613021 259538
rect 615600 259506 615652 259512
rect 616389 259470 616417 259708
rect 617311 259470 617339 259708
rect 618648 259566 618676 260030
rect 619256 259748 619308 259754
rect 619256 259690 619308 259696
rect 618648 259538 618710 259566
rect 618682 259470 618710 259538
rect 619268 259470 619296 259690
rect 620028 259566 620056 260234
rect 625260 260156 625312 260162
rect 625260 260098 625312 260104
rect 620660 259952 620712 259958
rect 620660 259894 620712 259900
rect 620198 259716 620254 259725
rect 620198 259651 620254 259660
rect 619997 259538 620056 259566
rect 619997 259470 620025 259538
rect 620212 259470 620240 259651
rect 620672 259470 620700 259894
rect 621856 259816 621908 259822
rect 621908 259764 621917 259804
rect 621856 259758 621917 259764
rect 621026 259716 621082 259725
rect 621026 259651 621082 259660
rect 621040 259470 621068 259651
rect 621889 259470 621917 259758
rect 623788 259748 623840 259754
rect 623084 259716 623140 259725
rect 623788 259690 623840 259696
rect 625120 259716 625176 259725
rect 623084 259651 623140 259660
rect 623098 259470 623126 259651
rect 623800 259470 623828 259690
rect 625120 259651 625176 259660
rect 625134 259566 625162 259651
rect 625272 259566 625300 260098
rect 627756 259618 627784 647251
rect 628860 635182 628888 648378
rect 631056 646872 631108 646878
rect 631056 646814 631108 646820
rect 628848 635176 628900 635182
rect 628848 635118 628900 635124
rect 629768 568468 629820 568474
rect 629768 568410 629820 568416
rect 629780 566706 629808 568410
rect 629768 566700 629820 566706
rect 629768 566642 629820 566648
rect 631068 530870 631096 646814
rect 631056 530864 631108 530870
rect 631056 530806 631108 530812
rect 627836 446340 627888 446346
rect 627836 446282 627888 446288
rect 627848 437166 627876 446282
rect 627836 437160 627888 437166
rect 627836 437102 627888 437108
rect 633276 280086 633304 652254
rect 635484 648442 635512 667146
rect 637232 666598 637260 728987
rect 637508 728682 637536 729366
rect 649308 729342 649916 729373
rect 650053 729486 650321 729514
rect 637678 729324 637734 729333
rect 637678 729259 637734 729268
rect 637692 728818 637720 729259
rect 637680 728812 637732 728818
rect 637680 728754 637732 728760
rect 637496 728676 637548 728682
rect 637496 728618 637548 728624
rect 649308 725492 649339 729342
rect 650053 729310 650081 729486
rect 650204 729430 650232 729486
rect 650434 729430 650462 729514
rect 650192 729424 650244 729430
rect 650192 729366 650244 729372
rect 650422 729424 650474 729430
rect 650422 729366 650474 729372
rect 651768 729362 651796 729514
rect 652474 729430 652502 729514
rect 653671 729494 653723 729552
rect 653424 729466 653723 729494
rect 652462 729424 652514 729430
rect 652462 729366 652514 729372
rect 649560 729282 650081 729310
rect 651756 729356 651808 729362
rect 652474 729333 652502 729366
rect 651756 729298 651808 729304
rect 652460 729324 652516 729333
rect 649560 728682 649588 729282
rect 649548 728676 649600 728682
rect 649548 728618 649600 728624
rect 651768 728546 651796 729298
rect 652460 729259 652516 729268
rect 651756 728540 651808 728546
rect 651756 728482 651808 728488
rect 649292 725440 649298 725492
rect 649350 725440 649356 725492
rect 653424 721270 653452 729466
rect 653671 729465 653723 729466
rect 654532 729333 654560 729514
rect 654896 729430 654924 729514
rect 654884 729424 654936 729430
rect 654884 729366 654936 729372
rect 654518 729324 654574 729333
rect 654518 729259 654574 729268
rect 654896 728818 654924 729366
rect 655362 729333 655390 729514
rect 655448 729486 655603 729514
rect 656276 729486 656332 729514
rect 655348 729324 655404 729333
rect 655348 729259 655404 729268
rect 654884 728812 654936 728818
rect 654884 728754 654936 728760
rect 655448 728750 655476 729486
rect 656276 729362 656304 729486
rect 656264 729356 656316 729362
rect 656264 729298 656316 729304
rect 655436 728744 655488 728750
rect 655436 728686 655488 728692
rect 654884 728676 654936 728682
rect 654884 728618 654936 728624
rect 652676 721264 652728 721270
rect 652676 721206 652728 721212
rect 653412 721264 653464 721270
rect 653412 721206 653464 721212
rect 646512 702020 646564 702026
rect 646512 701962 646564 701968
rect 643200 675976 643252 675982
rect 643200 675918 643252 675924
rect 643212 667210 643240 675918
rect 643200 667204 643252 667210
rect 643200 667146 643252 667152
rect 637220 666592 637272 666598
rect 637220 666534 637272 666540
rect 637680 657820 637732 657826
rect 637680 657762 637732 657768
rect 635472 648436 635524 648442
rect 635472 648378 635524 648384
rect 635472 646940 635524 646946
rect 635472 646882 635524 646888
rect 635484 529782 635512 646882
rect 635564 581932 635616 581938
rect 635564 581874 635616 581880
rect 635576 568406 635604 581874
rect 635564 568400 635616 568406
rect 635564 568342 635616 568348
rect 635472 529776 635524 529782
rect 635472 529718 635524 529724
rect 635472 426688 635524 426694
rect 635472 426630 635524 426636
rect 635484 423226 635512 426630
rect 635472 423220 635524 423226
rect 635472 423162 635524 423168
rect 634912 281126 636294 281152
rect 634912 280890 634944 281126
rect 636264 280890 636294 281126
rect 634912 280868 636294 280890
rect 633264 280080 633316 280086
rect 633264 280022 633316 280028
rect 637692 279882 637720 657762
rect 639518 650580 639574 650589
rect 639518 650515 639574 650524
rect 638784 646804 638836 646810
rect 638784 646746 638836 646752
rect 637772 587236 637824 587242
rect 637772 587178 637824 587184
rect 637784 581938 637812 587178
rect 637772 581932 637824 581938
rect 637772 581874 637824 581880
rect 637680 279876 637732 279882
rect 637680 279818 637732 279824
rect 638796 260094 638824 646746
rect 638876 473880 638928 473886
rect 638876 473822 638928 473828
rect 638888 446346 638916 473822
rect 638876 446340 638928 446346
rect 638876 446282 638928 446288
rect 639532 280766 639560 650515
rect 645408 647416 645460 647422
rect 645408 647358 645460 647364
rect 642096 647280 642148 647286
rect 642096 647222 642148 647228
rect 640992 647144 641044 647150
rect 640992 647086 641044 647092
rect 639888 601448 639940 601454
rect 639888 601390 639940 601396
rect 639900 587242 639928 601390
rect 639888 587236 639940 587242
rect 639888 587178 639940 587184
rect 639520 280760 639572 280766
rect 639520 280702 639572 280708
rect 640256 261992 640308 261998
rect 640256 261934 640308 261940
rect 638876 260904 638928 260910
rect 638876 260846 638928 260852
rect 638784 260088 638836 260094
rect 638784 260030 638836 260036
rect 638888 259822 638916 260846
rect 638876 259816 638928 259822
rect 638876 259758 638928 259764
rect 632526 259716 632582 259725
rect 632526 259651 632582 259660
rect 632540 259618 632568 259651
rect 625134 259538 625300 259566
rect 625674 259612 625726 259618
rect 625674 259554 625726 259560
rect 627744 259612 627796 259618
rect 627744 259554 627796 259560
rect 632528 259612 632580 259618
rect 640268 259589 640296 261934
rect 641004 259890 641032 647086
rect 641912 632456 641964 632462
rect 641912 632398 641964 632404
rect 641924 630762 641952 632398
rect 641912 630756 641964 630762
rect 641912 630698 641964 630704
rect 641084 547456 641136 547462
rect 641084 547398 641136 547404
rect 641096 541954 641124 547398
rect 641084 541948 641136 541954
rect 641084 541890 641136 541896
rect 641084 483264 641136 483270
rect 641084 483206 641136 483212
rect 641096 473886 641124 483206
rect 641084 473880 641136 473886
rect 641084 473822 641136 473828
rect 641084 436888 641136 436894
rect 641084 436830 641136 436836
rect 641096 426694 641124 436830
rect 641084 426688 641136 426694
rect 641084 426630 641136 426636
rect 642108 259958 642136 647222
rect 643200 617020 643252 617026
rect 643200 616962 643252 616968
rect 642298 280916 643130 280936
rect 642298 280712 642326 280916
rect 643110 280712 643130 280916
rect 642298 280692 643130 280712
rect 643212 280154 643240 616962
rect 643292 605392 643344 605398
rect 643292 605334 643344 605340
rect 643304 601454 643332 605334
rect 643292 601448 643344 601454
rect 643292 601390 643344 601396
rect 644304 541948 644356 541954
rect 644304 541890 644356 541896
rect 644316 538758 644344 541890
rect 644304 538752 644356 538758
rect 644304 538694 644356 538700
rect 645420 494490 645448 647358
rect 645500 626336 645552 626342
rect 645500 626278 645552 626284
rect 645512 605398 645540 626278
rect 645500 605392 645552 605398
rect 645500 605334 645552 605340
rect 645500 566700 645552 566706
rect 645500 566642 645552 566648
rect 645512 561946 645540 566642
rect 645500 561940 645552 561946
rect 645500 561882 645552 561888
rect 645408 494484 645460 494490
rect 645408 494426 645460 494432
rect 645408 491628 645460 491634
rect 645408 491570 645460 491576
rect 645420 483270 645448 491570
rect 645408 483264 645460 483270
rect 645408 483206 645460 483212
rect 644488 458512 644540 458518
rect 644488 458454 644540 458460
rect 644500 454710 644528 458454
rect 644488 454704 644540 454710
rect 644488 454646 644540 454652
rect 645408 444164 645460 444170
rect 645408 444106 645460 444112
rect 645420 436894 645448 444106
rect 645408 436888 645460 436894
rect 645408 436830 645460 436836
rect 643200 280148 643252 280154
rect 643200 280090 643252 280096
rect 646524 280018 646552 701962
rect 650928 681008 650980 681014
rect 650928 680950 650980 680956
rect 650940 675982 650968 680950
rect 650928 675976 650980 675982
rect 650928 675918 650980 675924
rect 652688 651706 652716 721206
rect 654240 698688 654292 698694
rect 654240 698630 654292 698636
rect 654252 681014 654280 698630
rect 654896 696518 654924 728618
rect 656276 728478 656304 729298
rect 656264 728472 656316 728478
rect 656264 728414 656316 728420
rect 658260 728246 658288 729521
rect 659183 729430 659211 729514
rect 659171 729424 659223 729430
rect 659171 729366 659223 729372
rect 659183 729333 659211 729366
rect 662579 729362 662607 729514
rect 664740 729430 664768 729514
rect 664728 729424 664780 729430
rect 664728 729366 664780 729372
rect 662567 729356 662619 729362
rect 659169 729324 659225 729333
rect 659169 729259 659225 729268
rect 662565 729324 662567 729333
rect 662619 729324 662621 729333
rect 662565 729259 662621 729268
rect 662579 729233 662607 729259
rect 664740 728614 664768 729366
rect 664818 729324 664874 729333
rect 664818 729259 664874 729268
rect 664728 728608 664780 728614
rect 664728 728550 664780 728556
rect 658242 728194 658248 728246
rect 658300 728194 658306 728246
rect 664832 696994 664860 729259
rect 675952 728608 676004 728614
rect 675952 728550 676004 728556
rect 675860 728472 675912 728478
rect 675860 728414 675912 728420
rect 673117 728192 673124 728244
rect 673176 728192 673182 728244
rect 664820 696988 664872 696994
rect 664820 696930 664872 696936
rect 667488 696988 667540 696994
rect 667488 696930 667540 696936
rect 654884 696512 654936 696518
rect 654884 696454 654936 696460
rect 667500 687678 667528 696930
rect 667488 687672 667540 687678
rect 667488 687614 667540 687620
rect 654240 681008 654292 681014
rect 654240 680950 654292 680956
rect 671352 661968 671404 661974
rect 671352 661910 671404 661916
rect 671364 661158 671392 661910
rect 671352 661152 671404 661158
rect 671352 661094 671404 661100
rect 652676 651700 652728 651706
rect 652676 651642 652728 651648
rect 668592 651700 668644 651706
rect 668592 651642 668644 651648
rect 666750 647452 666806 647461
rect 666750 647387 666806 647396
rect 666764 645994 666792 647387
rect 666752 645988 666804 645994
rect 666752 645930 666804 645936
rect 668604 637902 668632 651642
rect 671076 647892 671128 647898
rect 671076 647834 671128 647840
rect 671088 646198 671116 647834
rect 671904 647076 671956 647082
rect 671904 647018 671956 647024
rect 671076 646192 671128 646198
rect 671076 646134 671128 646140
rect 661968 637896 662020 637902
rect 661968 637838 662020 637844
rect 668592 637896 668644 637902
rect 668592 637838 668644 637844
rect 652032 630756 652084 630762
rect 652032 630698 652084 630704
rect 652044 615666 652072 630698
rect 661980 626342 662008 637838
rect 661968 626336 662020 626342
rect 661968 626278 662020 626284
rect 652032 615660 652084 615666
rect 652032 615602 652084 615608
rect 654240 615660 654292 615666
rect 654240 615602 654292 615608
rect 654252 602066 654280 615602
rect 669694 606244 669750 606253
rect 669694 606179 669750 606188
rect 669708 605942 669736 606179
rect 669696 605936 669748 605942
rect 669696 605878 669748 605884
rect 654240 602060 654292 602066
rect 654240 602002 654292 602008
rect 659760 602060 659812 602066
rect 659760 602002 659812 602008
rect 659772 587718 659800 602002
rect 659760 587712 659812 587718
rect 659760 587654 659812 587660
rect 667488 587712 667540 587718
rect 667488 587654 667540 587660
rect 667500 570650 667528 587654
rect 667488 570644 667540 570650
rect 667488 570586 667540 570592
rect 670798 565444 670854 565453
rect 670798 565379 670854 565388
rect 649824 561940 649876 561946
rect 649824 561882 649876 561888
rect 649836 545762 649864 561882
rect 670812 558954 670840 565379
rect 664176 558948 664228 558954
rect 664176 558890 664228 558896
rect 670800 558948 670852 558954
rect 670800 558890 670852 558896
rect 649824 545756 649876 545762
rect 649824 545698 649876 545704
rect 651296 545756 651348 545762
rect 651296 545698 651348 545704
rect 651308 543178 651336 545698
rect 651296 543172 651348 543178
rect 651296 543114 651348 543120
rect 661968 543172 662020 543178
rect 661968 543114 662020 543120
rect 648720 538752 648772 538758
rect 648720 538694 648772 538700
rect 648732 521418 648760 538694
rect 659760 525152 659812 525158
rect 659760 525094 659812 525100
rect 648720 521412 648772 521418
rect 648720 521354 648772 521360
rect 658656 521412 658708 521418
rect 658656 521354 658708 521360
rect 650928 512640 650980 512646
rect 650928 512582 650980 512588
rect 650940 491634 650968 512582
rect 658668 509314 658696 521354
rect 659772 512646 659800 525094
rect 659760 512640 659812 512646
rect 659760 512582 659812 512588
rect 658656 509308 658708 509314
rect 658656 509250 658708 509256
rect 661980 497142 662008 543114
rect 664188 525158 664216 558890
rect 671916 539846 671944 647018
rect 671904 539840 671956 539846
rect 671904 539782 671956 539788
rect 664176 525152 664228 525158
rect 664176 525094 664228 525100
rect 668592 517060 668644 517066
rect 668592 517002 668644 517008
rect 668604 502378 668632 517002
rect 666384 502372 666436 502378
rect 666384 502314 666436 502320
rect 668592 502372 668644 502378
rect 668592 502314 668644 502320
rect 666396 499182 666424 502314
rect 662060 499176 662112 499182
rect 662060 499118 662112 499124
rect 666384 499176 666436 499182
rect 666384 499118 666436 499124
rect 661968 497136 662020 497142
rect 661968 497078 662020 497084
rect 662072 493306 662100 499118
rect 669696 497136 669748 497142
rect 669696 497078 669748 497084
rect 669708 493334 669736 497078
rect 673136 494143 673164 728192
rect 675872 701142 675900 728414
rect 675964 702570 675992 728550
rect 676056 702988 676437 703016
rect 675952 702564 676004 702570
rect 675952 702506 676004 702512
rect 676056 702026 676084 702988
rect 676332 702579 676437 702607
rect 676228 702564 676280 702570
rect 676228 702506 676280 702512
rect 676240 702462 676268 702506
rect 676332 702462 676360 702579
rect 676240 702434 676437 702462
rect 676044 702020 676096 702026
rect 676044 701962 676096 701968
rect 675860 701136 675912 701142
rect 675860 701078 675912 701084
rect 675676 697532 675728 697538
rect 675676 697474 675728 697480
rect 675584 696580 675636 696586
rect 675584 696522 675636 696528
rect 675596 694234 675624 696522
rect 675688 694546 675716 697474
rect 675872 696586 675900 701078
rect 676240 700426 676268 702434
rect 676320 701137 676372 701142
rect 676320 701136 676437 701137
rect 676372 701109 676437 701136
rect 676320 701078 676372 701084
rect 676240 700398 676437 700426
rect 676240 698650 676268 700398
rect 676332 699189 676437 699217
rect 676332 698762 676360 699189
rect 676320 698756 676372 698762
rect 676320 698698 676372 698704
rect 676172 698622 676268 698650
rect 676172 698370 676200 698622
rect 676172 698342 676437 698370
rect 675952 698000 676004 698006
rect 675952 697942 676004 697948
rect 675860 696580 675912 696586
rect 675860 696522 675912 696528
rect 675768 696104 675820 696110
rect 675768 696046 675820 696052
rect 675676 694540 675728 694546
rect 675676 694482 675728 694488
rect 675596 694206 675716 694234
rect 675688 687134 675716 694206
rect 675676 687128 675728 687134
rect 675676 687070 675728 687076
rect 675780 687066 675808 696046
rect 675860 695424 675912 695430
rect 675860 695366 675912 695372
rect 675872 694070 675900 695366
rect 675860 694064 675912 694070
rect 675860 694006 675912 694012
rect 675964 693950 675992 697942
rect 676172 697538 676200 698342
rect 676326 698002 676378 698008
rect 676378 697950 676452 698002
rect 676326 697944 676378 697950
rect 676044 697532 676437 697538
rect 676096 697510 676437 697532
rect 676044 697474 676096 697480
rect 676056 697297 676437 697325
rect 676056 696518 676084 697297
rect 676332 696586 676437 696596
rect 676320 696580 676437 696586
rect 676372 696568 676437 696580
rect 676320 696522 676372 696528
rect 676044 696512 676096 696518
rect 676044 696454 676096 696460
rect 676056 696110 676084 696454
rect 676044 696104 676096 696110
rect 676044 696046 676096 696052
rect 676056 695982 676437 696010
rect 676056 695430 676084 695982
rect 676044 695424 676096 695430
rect 676044 695366 676096 695372
rect 676056 694602 676437 694630
rect 676056 694274 676084 694602
rect 676136 694540 676188 694546
rect 676134 694508 676136 694517
rect 676188 694508 676190 694517
rect 676134 694443 676190 694452
rect 676044 694268 676096 694274
rect 676044 694210 676096 694216
rect 676148 694234 676176 694443
rect 676148 694206 676268 694234
rect 676136 694064 676188 694070
rect 676136 694006 676188 694012
rect 675872 693922 675992 693950
rect 675872 690330 675900 693922
rect 675860 690324 675912 690330
rect 675860 690266 675912 690272
rect 675872 689854 675900 690266
rect 675860 689848 675912 689854
rect 675860 689790 675912 689796
rect 676044 688148 676096 688154
rect 676044 688090 676096 688096
rect 676148 688102 676176 694006
rect 676240 691220 676268 694206
rect 676332 693689 676437 693717
rect 676332 693186 676360 693689
rect 676320 693180 676372 693186
rect 676320 693122 676372 693128
rect 676228 691214 676280 691220
rect 676228 691156 676280 691162
rect 676240 688238 676268 691156
rect 676320 690324 676372 690330
rect 676372 690293 676437 690321
rect 676320 690266 676372 690272
rect 676240 688210 676360 688238
rect 676332 688170 676360 688210
rect 676332 688154 676437 688170
rect 676320 688148 676437 688154
rect 675950 687980 676006 687989
rect 675950 687915 676006 687924
rect 675964 687678 675992 687915
rect 675952 687672 676004 687678
rect 675952 687614 676004 687620
rect 675768 687060 675820 687066
rect 675768 687002 675820 687008
rect 675676 664008 675728 664014
rect 675676 663950 675728 663956
rect 675688 662314 675716 663950
rect 675860 663668 675912 663674
rect 675860 663610 675912 663616
rect 675768 662988 675820 662994
rect 675768 662930 675820 662936
rect 675676 662308 675728 662314
rect 675676 662250 675728 662256
rect 675780 660342 675808 662930
rect 675768 660336 675820 660342
rect 675768 660278 675820 660284
rect 675676 658160 675728 658166
rect 675676 658102 675728 658108
rect 675584 657412 675636 657418
rect 675584 657354 675636 657360
rect 675596 656738 675624 657354
rect 675584 656732 675636 656738
rect 675584 656674 675636 656680
rect 675492 654284 675544 654290
rect 675492 654226 675544 654232
rect 675504 648986 675532 654226
rect 675596 653853 675624 656674
rect 675688 655650 675716 658102
rect 675780 656058 675808 660278
rect 675872 656262 675900 663610
rect 675860 656256 675912 656262
rect 675860 656198 675912 656204
rect 675768 656052 675820 656058
rect 675768 655994 675820 656000
rect 675676 655644 675728 655650
rect 675676 655586 675728 655592
rect 675582 653844 675638 653853
rect 675582 653779 675638 653788
rect 675584 651632 675636 651638
rect 675584 651574 675636 651580
rect 675492 648980 675544 648986
rect 675492 648922 675544 648928
rect 675214 646908 675270 646917
rect 675214 646843 675270 646852
rect 673376 581388 673428 581394
rect 673376 581330 673428 581336
rect 673388 580578 673416 581330
rect 673376 580572 673428 580578
rect 673376 580514 673428 580520
rect 674112 572344 674164 572350
rect 674112 572286 674164 572292
rect 673376 495164 673428 495170
rect 673376 495106 673428 495112
rect 673388 494490 673416 495106
rect 673376 494484 673428 494490
rect 673376 494426 673428 494432
rect 673136 494115 673359 494143
rect 661980 493278 662100 493306
rect 669696 493328 669748 493334
rect 660864 492240 660916 492246
rect 660864 492182 660916 492188
rect 650928 491628 650980 491634
rect 650928 491570 650980 491576
rect 659760 483400 659812 483406
rect 659760 483342 659812 483348
rect 657552 475580 657604 475586
rect 657552 475522 657604 475528
rect 656448 462932 656500 462938
rect 656448 462874 656500 462880
rect 656460 458518 656488 462874
rect 656448 458512 656500 458518
rect 656448 458454 656500 458460
rect 657564 444170 657592 475522
rect 657552 444164 657604 444170
rect 657552 444106 657604 444112
rect 646512 280012 646564 280018
rect 646512 279954 646564 279960
rect 652584 260292 652636 260298
rect 652584 260234 652636 260240
rect 643384 260156 643436 260162
rect 643384 260098 643436 260104
rect 643016 260020 643068 260026
rect 643016 259962 643068 259968
rect 642096 259952 642148 259958
rect 642096 259894 642148 259900
rect 640992 259884 641044 259890
rect 640992 259826 641044 259832
rect 632528 259554 632580 259560
rect 640254 259580 640310 259589
rect 625134 259470 625162 259538
rect 625272 259470 625300 259538
rect 625686 259470 625714 259554
rect 640254 259515 640310 259524
rect 643028 259470 643056 259962
rect 643396 259686 643424 260098
rect 645592 260088 645644 260094
rect 645592 260030 645644 260036
rect 643384 259680 643436 259686
rect 643384 259622 643436 259628
rect 643396 259566 643424 259622
rect 643396 259538 643466 259566
rect 643438 259470 643466 259538
rect 645604 259470 645632 260030
rect 649916 259952 649968 259958
rect 649916 259894 649968 259900
rect 648996 259884 649048 259890
rect 648996 259826 649048 259832
rect 646462 259740 646514 259746
rect 649008 259702 649036 259826
rect 649928 259804 649956 259894
rect 651296 259884 651348 259890
rect 651296 259826 651348 259832
rect 646462 259682 646514 259688
rect 646474 259598 646502 259682
rect 648989 259674 649036 259702
rect 649911 259776 649956 259804
rect 649640 259680 649692 259686
rect 646462 259592 646514 259598
rect 646462 259534 646514 259540
rect 648989 259470 649017 259674
rect 649640 259623 649692 259628
rect 649638 259614 649694 259623
rect 649638 259549 649694 259558
rect 649911 259470 649939 259776
rect 651308 259566 651336 259826
rect 651856 259748 651908 259754
rect 651854 259716 651856 259725
rect 651908 259716 651910 259725
rect 651854 259651 651910 259660
rect 651282 259538 651336 259566
rect 651282 259470 651310 259538
rect 651868 259470 651896 259651
rect 652596 259470 652624 260234
rect 653228 260088 653280 260094
rect 653228 260030 653280 260036
rect 653240 259804 653268 260030
rect 657828 259884 657880 259890
rect 657828 259826 657880 259832
rect 653240 259776 653290 259804
rect 652798 259680 652850 259686
rect 652798 259622 652850 259628
rect 652810 259470 652838 259622
rect 653262 259470 653290 259776
rect 654477 259748 654529 259754
rect 654477 259690 654529 259696
rect 656400 259716 656456 259725
rect 653628 259680 653680 259686
rect 653628 259622 653680 259628
rect 653640 259470 653668 259622
rect 654489 259470 654517 259690
rect 655686 259680 655738 259686
rect 657840 259686 657868 259826
rect 659772 259754 659800 483342
rect 659760 259748 659812 259754
rect 660876 259725 660904 492182
rect 661980 475586 662008 493278
rect 669696 493270 669748 493276
rect 661968 475580 662020 475586
rect 661968 475522 662020 475528
rect 671904 475444 671956 475450
rect 671904 475386 671956 475392
rect 671916 462938 671944 475386
rect 671904 462932 671956 462938
rect 671904 462874 671956 462880
rect 673331 277960 673359 494115
rect 674124 280533 674152 572286
rect 674202 524372 674258 524381
rect 674202 524307 674258 524316
rect 674216 517066 674244 524307
rect 674204 517060 674256 517066
rect 674204 517002 674256 517008
rect 674110 280524 674166 280533
rect 674110 280459 674166 280468
rect 675228 279746 675256 646843
rect 675596 643954 675624 651574
rect 675688 647014 675716 655586
rect 675768 654216 675820 654222
rect 675768 654158 675820 654164
rect 675780 651434 675808 654158
rect 675872 651638 675900 656198
rect 675964 654290 675992 687614
rect 676056 664014 676084 688090
rect 676148 688074 676268 688102
rect 676372 688142 676437 688148
rect 676320 688090 676372 688096
rect 676134 687844 676190 687853
rect 676134 687779 676190 687788
rect 676148 666093 676176 687779
rect 676240 687751 676268 688074
rect 676332 688059 676360 688090
rect 676240 687723 676437 687751
rect 676332 687660 676360 687723
rect 676332 687632 676728 687660
rect 676320 687128 676372 687134
rect 676320 687070 676372 687076
rect 676228 687060 676280 687066
rect 676228 687002 676280 687008
rect 676134 666084 676190 666093
rect 676134 666019 676190 666028
rect 676044 664008 676096 664014
rect 676044 663950 676096 663956
rect 676044 663872 676096 663878
rect 676044 663814 676096 663820
rect 676056 658166 676084 663814
rect 676240 663674 676268 687002
rect 676332 678778 676360 687070
rect 676332 678750 676636 678778
rect 676228 663668 676280 663674
rect 676228 663610 676280 663616
rect 676608 663054 676636 678750
rect 676700 663878 676728 687632
rect 676688 663872 676740 663878
rect 676688 663814 676740 663820
rect 676596 663048 676648 663054
rect 676596 662990 676648 662996
rect 676136 662308 676188 662314
rect 676136 662250 676188 662256
rect 676148 661650 676176 662250
rect 676332 662188 676437 662216
rect 676332 661974 676360 662188
rect 676320 661968 676372 661974
rect 676320 661910 676372 661916
rect 676332 661779 676437 661807
rect 676332 661650 676360 661779
rect 676148 661622 676437 661650
rect 676148 659626 676176 661622
rect 676320 660337 676372 660342
rect 676320 660336 676437 660337
rect 676372 660309 676437 660336
rect 676320 660278 676372 660284
rect 676148 659598 676437 659626
rect 676044 658160 676096 658166
rect 676044 658102 676096 658108
rect 676148 657568 676176 659598
rect 676240 658389 676437 658417
rect 676240 657826 676268 658389
rect 676228 657820 676280 657826
rect 676228 657762 676280 657768
rect 676148 657540 676437 657568
rect 676240 657418 676268 657540
rect 676228 657412 676280 657418
rect 676228 657354 676280 657360
rect 676332 657162 676437 657190
rect 676332 656822 676360 657162
rect 676056 656794 676360 656822
rect 675952 654284 676004 654290
rect 675952 654226 676004 654232
rect 676056 654222 676084 656794
rect 676320 656732 676437 656738
rect 676372 656710 676437 656732
rect 676320 656674 676372 656680
rect 676332 656497 676437 656525
rect 676332 656262 676360 656497
rect 676320 656256 676372 656262
rect 676320 656198 676372 656204
rect 676136 656052 676188 656058
rect 676136 655994 676188 656000
rect 676148 655802 676176 655994
rect 676148 655774 676437 655802
rect 676044 654216 676096 654222
rect 676044 654158 676096 654164
rect 676148 654102 676176 655774
rect 676320 655644 676372 655650
rect 676320 655586 676372 655592
rect 676332 655210 676360 655586
rect 676332 655182 676437 655210
rect 675964 654074 676176 654102
rect 675860 651632 675912 651638
rect 675860 651574 675912 651580
rect 675768 651428 675820 651434
rect 675768 651370 675820 651376
rect 675964 649206 675992 654074
rect 676056 653938 676268 653966
rect 676056 651706 676084 653938
rect 676134 653844 676190 653853
rect 676240 653839 676268 653938
rect 676240 653811 676437 653839
rect 676134 653779 676190 653788
rect 676044 651700 676096 651706
rect 676044 651642 676096 651648
rect 676148 650420 676176 653779
rect 676240 652889 676437 652917
rect 676240 652454 676268 652889
rect 676228 652448 676280 652454
rect 676228 652390 676280 652396
rect 676228 651428 676280 651434
rect 676228 651370 676280 651376
rect 676136 650414 676188 650420
rect 676136 650356 676188 650362
rect 675780 649178 675992 649206
rect 675676 647008 675728 647014
rect 675676 646950 675728 646956
rect 675780 644838 675808 649178
rect 675860 649048 675912 649054
rect 675860 648990 675912 648996
rect 675872 647302 675900 648990
rect 675952 648980 676004 648986
rect 675952 648922 676004 648928
rect 675964 647710 675992 648922
rect 676148 647866 676176 650356
rect 676240 649521 676268 651370
rect 676240 649493 676437 649521
rect 676240 649122 676268 649493
rect 676228 649116 676280 649122
rect 676228 649058 676280 649064
rect 676148 647838 676268 647866
rect 675964 647682 676176 647710
rect 675872 647274 675992 647302
rect 675768 644832 675820 644838
rect 675768 644774 675820 644780
rect 675584 643948 675636 643954
rect 675584 643890 675636 643896
rect 675860 631776 675912 631782
rect 675860 631718 675912 631724
rect 675768 628784 675820 628790
rect 675768 628726 675820 628732
rect 675676 628716 675728 628722
rect 675676 628658 675728 628664
rect 675584 622392 675636 622398
rect 675584 622334 675636 622340
rect 675308 621372 675360 621378
rect 675308 621314 675360 621320
rect 675320 614306 675348 621314
rect 675596 616142 675624 622334
rect 675688 621038 675716 628658
rect 675676 621032 675728 621038
rect 675676 620974 675728 620980
rect 675780 616954 675808 628726
rect 675872 621378 675900 631718
rect 675860 621372 675912 621378
rect 675860 621314 675912 621320
rect 675860 621236 675912 621242
rect 675860 621178 675912 621184
rect 675872 619542 675900 621178
rect 675860 619536 675912 619542
rect 675860 619478 675912 619484
rect 675688 616926 675808 616954
rect 675584 616136 675636 616142
rect 675584 616078 675636 616084
rect 675492 615932 675544 615938
rect 675492 615874 675544 615880
rect 675400 615796 675452 615802
rect 675400 615738 675452 615744
rect 675308 614300 675360 614306
rect 675308 614242 675360 614248
rect 675412 614118 675440 615738
rect 675504 615734 675532 615874
rect 675492 615728 675544 615734
rect 675492 615670 675544 615676
rect 675320 614090 675440 614118
rect 675320 613053 675348 614090
rect 675400 613552 675452 613558
rect 675400 613494 675452 613500
rect 675306 613044 675362 613053
rect 675306 612979 675362 612988
rect 675320 609614 675348 612979
rect 675308 609608 675360 609614
rect 675308 609550 675360 609556
rect 675320 606622 675348 609550
rect 675308 606616 675360 606622
rect 675308 606558 675360 606564
rect 675320 605262 675348 606558
rect 675412 606214 675440 613494
rect 675504 611382 675532 615670
rect 675688 613558 675716 616926
rect 675768 615864 675820 615870
rect 675768 615806 675820 615812
rect 675676 613552 675728 613558
rect 675676 613494 675728 613500
rect 675584 613144 675636 613150
rect 675584 613086 675636 613092
rect 675492 611376 675544 611382
rect 675492 611318 675544 611324
rect 675492 609064 675544 609070
rect 675492 609006 675544 609012
rect 675400 606208 675452 606214
rect 675400 606150 675452 606156
rect 675308 605256 675360 605262
rect 675308 605198 675360 605204
rect 675504 605194 675532 609006
rect 675596 606389 675624 613086
rect 675676 612260 675728 612266
rect 675676 612202 675728 612208
rect 675582 606380 675638 606389
rect 675582 606315 675638 606324
rect 675596 605874 675624 606315
rect 675584 605868 675636 605874
rect 675584 605810 675636 605816
rect 675688 605330 675716 612202
rect 675780 609002 675808 615806
rect 675872 614986 675900 619478
rect 675860 614980 675912 614986
rect 675860 614922 675912 614928
rect 675872 611994 675900 614922
rect 675860 611988 675912 611994
rect 675860 611930 675912 611936
rect 675860 609132 675912 609138
rect 675860 609074 675912 609080
rect 675768 608996 675820 609002
rect 675768 608938 675820 608944
rect 675768 608180 675820 608186
rect 675768 608122 675820 608128
rect 675676 605324 675728 605330
rect 675676 605266 675728 605272
rect 675492 605188 675544 605194
rect 675492 605130 675544 605136
rect 675780 605126 675808 608122
rect 675872 605398 675900 609074
rect 675964 609070 675992 647274
rect 676148 647189 676176 647682
rect 676240 647370 676268 647838
rect 676240 647342 676437 647370
rect 676134 647180 676190 647189
rect 676134 647115 676190 647124
rect 676042 647044 676098 647053
rect 676042 646979 676098 646988
rect 675952 609064 676004 609070
rect 675952 609006 676004 609012
rect 676056 606638 676084 646979
rect 676148 646622 676176 647115
rect 676240 646810 676268 647342
rect 676320 647008 676372 647014
rect 676320 646951 676372 646956
rect 676320 646950 676437 646951
rect 676332 646923 676437 646950
rect 676332 646860 676360 646923
rect 676332 646832 676728 646860
rect 676228 646804 676280 646810
rect 676228 646746 676280 646752
rect 676148 646594 676360 646622
rect 676228 646532 676280 646538
rect 676228 646474 676280 646480
rect 676136 646192 676188 646198
rect 676136 646134 676188 646140
rect 675964 606610 676084 606638
rect 676148 606638 676176 646134
rect 676240 628722 676268 646474
rect 676332 631782 676360 646594
rect 676596 645988 676648 645994
rect 676596 645930 676648 645936
rect 676504 644832 676556 644838
rect 676504 644774 676556 644780
rect 676412 643948 676464 643954
rect 676412 643890 676464 643896
rect 676320 631776 676372 631782
rect 676320 631718 676372 631724
rect 676320 631640 676372 631646
rect 676320 631582 676372 631588
rect 676332 628790 676360 631582
rect 676424 631390 676452 643890
rect 676516 631510 676544 644774
rect 676504 631504 676556 631510
rect 676504 631446 676556 631452
rect 676424 631362 676544 631390
rect 676320 628784 676372 628790
rect 676320 628726 676372 628732
rect 676228 628716 676280 628722
rect 676228 628658 676280 628664
rect 676228 628580 676280 628586
rect 676228 628522 676280 628528
rect 676240 621242 676268 628522
rect 676516 622398 676544 631362
rect 676504 622392 676556 622398
rect 676504 622334 676556 622340
rect 676608 622176 676636 645930
rect 676700 631646 676728 646832
rect 676688 631640 676740 631646
rect 676688 631582 676740 631588
rect 676688 631504 676740 631510
rect 676688 631446 676740 631452
rect 676700 628586 676728 631446
rect 676688 628580 676740 628586
rect 676688 628522 676740 628528
rect 676332 622148 676636 622176
rect 676332 621416 676360 622148
rect 676332 621388 676437 621416
rect 676228 621236 676280 621242
rect 676228 621178 676280 621184
rect 676320 621032 676372 621038
rect 676372 620980 676437 621007
rect 676320 620979 676437 620980
rect 676320 620974 676372 620979
rect 676332 620850 676360 620974
rect 676240 620822 676437 620850
rect 676240 618742 676268 620822
rect 676320 619537 676372 619542
rect 676320 619536 676437 619537
rect 676372 619509 676437 619536
rect 676320 619478 676372 619484
rect 676332 618798 676437 618826
rect 676332 618742 676360 618798
rect 676240 618714 676360 618742
rect 676240 616768 676268 618714
rect 676332 617589 676437 617617
rect 676332 617026 676360 617589
rect 676320 617020 676372 617026
rect 676320 616962 676372 616968
rect 676240 616740 676437 616768
rect 676240 616482 676268 616740
rect 676228 616476 676280 616482
rect 676228 616418 676280 616424
rect 676240 616362 676437 616390
rect 676240 615870 676268 616362
rect 676320 616272 676372 616278
rect 676320 616214 676372 616220
rect 676332 615938 676360 616214
rect 676332 615910 676437 615938
rect 676332 615870 676360 615910
rect 676228 615864 676280 615870
rect 676228 615806 676280 615812
rect 676320 615864 676372 615870
rect 676320 615806 676372 615812
rect 676228 615728 676280 615734
rect 676280 615697 676437 615725
rect 676228 615670 676280 615676
rect 676240 614986 676437 615002
rect 676228 614980 676437 614986
rect 676280 614974 676437 614980
rect 676228 614922 676280 614928
rect 676240 614382 676437 614410
rect 676240 613558 676268 614382
rect 676320 614300 676372 614306
rect 676320 614242 676372 614248
rect 676228 613552 676280 613558
rect 676228 613494 676280 613500
rect 676332 613150 676360 614242
rect 676320 613144 676372 613150
rect 676320 613086 676372 613092
rect 676240 613002 676437 613030
rect 676240 612266 676268 613002
rect 676228 612260 676280 612266
rect 676228 612202 676280 612208
rect 676240 612089 676437 612117
rect 676240 611518 676268 612089
rect 676320 611988 676372 611994
rect 676320 611930 676372 611936
rect 676228 611512 676280 611518
rect 676228 611454 676280 611460
rect 676228 611376 676280 611382
rect 676228 611318 676280 611324
rect 676240 608186 676268 611318
rect 676332 609138 676360 611930
rect 676320 609132 676372 609138
rect 676320 609074 676372 609080
rect 676320 608996 676372 609002
rect 676320 608938 676372 608944
rect 676332 608721 676360 608938
rect 676332 608693 676437 608721
rect 676228 608180 676280 608186
rect 676228 608122 676280 608128
rect 676148 606610 676268 606638
rect 675860 605392 675912 605398
rect 675964 605380 675992 606610
rect 676240 605380 676268 606610
rect 676320 606616 676372 606622
rect 676372 606564 676437 606570
rect 676320 606558 676437 606564
rect 676332 606542 676437 606558
rect 676320 606208 676372 606214
rect 676320 606151 676372 606156
rect 676320 606150 676437 606151
rect 676332 606123 676437 606150
rect 676332 605992 676360 606123
rect 676332 605964 676728 605992
rect 676320 605868 676372 605874
rect 676320 605810 676372 605816
rect 675964 605352 676084 605380
rect 675860 605334 675912 605340
rect 675860 605256 675912 605262
rect 675860 605198 675912 605204
rect 675768 605120 675820 605126
rect 675768 605062 675820 605068
rect 675768 582068 675820 582074
rect 675768 582010 675820 582016
rect 675584 581456 675636 581462
rect 675584 581398 675636 581404
rect 675400 580096 675452 580102
rect 675400 580038 675452 580044
rect 675412 578266 675440 580038
rect 675596 578742 675624 581398
rect 675676 578872 675728 578878
rect 675676 578814 675728 578820
rect 675584 578736 675636 578742
rect 675584 578678 675636 578684
rect 675400 578260 675452 578266
rect 675400 578202 675452 578208
rect 675492 578192 675544 578198
rect 675492 578134 675544 578140
rect 675504 575614 675532 578134
rect 675492 575608 675544 575614
rect 675492 575550 675544 575556
rect 675308 574996 675360 575002
rect 675308 574938 675360 574944
rect 675320 574186 675348 574938
rect 675308 574180 675360 574186
rect 675308 574122 675360 574128
rect 675504 574134 675532 575550
rect 675596 575002 675624 578678
rect 675688 575818 675716 578814
rect 675676 575812 675728 575818
rect 675676 575754 675728 575760
rect 675596 574996 675728 575002
rect 675596 574974 675676 574996
rect 675676 574938 675728 574944
rect 675780 574934 675808 582010
rect 675872 580102 675900 605198
rect 675952 605188 676004 605194
rect 675952 605130 676004 605136
rect 675860 580096 675912 580102
rect 675860 580038 675912 580044
rect 675964 578198 675992 605130
rect 675952 578192 676004 578198
rect 675952 578134 676004 578140
rect 676056 578078 676084 605352
rect 676148 605352 676268 605380
rect 676148 578130 676176 605352
rect 676228 605120 676280 605126
rect 676228 605062 676280 605068
rect 676240 578878 676268 605062
rect 676332 582278 676360 605810
rect 676504 605392 676556 605398
rect 676504 605334 676556 605340
rect 676320 582272 676372 582278
rect 676320 582214 676372 582220
rect 676516 581462 676544 605334
rect 676596 605324 676648 605330
rect 676596 605266 676648 605272
rect 676608 581501 676636 605266
rect 676700 581637 676728 605964
rect 676686 581628 676742 581637
rect 676686 581563 676742 581572
rect 676594 581492 676650 581501
rect 676504 581456 676556 581462
rect 676594 581427 676650 581436
rect 676504 581398 676556 581404
rect 676320 580640 676372 580646
rect 676372 580588 676437 580616
rect 676320 580582 676372 580588
rect 676320 580232 676372 580238
rect 676372 580180 676437 580207
rect 676320 580179 676437 580180
rect 676320 580174 676372 580179
rect 676320 580096 676372 580102
rect 676372 580044 676437 580062
rect 676320 580038 676437 580044
rect 676332 580034 676437 580038
rect 676228 578872 676280 578878
rect 676228 578814 676280 578820
rect 676228 578737 676280 578742
rect 676228 578736 676437 578737
rect 676280 578709 676437 578736
rect 676228 578678 676280 578684
rect 676228 578260 676280 578266
rect 676228 578202 676280 578208
rect 675872 578050 676084 578078
rect 676136 578124 676188 578130
rect 676136 578066 676188 578072
rect 675872 575902 675900 578050
rect 676240 578026 676268 578202
rect 676240 577998 676437 578026
rect 676136 577988 676188 577994
rect 676136 577930 676188 577936
rect 676148 576090 676176 577930
rect 676136 576084 676188 576090
rect 676136 576026 676188 576032
rect 676240 575968 676268 577998
rect 676332 576789 676437 576817
rect 676332 576158 676360 576789
rect 676320 576152 676372 576158
rect 676320 576094 676372 576100
rect 676136 575948 676188 575954
rect 675872 575874 676084 575902
rect 676136 575890 676188 575896
rect 676240 575940 676437 575968
rect 675952 575812 676004 575818
rect 675952 575754 676004 575760
rect 675860 575744 675912 575750
rect 675860 575686 675912 575692
rect 675872 575138 675900 575686
rect 675860 575132 675912 575138
rect 675860 575074 675912 575080
rect 675768 574928 675820 574934
rect 675768 574870 675820 574876
rect 675676 574860 675728 574866
rect 675676 574802 675728 574808
rect 675766 574828 675822 574837
rect 675320 563850 675348 574122
rect 675504 574106 675624 574134
rect 675490 574012 675546 574021
rect 675490 573947 675546 573956
rect 675504 573642 675532 573947
rect 675492 573636 675544 573642
rect 675492 573578 675544 573584
rect 675398 572244 675454 572253
rect 675398 572179 675454 572188
rect 675412 568814 675440 572179
rect 675400 568808 675452 568814
rect 675400 568750 675452 568756
rect 675400 567856 675452 567862
rect 675400 567798 675452 567804
rect 675412 565074 675440 567798
rect 675504 565414 675532 573578
rect 675596 571194 675624 574106
rect 675584 571188 675636 571194
rect 675584 571130 675636 571136
rect 675584 571052 675636 571058
rect 675584 570994 675636 571000
rect 675492 565408 675544 565414
rect 675492 565350 675544 565356
rect 675400 565068 675452 565074
rect 675400 565010 675452 565016
rect 675308 563844 675360 563850
rect 675308 563786 675360 563792
rect 675596 563442 675624 570994
rect 675688 567862 675716 574802
rect 675766 574763 675822 574772
rect 675676 567856 675728 567862
rect 675676 567798 675728 567804
rect 675676 567720 675728 567726
rect 675676 567662 675728 567668
rect 675688 565754 675716 567662
rect 675676 565748 675728 565754
rect 675676 565690 675728 565696
rect 675584 563436 675636 563442
rect 675584 563378 675636 563384
rect 675688 559546 675716 565690
rect 675780 564598 675808 574763
rect 675872 572253 675900 575074
rect 675964 574798 675992 575754
rect 676056 575002 676084 575874
rect 676148 575002 676176 575890
rect 676240 575750 676268 575940
rect 676228 575744 676280 575750
rect 676228 575686 676280 575692
rect 676228 575608 676280 575614
rect 676280 575562 676437 575590
rect 676228 575550 676280 575556
rect 676228 575472 676280 575478
rect 676228 575414 676280 575420
rect 676044 574996 676096 575002
rect 676044 574938 676096 574944
rect 676136 574996 676188 575002
rect 676136 574938 676188 574944
rect 676044 574860 676096 574866
rect 676044 574802 676096 574808
rect 676136 574860 676188 574866
rect 676136 574802 676188 574808
rect 675952 574792 676004 574798
rect 675952 574734 676004 574740
rect 675858 572244 675914 572253
rect 675858 572179 675914 572188
rect 675860 571528 675912 571534
rect 675860 571470 675912 571476
rect 675872 566790 675900 571470
rect 675964 571058 675992 574734
rect 675952 571052 676004 571058
rect 675952 570994 676004 571000
rect 675952 568808 676004 568814
rect 675952 568750 676004 568756
rect 675964 567726 675992 568750
rect 675952 567720 676004 567726
rect 675952 567662 676004 567668
rect 675872 566762 675992 566790
rect 675768 564592 675820 564598
rect 675768 564534 675820 564540
rect 675688 559518 675900 559546
rect 675872 547402 675900 559518
rect 675596 547374 675900 547402
rect 675596 544090 675624 547374
rect 675504 544062 675624 544090
rect 675400 540588 675452 540594
rect 675400 540530 675452 540536
rect 675412 536362 675440 540530
rect 675504 539234 675532 544062
rect 675860 543716 675912 543722
rect 675860 543658 675912 543664
rect 675768 543648 675820 543654
rect 675768 543590 675820 543596
rect 675584 540520 675636 540526
rect 675584 540462 675636 540468
rect 675492 539228 675544 539234
rect 675492 539170 675544 539176
rect 675596 537738 675624 540462
rect 675676 540452 675728 540458
rect 675676 540394 675728 540400
rect 675584 537732 675636 537738
rect 675584 537674 675636 537680
rect 675412 536334 675532 536362
rect 675400 535216 675452 535222
rect 675400 535158 675452 535164
rect 675412 533930 675440 535158
rect 675400 533924 675452 533930
rect 675400 533866 675452 533872
rect 675504 532638 675532 536334
rect 675596 533250 675624 537674
rect 675688 536854 675716 540394
rect 675676 536848 675728 536854
rect 675676 536790 675728 536796
rect 675676 536032 675728 536038
rect 675676 535974 675728 535980
rect 675688 534610 675716 535974
rect 675676 534604 675728 534610
rect 675676 534546 675728 534552
rect 675584 533244 675636 533250
rect 675584 533186 675636 533192
rect 675492 532632 675544 532638
rect 675492 532574 675544 532580
rect 675504 532518 675532 532574
rect 675504 532490 675624 532518
rect 675596 524682 675624 532490
rect 675688 530258 675716 534546
rect 675780 532541 675808 543590
rect 675872 535222 675900 543658
rect 675860 535216 675912 535222
rect 675860 535158 675912 535164
rect 675964 535068 675992 566762
rect 676056 535086 676084 574802
rect 676148 539710 676176 574802
rect 676240 572350 676268 575414
rect 676320 575132 676437 575138
rect 676372 575110 676437 575132
rect 676320 575074 676372 575080
rect 676332 574897 676437 574925
rect 676332 574798 676360 574897
rect 676320 574792 676372 574798
rect 676320 574734 676372 574740
rect 676332 574186 676437 574196
rect 676320 574180 676437 574186
rect 676372 574168 676437 574180
rect 676320 574122 676372 574128
rect 676320 573636 676372 573642
rect 676372 573584 676437 573610
rect 676320 573582 676437 573584
rect 676320 573578 676372 573582
rect 676228 572344 676280 572350
rect 676228 572286 676280 572292
rect 676240 572202 676437 572230
rect 676240 571534 676268 572202
rect 676228 571528 676280 571534
rect 676228 571470 676280 571476
rect 676240 571386 676360 571414
rect 676240 570650 676268 571386
rect 676332 571317 676360 571386
rect 676332 571289 676437 571317
rect 676320 571188 676372 571194
rect 676320 571130 676372 571136
rect 676228 570644 676280 570650
rect 676228 570586 676280 570592
rect 676332 567921 676360 571130
rect 676332 567893 676437 567921
rect 676240 565754 676437 565770
rect 676228 565748 676437 565754
rect 676280 565742 676437 565748
rect 676228 565690 676280 565696
rect 676226 565580 676282 565589
rect 676226 565515 676282 565524
rect 676240 565056 676268 565515
rect 676320 565408 676372 565414
rect 676320 565351 676372 565356
rect 676320 565350 676437 565351
rect 676332 565323 676437 565350
rect 676332 565192 676360 565323
rect 676332 565164 676452 565192
rect 676320 565068 676372 565074
rect 676240 565028 676320 565056
rect 676320 565010 676372 565016
rect 676228 563436 676280 563442
rect 676228 563378 676280 563384
rect 676240 543722 676268 563378
rect 676228 543716 676280 543722
rect 676228 543658 676280 543664
rect 676332 543654 676360 565010
rect 676424 558886 676452 565164
rect 676596 564592 676648 564598
rect 676596 564534 676648 564540
rect 676504 559016 676556 559022
rect 676504 558958 676556 558964
rect 676412 558880 676464 558886
rect 676412 558822 676464 558828
rect 676320 543648 676372 543654
rect 676320 543590 676372 543596
rect 676516 540526 676544 558958
rect 676504 540520 676556 540526
rect 676504 540462 676556 540468
rect 676608 540458 676636 564534
rect 676688 563844 676740 563850
rect 676688 563786 676740 563792
rect 676700 559022 676728 563786
rect 676688 559016 676740 559022
rect 676688 558958 676740 558964
rect 676688 558880 676740 558886
rect 676688 558822 676740 558828
rect 676700 540594 676728 558822
rect 676688 540588 676740 540594
rect 676688 540530 676740 540536
rect 676596 540452 676648 540458
rect 676596 540394 676648 540400
rect 676136 539704 676188 539710
rect 676136 539646 676188 539652
rect 676320 539704 676372 539710
rect 676320 539646 676372 539652
rect 676332 539616 676360 539646
rect 676332 539588 676437 539616
rect 676136 539500 676188 539506
rect 676136 539442 676188 539448
rect 676148 536038 676176 539442
rect 676228 539228 676280 539234
rect 676280 539179 676437 539207
rect 676228 539170 676280 539176
rect 676240 539062 676268 539170
rect 676240 539034 676437 539062
rect 676240 537845 676268 539034
rect 676226 537836 676282 537845
rect 676226 537771 676282 537780
rect 676320 537737 676372 537738
rect 676320 537732 676437 537737
rect 676226 537700 676282 537709
rect 676372 537709 676437 537732
rect 676320 537674 676372 537680
rect 676226 537635 676282 537644
rect 676240 537058 676268 537635
rect 676228 537052 676280 537058
rect 676228 536994 676280 537000
rect 676320 537052 676372 537058
rect 676372 537000 676437 537026
rect 676320 536998 676437 537000
rect 676320 536994 676372 536998
rect 676240 536213 676268 536994
rect 676320 536848 676372 536854
rect 676320 536790 676372 536796
rect 676226 536204 676282 536213
rect 676226 536139 676282 536148
rect 676332 536122 676360 536790
rect 676322 536077 676360 536122
rect 676308 536068 676364 536077
rect 676136 536032 676188 536038
rect 676308 536003 676364 536012
rect 676136 535974 676188 535980
rect 676148 535890 676360 535918
rect 676148 535290 676176 535890
rect 676332 535817 676360 535890
rect 676332 535789 676437 535817
rect 676136 535284 676188 535290
rect 676136 535226 676188 535232
rect 675872 535040 675992 535068
rect 676044 535080 676096 535086
rect 675766 532532 675822 532541
rect 675766 532467 675822 532476
rect 675768 532428 675820 532434
rect 675768 532370 675820 532376
rect 675676 530252 675728 530258
rect 675676 530194 675728 530200
rect 675674 530084 675730 530093
rect 675674 530019 675730 530028
rect 675688 527810 675716 530019
rect 675676 527804 675728 527810
rect 675676 527746 675728 527752
rect 675780 524766 675808 532370
rect 675872 528634 675900 535040
rect 676044 535022 676096 535028
rect 676226 534980 676282 534989
rect 676044 534944 676096 534950
rect 676282 534938 676437 534966
rect 676226 534915 676282 534924
rect 676044 534886 676096 534892
rect 676056 534270 676084 534886
rect 676228 534604 676280 534610
rect 676280 534562 676437 534590
rect 676228 534546 676280 534552
rect 676044 534264 676096 534270
rect 676044 534206 676096 534212
rect 676226 534152 676282 534161
rect 676044 534128 676096 534134
rect 676282 534110 676437 534138
rect 676226 534087 676282 534096
rect 676044 534070 676096 534076
rect 675952 533924 676004 533930
rect 675952 533866 676004 533872
rect 675964 529646 675992 533866
rect 675952 529640 676004 529646
rect 675952 529582 676004 529588
rect 675872 528606 675992 528634
rect 675780 524738 675900 524766
rect 675584 524676 675636 524682
rect 675584 524618 675636 524624
rect 675766 524644 675822 524653
rect 675766 524579 675822 524588
rect 675780 520330 675808 524579
rect 675872 524002 675900 524738
rect 675860 523996 675912 524002
rect 675860 523938 675912 523944
rect 675768 520324 675820 520330
rect 675768 520266 675820 520272
rect 675768 509308 675820 509314
rect 675768 509250 675820 509256
rect 675492 502712 675544 502718
rect 675492 502654 675544 502660
rect 675400 495504 675452 495510
rect 675400 495446 675452 495452
rect 675308 494212 675360 494218
rect 675308 494154 675360 494160
rect 675320 490381 675348 494154
rect 675412 493130 675440 495446
rect 675400 493124 675452 493130
rect 675400 493066 675452 493072
rect 675504 491634 675532 502654
rect 675780 502106 675808 509250
rect 675860 504888 675912 504894
rect 675860 504830 675912 504836
rect 675768 502100 675820 502106
rect 675768 502042 675820 502048
rect 675768 501624 675820 501630
rect 675768 501566 675820 501572
rect 675676 500468 675728 500474
rect 675676 500410 675728 500416
rect 675584 498904 675636 498910
rect 675584 498846 675636 498852
rect 675596 491838 675624 498846
rect 675688 497722 675716 500410
rect 675780 498774 675808 501566
rect 675768 498768 675820 498774
rect 675768 498710 675820 498716
rect 675688 497694 675808 497722
rect 675780 496938 675808 497694
rect 675768 496932 675820 496938
rect 675768 496874 675820 496880
rect 675676 496252 675728 496258
rect 675676 496194 675728 496200
rect 675688 494218 675716 496194
rect 675676 494212 675728 494218
rect 675676 494154 675728 494160
rect 675676 493804 675728 493810
rect 675676 493746 675728 493752
rect 675688 493334 675716 493746
rect 675676 493328 675728 493334
rect 675676 493270 675728 493276
rect 675584 491832 675636 491838
rect 675584 491774 675636 491780
rect 675492 491628 675544 491634
rect 675492 491570 675544 491576
rect 675306 490372 675362 490381
rect 675306 490307 675362 490316
rect 675596 489994 675624 491774
rect 675504 489966 675624 489994
rect 675504 483610 675532 489966
rect 675688 486126 675716 493270
rect 675780 492246 675808 496874
rect 675872 495510 675900 504830
rect 675860 495504 675912 495510
rect 675860 495446 675912 495452
rect 675860 495368 675912 495374
rect 675860 495310 675912 495316
rect 675768 492240 675820 492246
rect 675768 492182 675820 492188
rect 675872 490478 675900 495310
rect 675860 490472 675912 490478
rect 675860 490414 675912 490420
rect 675768 489452 675820 489458
rect 675768 489394 675820 489400
rect 675676 486120 675728 486126
rect 675676 486062 675728 486068
rect 675492 483604 675544 483610
rect 675492 483546 675544 483552
rect 675504 481570 675532 483546
rect 675780 483474 675808 489394
rect 675860 487004 675912 487010
rect 675860 486946 675912 486952
rect 675872 484018 675900 486946
rect 675860 484012 675912 484018
rect 675860 483954 675912 483960
rect 675768 483468 675820 483474
rect 675768 483410 675820 483416
rect 675872 483406 675900 483954
rect 675860 483400 675912 483406
rect 675860 483342 675912 483348
rect 675492 481564 675544 481570
rect 675492 481506 675544 481512
rect 675964 280222 675992 528606
rect 676056 495374 676084 534070
rect 676320 533925 676372 533930
rect 676320 533924 676437 533925
rect 676372 533897 676437 533924
rect 676320 533866 676372 533872
rect 676136 533244 676188 533250
rect 676188 533192 676437 533196
rect 676136 533186 676437 533192
rect 676148 533168 676437 533186
rect 676148 532434 676176 533168
rect 676320 532632 676372 532638
rect 676372 532582 676437 532610
rect 676320 532574 676372 532580
rect 676136 532428 676188 532434
rect 676136 532370 676188 532376
rect 676148 531211 676437 531239
rect 676148 530870 676176 531211
rect 676136 530864 676188 530870
rect 676136 530806 676188 530812
rect 676148 530289 676437 530317
rect 676148 529782 676176 530289
rect 676320 530252 676372 530258
rect 676320 530194 676372 530200
rect 676136 529776 676188 529782
rect 676136 529718 676188 529724
rect 676136 529640 676188 529646
rect 676136 529582 676188 529588
rect 676148 520414 676176 529582
rect 676228 527804 676280 527810
rect 676228 527746 676280 527752
rect 676240 524766 676268 527746
rect 676332 526921 676360 530194
rect 676332 526893 676437 526921
rect 676240 524738 676437 524766
rect 676240 524120 676268 524738
rect 676320 524676 676372 524682
rect 676320 524618 676372 524624
rect 676332 524351 676360 524618
rect 676332 524323 676437 524351
rect 676332 524222 676360 524323
rect 676332 524194 676728 524222
rect 676240 524092 676360 524120
rect 676228 523996 676280 524002
rect 676228 523938 676280 523944
rect 676240 520550 676268 523938
rect 676332 520670 676360 524092
rect 676594 524100 676650 524109
rect 676594 524035 676650 524044
rect 676320 520664 676372 520670
rect 676320 520606 676372 520612
rect 676240 520522 676544 520550
rect 676412 520460 676464 520466
rect 676148 520386 676268 520414
rect 676412 520402 676464 520408
rect 676136 520324 676188 520330
rect 676136 520266 676188 520272
rect 676148 502718 676176 520266
rect 676240 504894 676268 520386
rect 676228 504888 676280 504894
rect 676228 504830 676280 504836
rect 676136 502712 676188 502718
rect 676136 502654 676188 502660
rect 676228 502712 676280 502718
rect 676228 502654 676280 502660
rect 676136 502168 676188 502174
rect 676136 502110 676188 502116
rect 676148 500474 676176 502110
rect 676136 500468 676188 500474
rect 676136 500410 676188 500416
rect 676136 499992 676188 499998
rect 676136 499934 676188 499940
rect 676148 498298 676176 499934
rect 676240 498910 676268 502654
rect 676320 502100 676372 502106
rect 676320 502042 676372 502048
rect 676332 498978 676360 502042
rect 676424 499998 676452 520402
rect 676516 502174 676544 520522
rect 676504 502168 676556 502174
rect 676504 502110 676556 502116
rect 676608 501630 676636 524035
rect 676700 502718 676728 524194
rect 676688 502712 676740 502718
rect 676688 502654 676740 502660
rect 676596 501624 676648 501630
rect 676596 501566 676648 501572
rect 676412 499992 676464 499998
rect 676412 499934 676464 499940
rect 676320 498972 676372 498978
rect 676320 498914 676372 498920
rect 676228 498904 676280 498910
rect 676228 498846 676280 498852
rect 676320 498836 676372 498842
rect 676372 498788 676437 498816
rect 676320 498778 676372 498784
rect 676228 498768 676280 498774
rect 676228 498710 676280 498716
rect 676136 498292 676188 498298
rect 676136 498234 676188 498240
rect 676148 496258 676176 498234
rect 676136 496252 676188 496258
rect 676136 496194 676188 496200
rect 676044 495368 676096 495374
rect 676044 495310 676096 495316
rect 676240 495254 676268 498710
rect 676320 498428 676372 498434
rect 676372 498379 676437 498407
rect 676320 498370 676372 498376
rect 676320 498292 676372 498298
rect 676372 498240 676437 498262
rect 676320 498234 676437 498240
rect 676320 496937 676372 496938
rect 676320 496932 676437 496937
rect 676372 496909 676437 496932
rect 676320 496874 676372 496880
rect 676320 496252 676372 496258
rect 676372 496200 676437 496226
rect 676320 496198 676437 496200
rect 676320 496194 676372 496198
rect 676056 495226 676268 495254
rect 676056 491718 676084 495226
rect 676136 495164 676188 495170
rect 676136 495106 676188 495112
rect 676148 495017 676176 495106
rect 676148 494989 676437 495017
rect 676228 494212 676280 494218
rect 676280 494160 676437 494166
rect 676228 494154 676437 494160
rect 676240 494138 676437 494154
rect 676240 493452 676268 494138
rect 676320 493804 676372 493810
rect 676372 493762 676437 493790
rect 676320 493746 676372 493752
rect 676240 493424 676360 493452
rect 676332 493350 676360 493424
rect 676332 493322 676437 493350
rect 676320 493125 676372 493130
rect 676320 493124 676437 493125
rect 676372 493097 676437 493124
rect 676320 493066 676372 493072
rect 676148 492370 676437 492398
rect 676148 492246 676176 492370
rect 676136 492240 676188 492246
rect 676136 492182 676188 492188
rect 676320 491832 676372 491838
rect 676372 491782 676437 491810
rect 676320 491774 676372 491780
rect 676056 491690 676268 491718
rect 676136 491628 676188 491634
rect 676136 491570 676188 491576
rect 676042 490322 676098 490331
rect 676042 490257 676098 490266
rect 676056 487010 676084 490257
rect 676044 487004 676096 487010
rect 676044 486946 676096 486952
rect 676148 486437 676176 491570
rect 676134 486428 676190 486437
rect 676134 486363 676190 486372
rect 676240 486278 676268 491690
rect 676320 490472 676372 490478
rect 676372 490420 676437 490439
rect 676320 490414 676437 490420
rect 676332 490411 676437 490414
rect 676332 489489 676437 489517
rect 676332 489458 676360 489489
rect 676320 489452 676372 489458
rect 676320 489394 676372 489400
rect 676056 486250 676268 486278
rect 676056 481706 676084 486250
rect 676320 486121 676372 486126
rect 676320 486120 676437 486121
rect 676372 486093 676437 486120
rect 676320 486062 676372 486068
rect 676320 484012 676372 484018
rect 676372 483960 676437 483966
rect 676320 483954 676437 483960
rect 676332 483938 676437 483954
rect 676228 483604 676280 483610
rect 676228 483551 676280 483552
rect 676228 483546 676437 483551
rect 676240 483523 676437 483546
rect 676228 483468 676280 483474
rect 676134 483436 676190 483445
rect 676228 483410 676280 483416
rect 676134 483371 676190 483380
rect 676044 481700 676096 481706
rect 676044 481642 676096 481648
rect 676044 481564 676096 481570
rect 676044 481506 676096 481512
rect 675952 280216 676004 280222
rect 675952 280158 676004 280164
rect 675216 279740 675268 279746
rect 675216 279682 675268 279688
rect 673312 277908 673318 277960
rect 673370 277908 673376 277960
rect 659760 259690 659812 259696
rect 660862 259716 660918 259725
rect 656400 259651 656456 259660
rect 657722 259680 657774 259686
rect 655686 259622 655738 259628
rect 655698 259470 655726 259622
rect 656414 259470 656442 259651
rect 657722 259622 657774 259628
rect 657828 259680 657880 259686
rect 676056 259686 676084 481506
rect 676148 279134 676176 483371
rect 676240 475450 676268 483410
rect 676576 481700 676628 481706
rect 676576 481642 676628 481648
rect 676228 475444 676280 475450
rect 676228 475386 676280 475392
rect 676588 423754 676616 481642
rect 676312 423726 676616 423754
rect 676312 400570 676340 423726
rect 676312 400542 676616 400570
rect 676588 385114 676616 400542
rect 676292 385086 676616 385114
rect 676292 361930 676320 385086
rect 676292 361902 676616 361930
rect 676588 300106 676616 361902
rect 676312 300078 676616 300106
rect 676136 279128 676188 279134
rect 676136 279070 676188 279076
rect 676312 279066 676340 300078
rect 676300 279060 676352 279066
rect 676300 279002 676352 279008
rect 660862 259651 660918 259660
rect 676044 259680 676096 259686
rect 657828 259622 657880 259628
rect 676044 259622 676096 259628
rect 657734 259566 657762 259622
rect 658276 259612 658328 259618
rect 657734 259538 657907 259566
rect 658276 259554 658328 259560
rect 657734 259470 657762 259538
rect 657879 259470 657907 259538
rect 658288 259470 658316 259554
rect 577602 259439 577658 259448
rect 414856 259340 414908 259346
rect 414856 259282 414908 259288
<< via2 >>
rect 208130 715729 208186 715785
rect 208222 715559 208278 715615
rect 208130 714793 208186 714849
rect 208130 711413 208186 711469
rect 208130 709078 208186 709134
rect 208866 709004 208922 709060
rect 208130 704729 208186 704785
rect 208222 702952 208278 703008
rect 208222 700237 208278 700293
rect 208222 699147 208278 699203
rect 209970 707236 210026 707292
rect 209970 703292 210026 703348
rect 209970 699076 210026 699132
rect 208866 698668 208922 698724
rect 208222 695376 208278 695432
rect 208130 694331 208186 694387
rect 208130 693833 208186 693889
rect 208314 691732 208370 691788
rect 208222 691529 208278 691585
rect 208222 691113 208278 691169
rect 209970 695404 210026 695460
rect 208222 676329 208278 676385
rect 208866 676364 208922 676420
rect 208130 676161 208186 676217
rect 208130 675534 208186 675590
rect 208222 675393 208278 675449
rect 208130 672185 208186 672241
rect 208130 672012 208186 672068
rect 208130 669673 208186 669729
rect 208314 672185 208370 672241
rect 208314 668038 208370 668094
rect 208314 667868 208370 667924
rect 208222 665331 208278 665387
rect 208130 663893 208186 663949
rect 208130 660837 208186 660893
rect 208130 659746 208186 659802
rect 208130 655976 208186 656032
rect 209326 691732 209382 691788
rect 209970 691052 210026 691108
rect 208130 654933 208186 654989
rect 208866 654332 208922 654388
rect 208130 652312 208186 652316
rect 208130 652260 208132 652312
rect 208132 652260 208184 652312
rect 208184 652260 208186 652312
rect 208130 652127 208186 652183
rect 208130 651663 208186 651719
rect 208222 638964 208278 639020
rect 208406 638828 208462 638884
rect 208958 651612 209014 651668
rect 208038 628220 208094 628276
rect 208038 625649 208094 625705
rect 208222 625636 208278 625692
rect 208590 625636 208646 625692
rect 208038 623770 208094 623826
rect 208498 611593 208554 611649
rect 208314 611471 208370 611527
rect 208038 605669 208094 605725
rect 208222 604828 208278 604884
rect 208224 604673 208280 604729
rect 208038 603376 208094 603432
rect 208038 602061 208094 602117
rect 208958 632164 209014 632220
rect 208958 623732 209014 623788
rect 208682 609180 208738 609236
rect 208498 602108 208554 602164
rect 208038 600169 208094 600225
rect 208038 596370 208094 596426
rect 208406 596396 208462 596452
rect 208314 584020 208370 584076
rect 208038 575976 208094 576032
rect 208038 575384 208094 575440
rect 208314 575316 208370 575372
rect 208038 574448 208094 574504
rect 208038 573996 208094 574052
rect 208498 575996 208554 576052
rect 208406 573956 208462 574012
rect 208038 571560 208094 571616
rect 208038 556621 208094 556677
rect 208866 577356 208922 577412
rect 208130 550078 208186 550134
rect 208866 574500 208922 574556
rect 208866 571508 208922 571564
rect 210062 659364 210118 659420
rect 209784 658153 210076 658661
rect 209142 655964 209198 656020
rect 209326 612988 209382 613044
rect 208038 546756 208094 546812
rect 208038 546484 208094 546540
rect 208038 545369 208094 545425
rect 208038 544172 208094 544228
rect 208038 543449 208094 543505
rect 208038 541570 208094 541626
rect 208038 529484 208094 529540
rect 208774 544172 208830 544228
rect 208590 543492 208646 543548
rect 208498 541588 208554 541644
rect 208038 526865 208094 526921
rect 208682 529222 208738 529278
rect 208222 522548 208278 522604
rect 208498 522548 208554 522604
rect 208038 519420 208094 519476
rect 208038 518808 208094 518864
rect 208314 518876 208370 518932
rect 208682 526900 208738 526956
rect 208038 516049 208094 516105
rect 208314 516020 208370 516076
rect 208682 519420 208738 519476
rect 208094 501950 208150 502006
rect 208498 501821 208554 501877
rect 208038 499465 208094 499521
rect 208038 496069 208094 496125
rect 208682 499428 208738 499484
rect 208406 495076 208462 495132
rect 208038 493172 208094 493228
rect 208038 492461 208094 492517
rect 208682 496028 208738 496084
rect 208682 495076 208738 495132
rect 208590 493264 208646 493320
rect 208038 486770 208094 486826
rect 208866 496028 208922 496084
rect 208774 492492 208830 492548
rect 208866 486780 208922 486836
rect 208590 474132 208646 474188
rect 208866 474132 208922 474188
rect 208038 461756 208094 461812
rect 208038 459724 208094 459780
rect 208038 459580 208094 459636
rect 208130 459040 208186 459096
rect 209050 467876 209106 467932
rect 208590 459580 208646 459636
rect 208682 459308 208738 459364
rect 208866 461756 208922 461812
rect 208866 459580 208922 459636
rect 208038 441069 208094 441125
rect 208222 440278 208278 440334
rect 208038 438776 208094 438832
rect 208590 446796 208646 446852
rect 209080 457810 209136 457866
rect 208406 438772 208462 438828
rect 208590 441084 208646 441140
rect 208038 431768 208094 431824
rect 208774 440278 208830 440334
rect 208682 431700 208738 431756
rect 208866 431700 208922 431756
rect 208866 393076 208922 393132
rect 208130 386478 208186 386534
rect 208038 383661 208094 383717
rect 208498 383692 208554 383748
rect 210154 655148 210210 655204
rect 209418 555596 209474 555652
rect 209694 584156 209750 584212
rect 226265 692383 226757 692698
rect 220076 667552 222120 667728
rect 236536 665954 242984 667020
rect 213466 654604 213522 654660
rect 211534 623732 211590 623788
rect 211534 556684 211590 556740
rect 211166 474540 211222 474596
rect 210430 447068 210486 447124
rect 231222 284684 231278 284740
rect 244654 599524 244710 599580
rect 244654 557092 244710 557148
rect 233614 284684 233670 284740
rect 232234 283732 232290 283788
rect 226990 280468 227046 280524
rect 230210 280468 230266 280524
rect 232326 279924 232382 279980
rect 240238 280060 240294 280116
rect 244654 279924 244710 279980
rect 246793 542964 246889 543064
rect 246862 500244 246918 500300
rect 247414 613668 247470 613724
rect 247322 436596 247378 436652
rect 246310 316100 246366 316156
rect 248058 550020 248114 550076
rect 248978 493172 249034 493228
rect 249254 415380 249310 415436
rect 249346 358532 249402 358588
rect 250082 585380 250138 585436
rect 250082 386820 250138 386876
rect 250726 699076 250782 699132
rect 250266 400964 250322 401020
rect 250450 648348 250506 648404
rect 250358 365604 250414 365660
rect 250818 514388 250874 514444
rect 250818 479028 250874 479084
rect 250818 422452 250874 422508
rect 251002 521460 251058 521516
rect 251094 464884 251150 464940
rect 251278 393892 251334 393948
rect 251830 627812 251886 627868
rect 252014 606596 252070 606652
rect 252014 535604 252070 535660
rect 251922 337316 251978 337372
rect 252382 620740 252438 620796
rect 252382 606596 252438 606652
rect 252290 486100 252346 486156
rect 252198 471956 252254 472012
rect 252566 642228 252622 642284
rect 252474 507588 252530 507644
rect 252382 443668 252438 443724
rect 252106 429524 252162 429580
rect 252106 351460 252162 351516
rect 252658 344660 252714 344716
rect 252290 330244 252346 330300
rect 252198 323172 252254 323228
rect 252198 309028 252254 309084
rect 252382 294884 252438 294940
rect 252290 280468 252346 280524
rect 254406 646852 254462 646908
rect 286606 698804 286662 698860
rect 279890 687380 279946 687436
rect 279982 681396 280038 681452
rect 286422 671060 286478 671116
rect 314942 699892 314998 699948
rect 288538 699756 288594 699812
rect 288262 695132 288318 695188
rect 288170 679084 288226 679140
rect 288078 676908 288134 676964
rect 287986 674732 288042 674788
rect 287894 672828 287950 672884
rect 288446 693228 288502 693284
rect 288538 686156 288594 686212
rect 288538 682892 288594 682948
rect 298382 699212 298438 699268
rect 301694 699212 301750 699268
rect 291482 698940 291538 698996
rect 290010 698804 290066 698860
rect 306846 699212 306902 699268
rect 310802 699076 310858 699132
rect 312090 698804 312146 698860
rect 313562 698804 313618 698860
rect 319082 698804 319138 698860
rect 289090 698668 289146 698724
rect 288814 691052 288870 691108
rect 288722 690508 288778 690564
rect 288630 682348 288686 682404
rect 288630 681396 288686 681452
rect 289090 668748 289146 668804
rect 289366 666744 289368 666764
rect 289368 666744 289420 666764
rect 289420 666744 289422 666764
rect 289366 666708 289422 666744
rect 290838 667252 290894 667308
rect 311354 667252 311410 667308
rect 311538 667252 311594 667308
rect 257902 646852 257958 646908
rect 258546 646852 258602 646908
rect 259190 646852 259246 646908
rect 278510 646852 278566 646908
rect 279982 646852 280038 646908
rect 287250 646852 287306 646908
rect 288078 646852 288134 646908
rect 301602 667116 301658 667172
rect 308226 667136 308282 667172
rect 308226 667116 308228 667136
rect 308228 667116 308280 667136
rect 308280 667116 308282 667136
rect 308594 667116 308650 667172
rect 307122 666844 307178 666900
rect 311538 648484 311594 648540
rect 320646 695948 320702 696004
rect 320646 691324 320702 691380
rect 320646 686292 320702 686348
rect 320646 684116 320702 684172
rect 322578 700028 322634 700084
rect 321014 698940 321070 698996
rect 320830 694180 320886 694236
rect 320738 676908 320794 676964
rect 320738 673644 320794 673700
rect 320922 691868 320978 691924
rect 321106 684116 321162 684172
rect 321014 680988 321070 681044
rect 321014 669564 321070 669620
rect 321198 677724 321254 677780
rect 321290 671604 321346 671660
rect 323682 698804 323738 698860
rect 325246 667388 325302 667444
rect 325246 666572 325302 666628
rect 341500 669822 341796 670342
rect 343162 669782 343450 670294
rect 301602 646852 301658 646908
rect 302430 646852 302486 646908
rect 315954 646852 316010 646908
rect 316782 646852 316838 646908
rect 356748 729268 356804 729324
rect 361034 729268 361090 729324
rect 365634 728860 365690 728916
rect 356986 693500 357042 693556
rect 367658 728996 367714 729052
rect 368026 728860 368082 728916
rect 386978 729424 387034 729426
rect 386978 729372 386980 729424
rect 386980 729372 387032 729424
rect 387032 729372 387034 729424
rect 386978 729370 387034 729372
rect 392222 728996 392278 729052
rect 394522 728996 394578 729052
rect 379066 700028 379122 700084
rect 360666 684932 360722 684988
rect 359838 681940 359894 681996
rect 360758 673508 360814 673564
rect 361126 666980 361182 667036
rect 361310 666980 361366 667036
rect 367106 698668 367162 698724
rect 385138 699892 385194 699948
rect 381090 699756 381146 699812
rect 370786 694588 370842 694644
rect 371154 694588 371210 694644
rect 375018 694588 375074 694644
rect 375202 694588 375258 694644
rect 365082 694452 365138 694508
rect 383114 694452 383170 694508
rect 362874 690508 362930 690564
rect 362414 687516 362470 687572
rect 362322 675548 362378 675604
rect 362506 684932 362562 684988
rect 362598 678948 362654 679004
rect 362690 673508 362746 673564
rect 390290 689148 390346 689204
rect 390382 687108 390438 687164
rect 365266 664940 365322 664996
rect 381090 667136 381146 667172
rect 381090 667116 381092 667136
rect 381092 667116 381144 667136
rect 381144 667116 381146 667136
rect 381274 667116 381330 667172
rect 385322 666436 385378 666492
rect 390290 680172 390346 680228
rect 390658 677724 390714 677780
rect 390290 674188 390346 674244
rect 390198 667252 390254 667308
rect 390474 671468 390530 671524
rect 390382 668884 390438 668940
rect 390382 666844 390438 666900
rect 344658 646852 344714 646908
rect 345486 646852 345542 646908
rect 410116 729268 410172 729324
rect 410948 729268 411004 729324
rect 414302 729268 414358 729324
rect 420190 729404 420246 729460
rect 419914 729268 419970 729324
rect 438148 729268 438204 729324
rect 441258 729268 441314 729324
rect 447698 729268 447754 729324
rect 448066 728996 448122 729052
rect 417338 647260 417394 647316
rect 446226 647124 446282 647180
rect 468582 729268 468638 729324
rect 474930 729268 474986 729324
rect 476402 728996 476458 729052
rect 495446 729268 495502 729324
rect 501610 729404 501666 729460
rect 501426 728996 501482 729052
rect 522678 729268 522734 729324
rect 529118 729268 529174 729324
rect 529210 728996 529266 729052
rect 546736 729268 546792 729324
rect 553038 729268 553094 729324
rect 554694 729132 554750 729188
rect 556258 729132 556314 729188
rect 577050 729268 577106 729324
rect 578430 728996 578486 729052
rect 583582 728860 583638 728916
rect 600948 729288 601004 729324
rect 600948 729268 600950 729288
rect 600950 729268 601002 729288
rect 601002 729268 601004 729288
rect 604769 729268 604825 729324
rect 608165 729304 608167 729324
rect 608167 729304 608219 729324
rect 608219 729304 608221 729324
rect 608165 729268 608221 729304
rect 611458 729268 611514 729324
rect 612194 651476 612250 651532
rect 612378 651612 612434 651668
rect 612286 650796 612342 650852
rect 614402 651884 614458 651940
rect 616794 651748 616850 651804
rect 402066 646852 402122 646908
rect 403078 646852 403134 646908
rect 474286 646852 474342 646908
rect 475022 646852 475078 646908
rect 512466 646852 512522 646908
rect 513294 646852 513350 646908
rect 536754 646852 536810 646908
rect 537398 646852 537454 646908
rect 541170 646852 541226 646908
rect 542182 646852 542238 646908
rect 569874 646852 569930 646908
rect 570886 646852 570942 646908
rect 584226 646852 584282 646908
rect 585238 646852 585294 646908
rect 598578 646852 598634 646908
rect 599590 646852 599646 646908
rect 612930 646852 612986 646908
rect 613942 646852 613998 646908
rect 617898 646852 617954 646908
rect 618726 646852 618782 646908
rect 619094 624412 619150 624468
rect 619094 621284 619150 621340
rect 619094 611764 619150 611820
rect 619094 611628 619150 611684
rect 619094 610676 619150 610732
rect 619094 551244 619150 551300
rect 619370 605372 619426 605428
rect 619462 604148 619518 604204
rect 619370 603876 619426 603932
rect 619370 583748 619426 583804
rect 619278 583476 619334 583532
rect 619278 575316 619334 575372
rect 619370 571916 619426 571972
rect 619278 541996 619334 542052
rect 619186 526900 619242 526956
rect 619094 519828 619150 519884
rect 619462 504868 619518 504924
rect 619094 490180 619150 490236
rect 276854 279652 276910 279708
rect 396638 279788 396694 279844
rect 478150 278972 478206 279028
rect 384310 259680 384366 259736
rect 384494 259680 384550 259736
rect 388375 259696 388377 259716
rect 388377 259696 388429 259716
rect 388429 259696 388431 259716
rect 388375 259660 388431 259696
rect 392196 259660 392252 259716
rect 392636 259660 392692 259716
rect 393026 259660 393082 259716
rect 393875 259660 393931 259716
rect 395074 259660 395130 259716
rect 414854 259660 414910 259716
rect 415424 259660 415480 259716
rect 417579 259660 417635 259716
rect 420972 259660 421028 259716
rect 424790 259660 424846 259716
rect 425248 259660 425304 259716
rect 425618 259660 425674 259716
rect 426446 259660 426502 259716
rect 446318 259660 446374 259716
rect 451010 259660 451066 259716
rect 454414 259584 454470 259640
rect 480266 259660 480322 259716
rect 482579 259696 482581 259716
rect 482581 259696 482633 259716
rect 482633 259696 482635 259716
rect 482579 259660 482635 259696
rect 485970 259660 486026 259716
rect 489788 259660 489844 259716
rect 490248 259660 490304 259716
rect 490616 259660 490672 259716
rect 491475 259660 491531 259716
rect 492684 259660 492740 259716
rect 494710 259660 494766 259716
rect 512834 259660 512890 259716
rect 516146 259716 516148 259736
rect 516148 259716 516200 259736
rect 516200 259716 516202 259736
rect 516146 259680 516202 259716
rect 518538 259660 518594 259716
rect 522402 259660 522458 259716
rect 545034 259588 545090 259644
rect 551175 259660 551231 259716
rect 554996 259680 555052 259716
rect 554996 259660 554998 259680
rect 554998 259660 555050 259680
rect 555050 259660 555052 259680
rect 619186 406404 619242 406460
rect 620014 636652 620070 636708
rect 620014 632028 620070 632084
rect 620014 597076 620070 597132
rect 620014 547572 620070 547628
rect 619922 292436 619978 292492
rect 620106 469508 620162 469564
rect 620198 441220 620254 441276
rect 620198 420004 620254 420060
rect 620198 370228 620254 370284
rect 620106 313652 620162 313708
rect 577602 259448 577658 259504
rect 578062 259660 578118 259716
rect 580822 259660 580878 259716
rect 583775 259680 583831 259716
rect 583775 259660 583777 259680
rect 583777 259660 583829 259680
rect 583829 259660 583831 259680
rect 584502 259660 584558 259716
rect 587584 259660 587640 259716
rect 588044 259660 588100 259716
rect 588426 259660 588482 259716
rect 590482 259660 590538 259716
rect 621486 632164 621542 632220
rect 621394 497796 621450 497852
rect 621210 427076 621266 427132
rect 621026 384372 621082 384428
rect 620934 341940 620990 341996
rect 620842 334868 620898 334924
rect 631238 729268 631294 729324
rect 631974 729268 632030 729324
rect 637218 728996 637274 729052
rect 609710 259932 609766 259988
rect 610630 259796 610686 259852
rect 622590 561716 622646 561772
rect 622406 462436 622462 462492
rect 622314 412932 622370 412988
rect 622222 349012 622278 349068
rect 622130 320724 622186 320780
rect 623418 568788 623474 568844
rect 623326 455364 623382 455420
rect 623234 434148 623290 434204
rect 623142 398788 623198 398844
rect 627742 647260 627798 647316
rect 615598 259660 615654 259716
rect 620198 259660 620254 259716
rect 621026 259660 621082 259716
rect 623084 259660 623140 259716
rect 625120 259660 625176 259716
rect 637678 729268 637734 729324
rect 652460 729268 652516 729324
rect 654518 729268 654574 729324
rect 655348 729268 655404 729324
rect 634944 280890 636264 281126
rect 639518 650524 639574 650580
rect 632526 259660 632582 259716
rect 642326 280712 643110 280916
rect 659169 729268 659225 729324
rect 662565 729304 662567 729324
rect 662567 729304 662619 729324
rect 662619 729304 662621 729324
rect 662565 729268 662621 729304
rect 664818 729268 664874 729324
rect 666750 647396 666806 647452
rect 669694 606188 669750 606244
rect 670798 565388 670854 565444
rect 676134 694488 676136 694508
rect 676136 694488 676188 694508
rect 676188 694488 676190 694508
rect 676134 694452 676190 694488
rect 675950 687924 676006 687980
rect 675582 653788 675638 653844
rect 675214 646852 675270 646908
rect 640254 259524 640310 259580
rect 649638 259558 649694 259614
rect 651854 259696 651856 259716
rect 651856 259696 651908 259716
rect 651908 259696 651910 259716
rect 651854 259660 651910 259696
rect 656400 259660 656456 259716
rect 674202 524316 674258 524372
rect 674110 280468 674166 280524
rect 676134 687788 676190 687844
rect 676134 666028 676190 666084
rect 676134 653788 676190 653844
rect 675306 612988 675362 613044
rect 675582 606324 675638 606380
rect 676134 647124 676190 647180
rect 676042 646988 676098 647044
rect 676686 581572 676742 581628
rect 676594 581436 676650 581492
rect 675490 573956 675546 574012
rect 675398 572188 675454 572244
rect 675766 574772 675822 574828
rect 675858 572188 675914 572244
rect 676226 565524 676282 565580
rect 676226 537780 676282 537836
rect 676226 537644 676282 537700
rect 676226 536148 676282 536204
rect 676308 536012 676364 536068
rect 675766 532476 675822 532532
rect 675674 530028 675730 530084
rect 676226 534924 676282 534980
rect 676226 534096 676282 534152
rect 675766 524588 675822 524644
rect 675306 490316 675362 490372
rect 676594 524044 676650 524100
rect 676042 490266 676098 490322
rect 676134 486372 676190 486428
rect 676134 483380 676190 483436
rect 660862 259660 660918 259716
<< obsm2 >>
rect 519318 259446 519378 259450
<< metal3 >>
rect 210508 736476 215394 736602
rect 210508 735934 210592 736476
rect 215276 735934 215394 736476
rect 210508 733110 215394 735934
rect 210508 732568 210598 733110
rect 215282 732568 215394 733110
rect 210508 732456 215394 732568
rect 219899 721784 224679 729560
rect 229878 721784 234658 729560
rect 246100 721784 250900 730190
rect 256151 721784 260940 730190
rect 219899 718852 260940 721784
rect 219899 718282 260888 718852
rect 208125 715787 208191 715790
rect 207928 715785 208191 715787
rect 207928 715729 208130 715785
rect 208186 715729 208191 715785
rect 207928 715727 208191 715729
rect 208125 715724 208191 715727
rect 208217 715617 208283 715620
rect 207928 715615 208283 715617
rect 207928 715559 208222 715615
rect 208278 715559 208283 715615
rect 207928 715557 208283 715559
rect 208217 715554 208283 715557
rect 207928 714930 208050 714990
rect 207990 714851 208050 714930
rect 208125 714851 208191 714854
rect 207928 714849 208191 714851
rect 207928 714793 208130 714849
rect 208186 714793 208191 714849
rect 207928 714791 208191 714793
rect 208125 714788 208191 714791
rect 207928 711581 208050 711641
rect 207990 711471 208050 711581
rect 208125 711471 208191 711474
rect 207928 711469 208191 711471
rect 207928 711413 208130 711469
rect 208186 711413 208191 711469
rect 207928 711411 208191 711413
rect 208125 711408 208191 711411
rect 208125 709136 208191 709139
rect 207928 709134 208602 709136
rect 207928 709078 208130 709134
rect 208186 709078 208602 709134
rect 207928 709076 208602 709078
rect 208125 709073 208191 709076
rect 208542 709062 208602 709076
rect 208861 709062 208927 709065
rect 208542 709060 208927 709062
rect 208542 709004 208866 709060
rect 208922 709004 208927 709060
rect 208542 709002 208927 709004
rect 208861 708999 208927 709002
rect 207928 707435 208188 707495
rect 208128 707325 208188 707435
rect 207928 707294 208188 707325
rect 209965 707294 210031 707297
rect 207928 707292 210031 707294
rect 207928 707265 209970 707292
rect 208128 707236 209970 707265
rect 210026 707236 210031 707292
rect 208128 707234 210031 707236
rect 209965 707231 210031 707234
rect 208125 704787 208191 704790
rect 207928 704785 208191 704787
rect 207928 704729 208130 704785
rect 208186 704729 208191 704785
rect 207928 704727 208191 704729
rect 208125 704724 208191 704727
rect 209965 703350 210031 703353
rect 207928 703348 210031 703350
rect 207928 703292 209970 703348
rect 210026 703292 210031 703348
rect 207928 703290 210031 703292
rect 208128 703181 208188 703290
rect 209965 703287 210031 703290
rect 207928 703121 208418 703181
rect 208217 703010 208283 703013
rect 208358 703010 208418 703121
rect 207928 703008 208418 703010
rect 207928 702952 208222 703008
rect 208278 702952 208418 703008
rect 207928 702950 208418 702952
rect 208217 702947 208283 702950
rect 208217 700295 208283 700298
rect 207928 700293 208283 700295
rect 207928 700237 208222 700293
rect 208278 700237 208283 700293
rect 207928 700235 208283 700237
rect 208217 700232 208283 700235
rect 208217 699205 208283 699208
rect 207928 699203 208602 699205
rect 207928 699147 208222 699203
rect 208278 699147 208602 699203
rect 207928 699145 208602 699147
rect 208217 699142 208283 699145
rect 208542 699134 208602 699145
rect 209965 699134 210031 699137
rect 208542 699132 210031 699134
rect 208542 699076 209970 699132
rect 210026 699076 210031 699132
rect 208542 699074 210031 699076
rect 209965 699071 210031 699074
rect 207928 698974 208188 699034
rect 208128 698770 208188 698974
rect 207928 698726 208188 698770
rect 208861 698726 208927 698729
rect 207928 698724 208927 698726
rect 207928 698710 208866 698724
rect 208128 698668 208866 698710
rect 208922 698668 208927 698724
rect 208128 698666 208927 698668
rect 208861 698663 208927 698666
rect 209965 695462 210031 695465
rect 208358 695460 210031 695462
rect 208217 695434 208283 695437
rect 208358 695434 209970 695460
rect 207928 695432 209970 695434
rect 207928 695376 208222 695432
rect 208278 695404 209970 695432
rect 210026 695404 210031 695460
rect 208278 695402 210031 695404
rect 208278 695376 208418 695402
rect 209965 695399 210031 695402
rect 207928 695374 208418 695376
rect 208217 695371 208283 695374
rect 208125 694389 208191 694392
rect 207928 694387 208191 694389
rect 207928 694331 208130 694387
rect 208186 694331 208191 694387
rect 207928 694329 208191 694331
rect 208125 694326 208191 694329
rect 208125 693891 208191 693894
rect 207928 693889 208191 693891
rect 207928 693833 208130 693889
rect 208186 693833 208191 693889
rect 207928 693831 208191 693833
rect 208125 693828 208191 693831
rect 226248 692698 226784 718282
rect 229878 718254 234658 718282
rect 272299 714638 277079 730190
rect 272299 708222 272398 714638
rect 276856 708222 277079 714638
rect 272299 707726 277079 708222
rect 282278 714662 287058 730190
rect 298299 724720 303079 730190
rect 298299 718358 298404 724720
rect 302880 718358 303079 724720
rect 298299 717846 303079 718358
rect 308278 724748 313058 730190
rect 308278 718386 308406 724748
rect 312882 718386 313058 724748
rect 308278 717846 313058 718386
rect 324500 724586 328760 730190
rect 324500 718358 324690 724586
rect 328652 718358 328760 724586
rect 324500 717846 328760 718358
rect 335042 724614 339340 730190
rect 359773 729456 359850 729508
rect 356743 729326 356809 729329
rect 359790 729326 359850 729456
rect 361029 729326 361095 729329
rect 356743 729324 361095 729326
rect 356743 729268 356748 729324
rect 356804 729268 361034 729324
rect 361090 729268 361095 729324
rect 356743 729266 361095 729268
rect 356743 729263 356809 729266
rect 361029 729263 361095 729266
rect 365629 728918 365695 728921
rect 366319 728918 366379 729553
rect 366451 729054 366511 729553
rect 386976 729431 387036 729553
rect 386973 729426 387039 729431
rect 386973 729370 386978 729426
rect 387034 729370 387039 729426
rect 386973 729365 387039 729370
rect 367653 729054 367719 729057
rect 366451 729052 367719 729054
rect 366451 728996 367658 729052
rect 367714 728996 367719 729052
rect 366451 728994 367719 728996
rect 367653 728991 367719 728994
rect 392217 729054 392283 729057
rect 393519 729054 393579 729553
rect 392217 729052 393579 729054
rect 392217 728996 392222 729052
rect 392278 728996 393579 729052
rect 392217 728994 393579 728996
rect 393646 729054 393706 729553
rect 410111 729326 410177 729329
rect 410943 729326 411009 729329
rect 413976 729326 414036 729553
rect 420185 729462 420251 729465
rect 420516 729462 420576 729553
rect 420651 729493 420754 729553
rect 420185 729460 420576 729462
rect 420185 729404 420190 729460
rect 420246 729404 420576 729460
rect 420185 729402 420576 729404
rect 420185 729399 420251 729402
rect 414297 729326 414363 729329
rect 410111 729324 414363 729326
rect 410111 729268 410116 729324
rect 410172 729268 410948 729324
rect 411004 729268 414302 729324
rect 414358 729268 414363 729324
rect 410111 729266 414363 729268
rect 410111 729263 410177 729266
rect 410943 729263 411009 729266
rect 414297 729263 414363 729266
rect 419909 729326 419975 729329
rect 420694 729326 420754 729493
rect 441176 729329 441236 729553
rect 447716 729453 447782 729566
rect 447696 729389 447782 729453
rect 447696 729329 447756 729389
rect 419909 729324 420754 729326
rect 419909 729268 419914 729324
rect 419970 729268 420754 729324
rect 419909 729266 420754 729268
rect 438143 729326 438209 729329
rect 441176 729326 441319 729329
rect 438143 729324 441319 729326
rect 438143 729268 438148 729324
rect 438204 729268 441258 729324
rect 441314 729268 441319 729324
rect 438143 729266 441319 729268
rect 419909 729263 419975 729266
rect 438143 729263 438209 729266
rect 441253 729263 441319 729266
rect 447693 729324 447759 729329
rect 447693 729268 447698 729324
rect 447754 729268 447759 729324
rect 447693 729263 447759 729268
rect 394517 729054 394583 729057
rect 393646 729052 394583 729054
rect 393646 728996 394522 729052
rect 394578 728996 394583 729052
rect 393646 728994 394583 728996
rect 447851 729054 447911 729553
rect 468373 729422 468439 729566
rect 468350 729326 468439 729422
rect 474919 729329 474979 729553
rect 468577 729326 468643 729329
rect 468350 729324 468643 729326
rect 468350 729268 468582 729324
rect 468638 729268 468643 729324
rect 468350 729266 468643 729268
rect 474919 729324 474991 729329
rect 474919 729268 474930 729324
rect 474986 729268 474991 729324
rect 474919 729266 474991 729268
rect 468577 729263 468643 729266
rect 474925 729263 474991 729266
rect 448061 729054 448127 729057
rect 447851 729052 448127 729054
rect 447851 728996 448066 729052
rect 448122 728996 448127 729052
rect 447851 728994 448127 728996
rect 475051 729054 475111 729553
rect 495373 729460 495439 729566
rect 501916 729468 501982 729566
rect 502047 729493 502266 729553
rect 501605 729462 501671 729465
rect 501817 729462 501982 729468
rect 501605 729460 501982 729462
rect 495373 729402 495458 729460
rect 495398 729329 495458 729402
rect 501605 729404 501610 729460
rect 501666 729404 501982 729460
rect 501605 729402 501982 729404
rect 501605 729399 501671 729402
rect 495398 729324 495507 729329
rect 502206 729326 502266 729493
rect 495398 729268 495446 729324
rect 495502 729268 495507 729324
rect 495398 729266 495507 729268
rect 495441 729263 495507 729266
rect 502022 729266 502266 729326
rect 522576 729329 522636 729553
rect 529119 729329 529179 729553
rect 522576 729324 522739 729329
rect 522576 729268 522678 729324
rect 522734 729268 522739 729324
rect 522576 729266 522739 729268
rect 476397 729054 476463 729057
rect 475051 729052 476463 729054
rect 475051 728996 476402 729052
rect 476458 728996 476463 729052
rect 475051 728994 476463 728996
rect 392217 728991 392283 728994
rect 394517 728991 394583 728994
rect 448061 728991 448127 728994
rect 476397 728991 476463 728994
rect 501421 729054 501487 729057
rect 502022 729054 502082 729266
rect 522673 729263 522739 729266
rect 529113 729324 529179 729329
rect 529113 729268 529118 729324
rect 529174 729268 529179 729324
rect 529113 729263 529179 729268
rect 529254 729057 529314 729553
rect 546731 729326 546797 729329
rect 549776 729326 549836 729553
rect 553033 729326 553099 729329
rect 546731 729324 553099 729326
rect 546731 729268 546736 729324
rect 546792 729268 553038 729324
rect 553094 729268 553099 729324
rect 546731 729266 553099 729268
rect 546731 729263 546797 729266
rect 553033 729263 553099 729266
rect 556317 729193 556377 729553
rect 554689 729190 554755 729193
rect 556253 729190 556377 729193
rect 554689 729188 556377 729190
rect 554689 729132 554694 729188
rect 554750 729132 556258 729188
rect 556314 729132 556377 729188
rect 554689 729130 556377 729132
rect 554689 729127 554755 729130
rect 556253 729127 556319 729130
rect 501421 729052 502082 729054
rect 501421 728996 501426 729052
rect 501482 728996 502082 729052
rect 501421 728994 502082 728996
rect 529205 729052 529314 729057
rect 529205 728996 529210 729052
rect 529266 728996 529314 729052
rect 529205 728994 529314 728996
rect 501421 728991 501487 728994
rect 529205 728991 529271 728994
rect 368021 728918 368087 728921
rect 365629 728916 368087 728918
rect 365629 728860 365634 728916
rect 365690 728860 368026 728916
rect 368082 728860 368087 728916
rect 365629 728858 368087 728860
rect 365629 728855 365695 728858
rect 368021 728855 368087 728858
rect 335042 718386 335230 724614
rect 339192 718386 339340 724614
rect 335042 717846 339340 718386
rect 282278 708246 282478 714662
rect 286936 708246 287058 714662
rect 282278 707726 287058 708246
rect 252694 706184 252700 706248
rect 252764 706246 252770 706248
rect 556451 706246 556511 729553
rect 576976 729329 577036 729553
rect 583516 729405 583582 729566
rect 583511 729341 583517 729405
rect 583581 729341 583587 729405
rect 576976 729324 577111 729329
rect 576976 729268 577050 729324
rect 577106 729268 577111 729324
rect 576976 729266 577111 729268
rect 577045 729263 577111 729266
rect 578425 729054 578491 729057
rect 583651 729054 583711 729553
rect 600943 729326 601009 729329
rect 603973 729326 604039 729566
rect 604764 729326 604830 729329
rect 600943 729324 604830 729326
rect 600943 729268 600948 729324
rect 601004 729268 604769 729324
rect 604825 729268 604830 729324
rect 600943 729266 604830 729268
rect 600943 729263 601009 729266
rect 604764 729263 604830 729266
rect 608160 729326 608226 729329
rect 610519 729326 610579 729553
rect 631179 729329 631239 729553
rect 637719 729329 637779 729553
rect 611453 729326 611519 729329
rect 608160 729324 611519 729326
rect 608160 729268 608165 729324
rect 608221 729268 611458 729324
rect 611514 729268 611519 729324
rect 608160 729266 611519 729268
rect 608160 729263 608226 729266
rect 611453 729263 611519 729266
rect 631179 729324 631299 729329
rect 631179 729268 631238 729324
rect 631294 729268 631299 729324
rect 631179 729265 631299 729268
rect 631233 729263 631299 729265
rect 631969 729326 632035 729329
rect 637673 729326 637779 729329
rect 631969 729324 637779 729326
rect 631969 729268 631974 729324
rect 632030 729268 637678 729324
rect 637734 729268 637779 729324
rect 631969 729266 637779 729268
rect 631969 729263 632035 729266
rect 637673 729263 637739 729266
rect 578425 729052 583711 729054
rect 578425 728996 578430 729052
rect 578486 728996 583711 729052
rect 578425 728994 583711 728996
rect 637213 729054 637279 729057
rect 637851 729054 637911 729553
rect 652455 729326 652521 729329
rect 654513 729326 654579 729329
rect 655343 729326 655409 729329
rect 658376 729326 658436 729553
rect 664919 729329 664979 729553
rect 659164 729326 659230 729329
rect 652455 729324 659230 729326
rect 652455 729268 652460 729324
rect 652516 729268 654518 729324
rect 654574 729268 655348 729324
rect 655404 729268 659169 729324
rect 659225 729268 659230 729324
rect 652455 729266 659230 729268
rect 652455 729263 652521 729266
rect 654513 729263 654579 729266
rect 655343 729263 655409 729266
rect 659164 729263 659230 729266
rect 662560 729326 662626 729329
rect 664813 729326 664979 729329
rect 662560 729324 664979 729326
rect 662560 729268 662565 729324
rect 662621 729268 664818 729324
rect 664874 729268 664979 729324
rect 662560 729266 664979 729268
rect 662560 729263 662626 729266
rect 664813 729263 664879 729266
rect 637213 729052 637911 729054
rect 637213 728996 637218 729052
rect 637274 728996 637911 729052
rect 637213 728994 637911 728996
rect 578425 728991 578491 728994
rect 637213 728991 637279 728994
rect 583577 728918 583643 728921
rect 583534 728916 583643 728918
rect 583534 728860 583582 728916
rect 583638 728860 583643 728916
rect 583534 728855 583643 728860
rect 583534 728784 583594 728855
rect 583526 728720 583532 728784
rect 583596 728720 583602 728784
rect 252764 706186 556511 706246
rect 252764 706184 252770 706186
rect 322573 700086 322639 700089
rect 379061 700086 379127 700089
rect 322573 700084 379127 700086
rect 322573 700028 322578 700084
rect 322634 700028 379066 700084
rect 379122 700028 379127 700084
rect 322573 700026 379127 700028
rect 322573 700023 322639 700026
rect 379061 700023 379127 700026
rect 314937 699950 315003 699953
rect 385133 699950 385199 699953
rect 314937 699948 385199 699950
rect 314937 699892 314942 699948
rect 314998 699892 385138 699948
rect 385194 699892 385199 699948
rect 314937 699890 385199 699892
rect 314937 699887 315003 699890
rect 385133 699887 385199 699890
rect 288533 699814 288599 699817
rect 381085 699814 381151 699817
rect 288533 699812 381151 699814
rect 288533 699756 288538 699812
rect 288594 699756 381090 699812
rect 381146 699756 381151 699812
rect 288533 699754 381151 699756
rect 288533 699751 288599 699754
rect 381085 699751 381151 699754
rect 290414 699208 290420 699272
rect 290484 699270 290490 699272
rect 298377 699270 298443 699273
rect 290484 699268 298443 699270
rect 290484 699212 298382 699268
rect 298438 699212 298443 699268
rect 290484 699210 298443 699212
rect 290484 699208 290490 699210
rect 298377 699207 298443 699210
rect 301689 699270 301755 699273
rect 306841 699270 306907 699273
rect 301689 699268 306907 699270
rect 301689 699212 301694 699268
rect 301750 699212 306846 699268
rect 306902 699212 306907 699268
rect 301689 699210 306907 699212
rect 301689 699207 301755 699210
rect 306841 699207 306907 699210
rect 250721 699134 250787 699137
rect 310797 699134 310863 699137
rect 250721 699132 310863 699134
rect 250721 699076 250726 699132
rect 250782 699076 310802 699132
rect 310858 699076 310863 699132
rect 250721 699074 310863 699076
rect 250721 699071 250787 699074
rect 310797 699071 310863 699074
rect 291477 698998 291543 699001
rect 321009 698998 321075 699001
rect 279474 698938 291034 698998
rect 252510 698800 252516 698864
rect 252580 698862 252586 698864
rect 279474 698862 279534 698938
rect 252580 698802 279534 698862
rect 286601 698862 286667 698865
rect 290005 698862 290071 698865
rect 286601 698860 290071 698862
rect 286601 698804 286606 698860
rect 286662 698804 290010 698860
rect 290066 698804 290071 698860
rect 286601 698802 290071 698804
rect 252580 698800 252586 698802
rect 286601 698799 286667 698802
rect 290005 698799 290071 698802
rect 289085 698726 289151 698729
rect 288950 698724 289151 698726
rect 288950 698668 289090 698724
rect 289146 698668 289151 698724
rect 288950 698666 289151 698668
rect 290974 698726 291034 698938
rect 291477 698996 321075 698998
rect 291477 698940 291482 698996
rect 291538 698940 321014 698996
rect 321070 698940 321075 698996
rect 291477 698938 321075 698940
rect 291477 698935 291543 698938
rect 321009 698935 321075 698938
rect 312085 698862 312151 698865
rect 311030 698860 312151 698862
rect 311030 698804 312090 698860
rect 312146 698804 312151 698860
rect 311030 698802 312151 698804
rect 311030 698726 311090 698802
rect 312085 698799 312151 698802
rect 313557 698860 313623 698865
rect 313557 698804 313562 698860
rect 313618 698804 313623 698860
rect 313557 698799 313623 698804
rect 319077 698862 319143 698865
rect 323677 698862 323743 698865
rect 319077 698860 323743 698862
rect 319077 698804 319082 698860
rect 319138 698804 323682 698860
rect 323738 698804 323743 698860
rect 319077 698802 323743 698804
rect 319077 698799 319143 698802
rect 323677 698799 323743 698802
rect 290974 698666 311090 698726
rect 313560 698726 313620 698799
rect 367101 698726 367167 698729
rect 313560 698724 367167 698726
rect 313560 698668 367106 698724
rect 367162 698668 367167 698724
rect 313560 698666 367167 698668
rect 288950 698054 289010 698666
rect 289085 698663 289151 698666
rect 367101 698663 367167 698666
rect 320598 696009 320658 696618
rect 320598 696004 320707 696009
rect 320598 695948 320646 696004
rect 320702 695948 320707 696004
rect 320598 695946 320707 695948
rect 320641 695943 320707 695946
rect 288257 695190 288323 695193
rect 288950 695190 289010 695802
rect 288257 695188 289010 695190
rect 288257 695132 288262 695188
rect 288318 695132 289010 695188
rect 288257 695130 289010 695132
rect 288257 695127 288323 695130
rect 320782 694241 320842 694714
rect 370781 694646 370847 694649
rect 371149 694646 371215 694649
rect 370781 694644 371215 694646
rect 370781 694588 370786 694644
rect 370842 694588 371154 694644
rect 371210 694588 371215 694644
rect 370781 694586 371215 694588
rect 370781 694583 370847 694586
rect 371149 694583 371215 694586
rect 375013 694646 375079 694649
rect 375197 694646 375263 694649
rect 375013 694644 375263 694646
rect 375013 694588 375018 694644
rect 375074 694588 375202 694644
rect 375258 694588 375263 694644
rect 375013 694586 375263 694588
rect 375013 694583 375079 694586
rect 375197 694583 375263 694586
rect 364566 694448 364572 694512
rect 364636 694510 364642 694512
rect 365077 694510 365143 694513
rect 364636 694508 365143 694510
rect 364636 694452 365082 694508
rect 365138 694452 365143 694508
rect 364636 694450 365143 694452
rect 364636 694448 364642 694450
rect 365077 694447 365143 694450
rect 382230 694448 382236 694512
rect 382300 694510 382306 694512
rect 383109 694510 383175 694513
rect 382300 694508 383175 694510
rect 382300 694452 383114 694508
rect 383170 694452 383175 694508
rect 382300 694450 383175 694452
rect 382300 694448 382306 694450
rect 383109 694447 383175 694450
rect 676129 694510 676195 694513
rect 676299 694510 676466 694527
rect 676129 694508 676466 694510
rect 676129 694452 676134 694508
rect 676190 694461 676466 694508
rect 676190 694452 676369 694461
rect 676129 694450 676369 694452
rect 676129 694447 676195 694450
rect 320782 694236 320891 694241
rect 320782 694180 320830 694236
rect 320886 694180 320891 694236
rect 320782 694178 320891 694180
rect 320825 694175 320891 694178
rect 288441 693286 288507 693289
rect 288950 693286 289010 693898
rect 356981 693558 357047 693561
rect 362918 693558 362978 694102
rect 356981 693556 362978 693558
rect 356981 693500 356986 693556
rect 357042 693500 362978 693556
rect 356981 693498 362978 693500
rect 356981 693495 357047 693498
rect 288441 693284 289010 693286
rect 288441 693228 288446 693284
rect 288502 693228 289010 693284
rect 288441 693226 289010 693228
rect 288441 693223 288507 693226
rect 226248 692383 226265 692698
rect 226757 692383 226784 692698
rect 226248 692358 226784 692383
rect 320782 691926 320842 692538
rect 320917 691926 320983 691929
rect 320782 691924 320983 691926
rect 320782 691868 320922 691924
rect 320978 691868 320983 691924
rect 320782 691866 320983 691868
rect 320917 691863 320983 691866
rect 208309 691790 208375 691793
rect 209321 691790 209387 691793
rect 208128 691788 209387 691790
rect 208128 691732 208314 691788
rect 208370 691732 209326 691788
rect 209382 691732 209387 691788
rect 208128 691730 209387 691732
rect 208128 691716 208188 691730
rect 208309 691727 208375 691730
rect 209321 691727 209387 691730
rect 207928 691656 208188 691716
rect 208217 691587 208283 691590
rect 207928 691585 208283 691587
rect 207928 691529 208222 691585
rect 208278 691529 208283 691585
rect 207928 691527 208283 691529
rect 208217 691524 208283 691527
rect 207903 691322 208118 691388
rect 208217 691171 208283 691174
rect 207928 691169 208283 691171
rect 207928 691113 208222 691169
rect 208278 691113 208283 691169
rect 207928 691111 208283 691113
rect 208217 691110 208283 691111
rect 209965 691110 210031 691113
rect 208217 691108 210031 691110
rect 208220 691052 209970 691108
rect 210026 691052 210031 691108
rect 208220 691050 210031 691052
rect 209965 691047 210031 691050
rect 288809 691110 288875 691113
rect 288950 691110 289010 691722
rect 320641 691382 320707 691385
rect 288809 691108 289010 691110
rect 288809 691052 288814 691108
rect 288870 691052 289010 691108
rect 288809 691050 289010 691052
rect 320598 691380 320707 691382
rect 320598 691324 320646 691380
rect 320702 691324 320707 691380
rect 320598 691319 320707 691324
rect 288809 691047 288875 691050
rect 320598 690710 320658 691319
rect 362918 690569 362978 691110
rect 288717 690566 288783 690569
rect 288717 690564 289010 690566
rect 288717 690508 288722 690564
rect 288778 690508 289010 690564
rect 288717 690506 289010 690508
rect 288717 690503 288783 690506
rect 288950 689894 289010 690506
rect 362869 690564 362978 690569
rect 362869 690508 362874 690564
rect 362930 690508 362978 690564
rect 362869 690506 362978 690508
rect 362869 690503 362935 690506
rect 390334 689209 390394 689750
rect 390285 689204 390394 689209
rect 390285 689148 390290 689204
rect 390346 689148 390394 689204
rect 390285 689146 390394 689148
rect 390285 689143 390351 689146
rect 320774 688396 320780 688460
rect 320844 688396 320850 688460
rect 279885 687438 279951 687441
rect 288950 687438 289010 687642
rect 362409 687574 362475 687577
rect 362918 687574 362978 688118
rect 675945 687982 676011 687985
rect 675945 687980 676453 687982
rect 675945 687924 675950 687980
rect 676006 687924 676453 687980
rect 675945 687922 676453 687924
rect 675945 687919 676011 687922
rect 676129 687846 676195 687849
rect 676129 687844 676453 687846
rect 676129 687788 676134 687844
rect 676190 687788 676453 687844
rect 676129 687786 676453 687788
rect 676129 687783 676195 687786
rect 362409 687572 362978 687574
rect 362409 687516 362414 687572
rect 362470 687516 362978 687572
rect 362409 687514 362978 687516
rect 362409 687511 362475 687514
rect 279885 687436 289010 687438
rect 279885 687380 279890 687436
rect 279946 687380 289010 687436
rect 279885 687378 289010 687380
rect 279885 687375 279951 687378
rect 390377 687166 390443 687169
rect 390334 687164 390443 687166
rect 390334 687108 390382 687164
rect 390438 687108 390443 687164
rect 390334 687103 390443 687108
rect 390334 686970 390394 687103
rect 320598 686353 320658 686512
rect 320598 686348 320707 686353
rect 320598 686292 320646 686348
rect 320702 686292 320707 686348
rect 320598 686290 320707 686292
rect 320641 686287 320707 686290
rect 288533 686214 288599 686217
rect 288533 686212 289010 686214
rect 288533 686156 288538 686212
rect 288594 686156 289010 686212
rect 288533 686154 289010 686156
rect 288533 686151 288599 686154
rect 288950 685814 289010 686154
rect 360661 684990 360727 684993
rect 362501 684990 362567 684993
rect 362918 684990 362978 685126
rect 360661 684988 362978 684990
rect 360661 684932 360666 684988
rect 360722 684932 362506 684988
rect 362562 684932 362978 684988
rect 360661 684930 362978 684932
rect 360661 684927 360727 684930
rect 362501 684927 362567 684930
rect 320598 684177 320658 684378
rect 320598 684174 320707 684177
rect 321101 684174 321167 684177
rect 320598 684172 321167 684174
rect 320598 684116 320646 684172
rect 320702 684116 321106 684172
rect 321162 684116 321167 684172
rect 320598 684114 321167 684116
rect 320641 684111 320707 684114
rect 321101 684111 321167 684114
rect 288533 682950 288599 682953
rect 288950 682950 289010 683562
rect 288533 682948 289010 682950
rect 288533 682892 288538 682948
rect 288594 682892 289010 682948
rect 288533 682890 289010 682892
rect 288533 682887 288599 682890
rect 288625 682406 288691 682409
rect 288625 682404 289010 682406
rect 288625 682348 288630 682404
rect 288686 682348 289010 682404
rect 288625 682346 289010 682348
rect 288625 682343 288691 682346
rect 288950 681734 289010 682346
rect 320782 681862 320842 682474
rect 359833 681998 359899 682001
rect 362918 681998 362978 682134
rect 359833 681996 362978 681998
rect 359833 681940 359838 681996
rect 359894 681940 362978 681996
rect 359833 681938 362978 681940
rect 359833 681935 359899 681938
rect 320958 681862 320964 681864
rect 320782 681802 320964 681862
rect 320958 681800 320964 681802
rect 321028 681800 321034 681864
rect 279977 681454 280043 681457
rect 288625 681454 288691 681457
rect 279977 681452 288691 681454
rect 279977 681396 279982 681452
rect 280038 681396 288630 681452
rect 288686 681396 288691 681452
rect 279977 681394 288691 681396
rect 279977 681391 280043 681394
rect 288625 681391 288691 681394
rect 321009 681046 321075 681049
rect 320782 681044 321075 681046
rect 320782 680988 321014 681044
rect 321070 680988 321075 681044
rect 320782 680986 321075 680988
rect 320782 680374 320842 680986
rect 321009 680983 321075 680986
rect 390334 680233 390394 680774
rect 390285 680228 390394 680233
rect 390285 680172 390290 680228
rect 390346 680172 390394 680228
rect 390285 680170 390394 680172
rect 390285 680167 390351 680170
rect 288165 679142 288231 679145
rect 288950 679142 289010 679482
rect 288165 679140 289010 679142
rect 288165 679084 288170 679140
rect 288226 679084 289010 679140
rect 288165 679082 289010 679084
rect 288165 679079 288231 679082
rect 362593 679006 362659 679009
rect 362918 679006 362978 679142
rect 362593 679004 362978 679006
rect 362593 678948 362598 679004
rect 362654 678948 362978 679004
rect 362593 678946 362978 678948
rect 362593 678943 362659 678946
rect 320782 677782 320842 678394
rect 321193 677782 321259 677785
rect 390653 677782 390719 677785
rect 320782 677780 321259 677782
rect 320782 677724 321198 677780
rect 321254 677724 321259 677780
rect 320782 677722 321259 677724
rect 390518 677780 390719 677782
rect 390518 677724 390658 677780
rect 390714 677724 390719 677780
rect 390518 677722 390719 677724
rect 321193 677719 321259 677722
rect 390653 677719 390719 677722
rect 288073 676966 288139 676969
rect 288950 676966 289010 677578
rect 288073 676964 289010 676966
rect 288073 676908 288078 676964
rect 288134 676908 289010 676964
rect 288073 676906 289010 676908
rect 320733 676966 320799 676969
rect 320733 676964 320842 676966
rect 320733 676908 320738 676964
rect 320794 676908 320842 676964
rect 288073 676903 288139 676906
rect 320733 676903 320842 676908
rect 208861 676422 208927 676425
rect 208542 676420 208927 676422
rect 208217 676387 208283 676390
rect 208542 676387 208866 676420
rect 207928 676385 208866 676387
rect 207928 676329 208222 676385
rect 208278 676364 208866 676385
rect 208922 676364 208927 676420
rect 208278 676362 208927 676364
rect 208278 676329 208602 676362
rect 208861 676359 208927 676362
rect 207928 676327 208602 676329
rect 208217 676324 208283 676327
rect 320782 676294 320842 676903
rect 208125 676219 208191 676222
rect 207928 676217 208191 676219
rect 207928 676161 208130 676217
rect 208186 676161 208191 676217
rect 207928 676159 208191 676161
rect 208125 676156 208191 676159
rect 362317 675606 362383 675609
rect 362918 675606 362978 676150
rect 362317 675604 362978 675606
rect 208125 675592 208191 675595
rect 207928 675590 208191 675592
rect 207928 675534 208130 675590
rect 208186 675534 208191 675590
rect 362317 675548 362322 675604
rect 362378 675548 362978 675604
rect 362317 675546 362978 675548
rect 362317 675543 362383 675546
rect 207928 675532 208191 675534
rect 208125 675529 208191 675532
rect 208217 675451 208283 675454
rect 207928 675449 208283 675451
rect 207928 675393 208222 675449
rect 208278 675393 208283 675449
rect 207928 675391 208283 675393
rect 208217 675388 208283 675391
rect 287981 674790 288047 674793
rect 288950 674790 289010 675402
rect 320774 675000 320780 675064
rect 320844 675062 320850 675064
rect 321142 675062 321148 675064
rect 320844 675002 321148 675062
rect 320844 675000 320850 675002
rect 321142 675000 321148 675002
rect 321212 675000 321218 675064
rect 287981 674788 289010 674790
rect 287981 674732 287986 674788
rect 288042 674732 289010 674788
rect 287981 674730 289010 674732
rect 287981 674727 288047 674730
rect 320782 673705 320842 674314
rect 390334 674249 390394 674790
rect 390285 674244 390394 674249
rect 390285 674188 390290 674244
rect 390346 674188 390394 674244
rect 390285 674186 390394 674188
rect 390285 674183 390351 674186
rect 320733 673700 320842 673705
rect 320733 673644 320738 673700
rect 320794 673644 320842 673700
rect 320733 673642 320842 673644
rect 320733 673639 320799 673642
rect 360753 673566 360819 673569
rect 362685 673566 362751 673569
rect 360753 673564 362978 673566
rect 360753 673508 360758 673564
rect 360814 673508 362690 673564
rect 362746 673508 362978 673564
rect 360753 673506 362978 673508
rect 360753 673503 360819 673506
rect 362685 673503 362751 673506
rect 287889 672886 287955 672889
rect 288950 672886 289010 673498
rect 362918 673370 362978 673506
rect 287889 672884 289010 672886
rect 287889 672828 287894 672884
rect 287950 672828 289010 672884
rect 287889 672826 289010 672828
rect 287889 672823 287955 672826
rect 208125 672243 208191 672246
rect 208309 672243 208375 672246
rect 207928 672241 208375 672243
rect 207928 672185 208130 672241
rect 208186 672185 208314 672241
rect 208370 672185 208375 672241
rect 207928 672183 208375 672185
rect 208125 672180 208191 672183
rect 208309 672180 208375 672183
rect 208125 672070 208191 672073
rect 207928 672068 208191 672070
rect 207928 672012 208130 672068
rect 208186 672012 208191 672068
rect 207928 672010 208191 672012
rect 208125 672007 208191 672010
rect 320782 671662 320842 672138
rect 321285 671662 321351 671665
rect 320782 671660 321351 671662
rect 320782 671604 321290 671660
rect 321346 671604 321351 671660
rect 320782 671602 321351 671604
rect 321285 671599 321351 671602
rect 390518 671529 390578 672070
rect 390469 671524 390578 671529
rect 390469 671468 390474 671524
rect 390530 671468 390578 671524
rect 390469 671466 390578 671468
rect 390469 671463 390535 671466
rect 286417 671118 286483 671121
rect 288950 671118 289010 671322
rect 286417 671116 289010 671118
rect 286417 671060 286422 671116
rect 286478 671060 289010 671116
rect 286417 671058 289010 671060
rect 286417 671055 286483 671058
rect 323967 670342 341848 670358
rect 323967 670324 341500 670342
rect 208125 669731 208191 669734
rect 207928 669729 208191 669731
rect 207928 669673 208130 669729
rect 208186 669673 208191 669729
rect 207928 669671 208191 669673
rect 208125 669668 208191 669671
rect 320782 669622 320842 670234
rect 323967 669868 324036 670324
rect 326786 669868 341500 670324
rect 323967 669822 341500 669868
rect 341796 669822 341848 670342
rect 323967 669804 341848 669822
rect 343118 670294 362101 670318
rect 343118 669782 343162 670294
rect 343450 670284 362101 670294
rect 343450 669812 359258 670284
rect 362026 669812 362101 670284
rect 343450 669782 362101 669812
rect 343118 669764 362101 669782
rect 321009 669622 321075 669625
rect 320782 669620 321075 669622
rect 320782 669564 321014 669620
rect 321070 669564 321075 669620
rect 320782 669562 321075 669564
rect 321009 669559 321075 669562
rect 288950 668806 289010 669418
rect 390334 668945 390394 669078
rect 390334 668940 390443 668945
rect 390334 668884 390382 668940
rect 390438 668884 390443 668940
rect 390334 668882 390443 668884
rect 390377 668879 390443 668882
rect 289085 668806 289151 668809
rect 288950 668804 289151 668806
rect 288950 668748 289090 668804
rect 289146 668748 289151 668804
rect 288950 668746 289151 668748
rect 289085 668743 289151 668746
rect 208309 668096 208375 668099
rect 207928 668094 208375 668096
rect 207928 668038 208314 668094
rect 208370 668038 208375 668094
rect 207928 668036 208375 668038
rect 208309 668033 208375 668036
rect 208309 667926 208375 667929
rect 207928 667924 208375 667926
rect 207928 667868 208314 667924
rect 208370 667868 208375 667924
rect 207928 667866 208375 667868
rect 208309 667863 208375 667866
rect 220034 667728 222160 667758
rect 220034 667552 220076 667728
rect 222120 667552 222160 667728
rect 220034 667516 222160 667552
rect 320782 667446 320842 668058
rect 325241 667446 325307 667449
rect 320782 667444 325307 667446
rect 320782 667388 325246 667444
rect 325302 667388 325307 667444
rect 320782 667386 325307 667388
rect 325241 667383 325307 667386
rect 290414 667248 290420 667312
rect 290484 667310 290490 667312
rect 290833 667310 290899 667313
rect 290484 667308 290899 667310
rect 290484 667252 290838 667308
rect 290894 667252 290899 667308
rect 290484 667250 290899 667252
rect 290484 667248 290490 667250
rect 290833 667247 290899 667250
rect 311349 667310 311415 667313
rect 311533 667310 311599 667313
rect 390193 667310 390259 667313
rect 311349 667308 325902 667310
rect 311349 667252 311354 667308
rect 311410 667252 311538 667308
rect 311594 667252 325902 667308
rect 311349 667250 325902 667252
rect 311349 667247 311415 667250
rect 311533 667247 311599 667250
rect 301597 667174 301663 667177
rect 308221 667174 308287 667177
rect 308589 667174 308655 667177
rect 301597 667172 302718 667174
rect 236436 667020 243140 667120
rect 301597 667116 301602 667172
rect 301658 667116 302718 667172
rect 301597 667114 302718 667116
rect 301597 667111 301663 667114
rect 236436 665954 236536 667020
rect 242984 665954 243140 667020
rect 302658 667038 302718 667114
rect 308221 667172 308655 667174
rect 308221 667116 308226 667172
rect 308282 667116 308594 667172
rect 308650 667116 308655 667172
rect 308221 667114 308655 667116
rect 308221 667111 308287 667114
rect 308589 667111 308655 667114
rect 320590 667112 320596 667176
rect 320660 667174 320666 667176
rect 320958 667174 320964 667176
rect 320660 667114 320964 667174
rect 320660 667112 320666 667114
rect 320958 667112 320964 667114
rect 321028 667112 321034 667176
rect 325842 667174 325902 667250
rect 356754 667308 390259 667310
rect 356754 667252 390198 667308
rect 390254 667252 390259 667308
rect 356754 667250 390259 667252
rect 356754 667174 356814 667250
rect 390193 667247 390259 667250
rect 325842 667114 356814 667174
rect 381085 667174 381151 667177
rect 381269 667174 381335 667177
rect 381085 667172 381335 667174
rect 381085 667116 381090 667172
rect 381146 667116 381274 667172
rect 381330 667116 381335 667172
rect 381085 667114 381335 667116
rect 381085 667111 381151 667114
rect 381269 667111 381335 667114
rect 361121 667038 361187 667041
rect 302658 667036 361187 667038
rect 302658 666980 361126 667036
rect 361182 666980 361187 667036
rect 302658 666978 361187 666980
rect 361121 666975 361187 666978
rect 361305 667038 361371 667041
rect 364566 667038 364572 667040
rect 361305 667036 364572 667038
rect 361305 666980 361310 667036
rect 361366 666980 364572 667036
rect 361305 666978 364572 666980
rect 361305 666975 361371 666978
rect 364566 666976 364572 666978
rect 364636 666976 364642 667040
rect 307117 666902 307183 666905
rect 390377 666902 390443 666905
rect 307117 666900 390443 666902
rect 307117 666844 307122 666900
rect 307178 666844 390382 666900
rect 390438 666844 390443 666900
rect 307117 666842 390443 666844
rect 307117 666839 307183 666842
rect 390377 666839 390443 666842
rect 289361 666766 289427 666769
rect 382230 666766 382236 666768
rect 289361 666764 382236 666766
rect 289361 666708 289366 666764
rect 289422 666708 382236 666764
rect 289361 666706 382236 666708
rect 289361 666703 289427 666706
rect 382230 666704 382236 666706
rect 382300 666704 382306 666768
rect 325241 666630 325307 666633
rect 325241 666628 372270 666630
rect 325241 666572 325246 666628
rect 325302 666572 372270 666628
rect 325241 666570 372270 666572
rect 325241 666567 325307 666570
rect 372210 666494 372270 666570
rect 385317 666494 385383 666497
rect 372210 666492 385383 666494
rect 372210 666436 385322 666492
rect 385378 666436 385383 666492
rect 372210 666434 385383 666436
rect 385317 666431 385383 666434
rect 251774 666024 251780 666088
rect 251844 666086 251850 666088
rect 676129 666086 676195 666089
rect 251844 666084 676195 666086
rect 251844 666028 676134 666084
rect 676190 666028 676195 666084
rect 251844 666026 676195 666028
rect 251844 666024 251850 666026
rect 676129 666023 676195 666026
rect 236436 665890 243140 665954
rect 208217 665389 208283 665392
rect 207928 665387 208283 665389
rect 207928 665331 208222 665387
rect 208278 665331 208283 665387
rect 207928 665329 208283 665331
rect 208217 665326 208283 665329
rect 364566 664936 364572 665000
rect 364636 664998 364642 665000
rect 365261 664998 365327 665001
rect 364636 664996 365327 664998
rect 364636 664940 365266 664996
rect 365322 664940 365327 664996
rect 364636 664938 365327 664940
rect 364636 664936 364642 664938
rect 365261 664935 365327 664938
rect 208125 663951 208191 663954
rect 207928 663949 208191 663951
rect 207928 663893 208130 663949
rect 208186 663893 208191 663949
rect 207928 663891 208191 663893
rect 207990 663781 208050 663891
rect 208125 663888 208191 663891
rect 207928 663721 208050 663781
rect 207990 663611 208050 663721
rect 207928 663551 208050 663611
rect 208125 660895 208191 660898
rect 207928 660893 208191 660895
rect 207928 660837 208130 660893
rect 208186 660837 208191 660893
rect 207928 660835 208191 660837
rect 208125 660832 208191 660835
rect 208125 659804 208191 659807
rect 207928 659802 208191 659804
rect 207928 659746 208130 659802
rect 208186 659746 208191 659802
rect 207928 659744 208191 659746
rect 208125 659741 208191 659744
rect 207928 659573 208188 659633
rect 208128 659422 208188 659573
rect 210057 659422 210123 659425
rect 208128 659420 210123 659422
rect 208128 659371 210062 659420
rect 207928 659364 210062 659371
rect 210118 659364 210123 659420
rect 207928 659362 210123 659364
rect 207928 659311 208188 659362
rect 210057 659359 210123 659362
rect 209752 658662 216288 658690
rect 209752 658661 215274 658662
rect 209752 658153 209784 658661
rect 210076 658184 215274 658661
rect 216250 658184 216288 658662
rect 210076 658153 216288 658184
rect 209752 658128 216288 658153
rect 210342 657478 211698 657548
rect 210342 657472 210476 657478
rect 209752 656894 210476 657472
rect 208125 656034 208191 656037
rect 209763 656034 209937 656894
rect 210342 656586 210476 656894
rect 211618 656586 211698 657478
rect 210342 656482 211698 656586
rect 207928 656032 209937 656034
rect 207928 655976 208130 656032
rect 208186 656020 209937 656032
rect 208186 655976 209142 656020
rect 207928 655974 209142 655976
rect 208125 655971 209142 655974
rect 208128 655964 209142 655971
rect 209198 655964 209937 656020
rect 208128 655962 209937 655964
rect 209119 655863 209937 655962
rect 209763 655861 209937 655863
rect 210149 655206 210215 655209
rect 208128 655204 210215 655206
rect 208128 655148 210154 655204
rect 210210 655148 210215 655204
rect 208128 655146 210215 655148
rect 208128 654994 208188 655146
rect 210149 655143 210215 655146
rect 208125 654991 208191 654994
rect 207928 654989 208191 654991
rect 207928 654933 208130 654989
rect 208186 654933 208191 654989
rect 207928 654931 208191 654933
rect 208125 654928 208191 654931
rect 213461 654662 213527 654665
rect 208542 654660 213527 654662
rect 208542 654640 213466 654660
rect 207928 654604 213466 654640
rect 213522 654604 213527 654660
rect 207928 654602 213527 654604
rect 207928 654580 208602 654602
rect 213461 654599 213527 654602
rect 207928 654429 208188 654489
rect 208128 654390 208188 654429
rect 208861 654390 208927 654393
rect 208128 654388 208927 654390
rect 208128 654332 208866 654388
rect 208922 654332 208927 654388
rect 208128 654330 208927 654332
rect 208861 654327 208927 654330
rect 675577 653846 675643 653849
rect 676129 653846 676195 653849
rect 675577 653844 676318 653846
rect 675577 653788 675582 653844
rect 675638 653788 676134 653844
rect 676190 653788 676318 653844
rect 675577 653786 676318 653788
rect 675577 653783 675643 653786
rect 676129 653783 676195 653786
rect 676258 653727 676318 653786
rect 676258 653661 676466 653727
rect 208125 652318 208191 652321
rect 207928 652316 208191 652318
rect 207928 652260 208130 652316
rect 208186 652260 208191 652316
rect 207928 652258 208191 652260
rect 208125 652255 208191 652258
rect 208125 652185 208191 652188
rect 207928 652183 208191 652185
rect 207928 652127 208130 652183
rect 208186 652127 208191 652183
rect 207928 652125 208191 652127
rect 208125 652122 208191 652125
rect 207934 651922 208122 651988
rect 614397 651942 614463 651945
rect 619406 651942 619412 651944
rect 614397 651940 619412 651942
rect 614397 651884 614402 651940
rect 614458 651884 619412 651940
rect 614397 651882 619412 651884
rect 614397 651879 614463 651882
rect 619406 651880 619412 651882
rect 619476 651880 619482 651944
rect 616789 651806 616855 651809
rect 619038 651806 619044 651808
rect 616789 651804 619044 651806
rect 616789 651748 616794 651804
rect 616850 651748 619044 651804
rect 616789 651746 619044 651748
rect 616789 651743 616855 651746
rect 619038 651744 619044 651746
rect 619108 651744 619114 651808
rect 208125 651721 208191 651724
rect 207928 651719 208318 651721
rect 207928 651663 208130 651719
rect 208186 651670 208318 651719
rect 208953 651670 209019 651673
rect 208186 651668 209019 651670
rect 208186 651663 208958 651668
rect 207928 651661 208958 651663
rect 208125 651658 208958 651661
rect 208174 651612 208958 651658
rect 209014 651612 209019 651668
rect 208174 651610 209019 651612
rect 208953 651607 209019 651610
rect 612373 651670 612439 651673
rect 620694 651670 620700 651672
rect 612373 651668 620700 651670
rect 612373 651612 612378 651668
rect 612434 651612 620700 651668
rect 612373 651610 620700 651612
rect 612373 651607 612439 651610
rect 620694 651608 620700 651610
rect 620764 651608 620770 651672
rect 612189 651534 612255 651537
rect 619222 651534 619228 651536
rect 612189 651532 619228 651534
rect 612189 651476 612194 651532
rect 612250 651476 619228 651532
rect 612189 651474 619228 651476
rect 612189 651471 612255 651474
rect 619222 651472 619228 651474
rect 619292 651472 619298 651536
rect 612281 650854 612347 650857
rect 619590 650854 619596 650856
rect 612281 650852 619596 650854
rect 612281 650796 612286 650852
rect 612342 650796 619596 650852
rect 612281 650794 619596 650796
rect 612281 650791 612347 650794
rect 619590 650792 619596 650794
rect 619660 650792 619666 650856
rect 320590 650520 320596 650584
rect 320660 650582 320666 650584
rect 639513 650582 639579 650585
rect 320660 650580 639579 650582
rect 320660 650524 639518 650580
rect 639574 650524 639579 650580
rect 320660 650522 639579 650524
rect 320660 650520 320666 650522
rect 639513 650519 639579 650522
rect 252326 648480 252332 648544
rect 252396 648542 252402 648544
rect 311533 648542 311599 648545
rect 252396 648540 311599 648542
rect 252396 648484 311538 648540
rect 311594 648484 311599 648540
rect 252396 648482 311599 648484
rect 252396 648480 252402 648482
rect 311533 648479 311599 648482
rect 250445 648406 250511 648409
rect 320774 648406 320780 648408
rect 250445 648404 320780 648406
rect 250445 648348 250450 648404
rect 250506 648348 320780 648404
rect 250445 648346 320780 648348
rect 250445 648343 250511 648346
rect 320774 648344 320780 648346
rect 320844 648344 320850 648408
rect 252142 647392 252148 647456
rect 252212 647454 252218 647456
rect 666745 647454 666811 647457
rect 252212 647452 666811 647454
rect 252212 647396 666750 647452
rect 666806 647396 666811 647452
rect 252212 647394 666811 647396
rect 252212 647392 252218 647394
rect 666745 647391 666811 647394
rect 417333 647318 417399 647321
rect 627737 647318 627803 647321
rect 417333 647316 627803 647318
rect 417333 647260 417338 647316
rect 417394 647260 627742 647316
rect 627798 647260 627803 647316
rect 417333 647258 627803 647260
rect 417333 647255 417399 647258
rect 627737 647255 627803 647258
rect 208166 647120 208172 647184
rect 208236 647182 208242 647184
rect 446221 647182 446287 647185
rect 208236 647180 446287 647182
rect 208236 647124 446226 647180
rect 446282 647124 446287 647180
rect 208236 647122 446287 647124
rect 208236 647120 208242 647122
rect 446221 647119 446287 647122
rect 676129 647182 676195 647185
rect 676129 647180 676453 647182
rect 676129 647124 676134 647180
rect 676190 647124 676453 647180
rect 676129 647122 676453 647124
rect 676129 647119 676195 647122
rect 251958 646984 251964 647048
rect 252028 647046 252034 647048
rect 676037 647046 676103 647049
rect 252028 647044 676103 647046
rect 252028 646988 676042 647044
rect 676098 646988 676103 647044
rect 252028 646986 676103 646988
rect 252028 646984 252034 646986
rect 676037 646983 676103 646986
rect 676224 646986 676453 647046
rect 254401 646910 254467 646913
rect 257897 646910 257963 646913
rect 254401 646908 257963 646910
rect 254401 646852 254406 646908
rect 254462 646852 257902 646908
rect 257958 646852 257963 646908
rect 254401 646850 257963 646852
rect 254401 646847 254467 646850
rect 257897 646847 257963 646850
rect 258541 646910 258607 646913
rect 259185 646910 259251 646913
rect 258541 646908 259251 646910
rect 258541 646852 258546 646908
rect 258602 646852 259190 646908
rect 259246 646852 259251 646908
rect 258541 646850 259251 646852
rect 258541 646847 258607 646850
rect 259185 646847 259251 646850
rect 278505 646910 278571 646913
rect 279977 646910 280043 646913
rect 278505 646908 280043 646910
rect 278505 646852 278510 646908
rect 278566 646852 279982 646908
rect 280038 646852 280043 646908
rect 278505 646850 280043 646852
rect 278505 646847 278571 646850
rect 279977 646847 280043 646850
rect 287245 646910 287311 646913
rect 288073 646910 288139 646913
rect 287245 646908 288139 646910
rect 287245 646852 287250 646908
rect 287306 646852 288078 646908
rect 288134 646852 288139 646908
rect 287245 646850 288139 646852
rect 287245 646847 287311 646850
rect 288073 646847 288139 646850
rect 301597 646910 301663 646913
rect 302425 646910 302491 646913
rect 301597 646908 302491 646910
rect 301597 646852 301602 646908
rect 301658 646852 302430 646908
rect 302486 646852 302491 646908
rect 301597 646850 302491 646852
rect 301597 646847 301663 646850
rect 302425 646847 302491 646850
rect 315949 646910 316015 646913
rect 316777 646910 316843 646913
rect 315949 646908 316843 646910
rect 315949 646852 315954 646908
rect 316010 646852 316782 646908
rect 316838 646852 316843 646908
rect 315949 646850 316843 646852
rect 315949 646847 316015 646850
rect 316777 646847 316843 646850
rect 344653 646910 344719 646913
rect 345481 646910 345547 646913
rect 344653 646908 345547 646910
rect 344653 646852 344658 646908
rect 344714 646852 345486 646908
rect 345542 646852 345547 646908
rect 344653 646850 345547 646852
rect 344653 646847 344719 646850
rect 345481 646847 345547 646850
rect 402061 646910 402127 646913
rect 403073 646910 403139 646913
rect 402061 646908 403139 646910
rect 402061 646852 402066 646908
rect 402122 646852 403078 646908
rect 403134 646852 403139 646908
rect 402061 646850 403139 646852
rect 402061 646847 402127 646850
rect 403073 646847 403139 646850
rect 474281 646910 474347 646913
rect 475017 646910 475083 646913
rect 474281 646908 475083 646910
rect 474281 646852 474286 646908
rect 474342 646852 475022 646908
rect 475078 646852 475083 646908
rect 474281 646850 475083 646852
rect 474281 646847 474347 646850
rect 475017 646847 475083 646850
rect 512461 646910 512527 646913
rect 513289 646910 513355 646913
rect 512461 646908 513355 646910
rect 512461 646852 512466 646908
rect 512522 646852 513294 646908
rect 513350 646852 513355 646908
rect 512461 646850 513355 646852
rect 512461 646847 512527 646850
rect 513289 646847 513355 646850
rect 536749 646910 536815 646913
rect 537393 646910 537459 646913
rect 536749 646908 537459 646910
rect 536749 646852 536754 646908
rect 536810 646852 537398 646908
rect 537454 646852 537459 646908
rect 536749 646850 537459 646852
rect 536749 646847 536815 646850
rect 537393 646847 537459 646850
rect 541165 646910 541231 646913
rect 542177 646910 542243 646913
rect 541165 646908 542243 646910
rect 541165 646852 541170 646908
rect 541226 646852 542182 646908
rect 542238 646852 542243 646908
rect 541165 646850 542243 646852
rect 541165 646847 541231 646850
rect 542177 646847 542243 646850
rect 569869 646910 569935 646913
rect 570881 646910 570947 646913
rect 569869 646908 570947 646910
rect 569869 646852 569874 646908
rect 569930 646852 570886 646908
rect 570942 646852 570947 646908
rect 569869 646850 570947 646852
rect 569869 646847 569935 646850
rect 570881 646847 570947 646850
rect 584221 646910 584287 646913
rect 585233 646910 585299 646913
rect 584221 646908 585299 646910
rect 584221 646852 584226 646908
rect 584282 646852 585238 646908
rect 585294 646852 585299 646908
rect 584221 646850 585299 646852
rect 584221 646847 584287 646850
rect 585233 646847 585299 646850
rect 598573 646910 598639 646913
rect 599585 646910 599651 646913
rect 598573 646908 599651 646910
rect 598573 646852 598578 646908
rect 598634 646852 599590 646908
rect 599646 646852 599651 646908
rect 598573 646850 599651 646852
rect 598573 646847 598639 646850
rect 599585 646847 599651 646850
rect 612925 646910 612991 646913
rect 613937 646910 614003 646913
rect 612925 646908 614003 646910
rect 612925 646852 612930 646908
rect 612986 646852 613942 646908
rect 613998 646852 614003 646908
rect 612925 646850 614003 646852
rect 612925 646847 612991 646850
rect 613937 646847 614003 646850
rect 617893 646910 617959 646913
rect 618721 646910 618787 646913
rect 617893 646908 618787 646910
rect 617893 646852 617898 646908
rect 617954 646852 618726 646908
rect 618782 646852 618787 646908
rect 617893 646850 618787 646852
rect 617893 646847 617959 646850
rect 618721 646847 618787 646850
rect 675209 646910 675275 646913
rect 676224 646910 676284 646986
rect 675209 646908 676284 646910
rect 675209 646852 675214 646908
rect 675270 646852 676284 646908
rect 675209 646850 676284 646852
rect 675209 646847 675275 646850
rect 619406 644672 619412 644736
rect 619476 644672 619482 644736
rect 619414 644462 619474 644672
rect 619774 644462 619780 644464
rect 619414 644402 619780 644462
rect 619774 644400 619780 644402
rect 619844 644400 619850 644464
rect 252561 642286 252627 642289
rect 252334 642284 252627 642286
rect 252334 642228 252566 642284
rect 252622 642228 252627 642284
rect 252334 642226 252627 642228
rect 252334 642014 252394 642226
rect 252561 642223 252627 642226
rect 252334 641954 252578 642014
rect 208217 639022 208283 639025
rect 207946 639020 208283 639022
rect 207946 638964 208222 639020
rect 208278 638964 208283 639020
rect 207946 638962 208283 638964
rect 208217 638959 208283 638962
rect 208401 638886 208467 638889
rect 207946 638884 208467 638886
rect 207946 638828 208406 638884
rect 208462 638828 208467 638884
rect 207946 638826 208467 638828
rect 208401 638823 208467 638826
rect 619222 637464 619228 637528
rect 619292 637464 619298 637528
rect 619230 636710 619290 637464
rect 620009 636710 620075 636713
rect 619230 636708 620075 636710
rect 619230 636652 620014 636708
rect 620070 636652 620075 636708
rect 619230 636650 620075 636652
rect 620009 636647 620075 636650
rect 619038 632432 619044 632496
rect 619108 632432 619114 632496
rect 207934 632273 208126 632339
rect 208066 632222 208126 632273
rect 208953 632222 209019 632225
rect 208066 632220 209019 632222
rect 208066 632164 208958 632220
rect 209014 632164 209019 632220
rect 208066 632162 209019 632164
rect 208953 632159 209019 632162
rect 619038 632160 619044 632224
rect 619108 632222 619114 632224
rect 621481 632222 621547 632225
rect 619108 632220 621547 632222
rect 619108 632164 621486 632220
rect 621542 632164 621547 632220
rect 619108 632162 621547 632164
rect 619108 632160 619114 632162
rect 621481 632159 621547 632162
rect 619038 632024 619044 632088
rect 619108 632086 619114 632088
rect 620009 632086 620075 632089
rect 619108 632084 620075 632086
rect 619108 632028 620014 632084
rect 620070 632028 620075 632084
rect 619108 632026 620075 632028
rect 619108 632024 619114 632026
rect 620009 632023 620075 632026
rect 619038 628624 619044 628688
rect 619108 628686 619114 628688
rect 619108 628626 619290 628686
rect 619108 628624 619114 628626
rect 619230 628416 619290 628626
rect 619222 628352 619228 628416
rect 619292 628352 619298 628416
rect 208033 628278 208099 628281
rect 208166 628278 208172 628280
rect 208033 628276 208172 628278
rect 208033 628220 208038 628276
rect 208094 628220 208172 628276
rect 208033 628218 208172 628220
rect 208033 628215 208099 628218
rect 208166 628216 208172 628218
rect 208236 628216 208242 628280
rect 251825 627870 251891 627873
rect 251825 627868 252578 627870
rect 251825 627812 251830 627868
rect 251886 627812 252578 627868
rect 251825 627810 252578 627812
rect 251825 627807 251891 627810
rect 208033 625705 208099 625710
rect 208033 625649 208038 625705
rect 208094 625694 208099 625705
rect 208217 625694 208283 625697
rect 208585 625694 208651 625697
rect 208094 625692 208651 625694
rect 208094 625649 208222 625692
rect 208033 625644 208222 625649
rect 208036 625636 208222 625644
rect 208278 625636 208590 625692
rect 208646 625636 208651 625692
rect 208036 625634 208651 625636
rect 208217 625631 208283 625634
rect 208585 625631 208651 625634
rect 619089 624472 619155 624473
rect 619084 624408 619090 624472
rect 619154 624470 619160 624472
rect 619154 624410 619246 624470
rect 619154 624408 619160 624410
rect 619089 624407 619155 624408
rect 208033 623828 208099 623831
rect 208033 623826 208234 623828
rect 208033 623770 208038 623826
rect 208094 623790 208234 623826
rect 208953 623790 209019 623793
rect 211529 623790 211595 623793
rect 208094 623788 211595 623790
rect 208094 623770 208958 623788
rect 208033 623768 208958 623770
rect 208033 623765 208099 623768
rect 208174 623732 208958 623768
rect 209014 623732 211534 623788
rect 211590 623732 211595 623788
rect 208174 623730 211595 623732
rect 208953 623727 209019 623730
rect 211529 623727 211595 623730
rect 619089 621342 619155 621345
rect 619089 621340 619658 621342
rect 619089 621284 619094 621340
rect 619150 621284 619658 621340
rect 619089 621282 619658 621284
rect 619089 621279 619155 621282
rect 619598 621208 619658 621282
rect 619406 621206 619412 621208
rect 619230 621146 619412 621206
rect 619230 620936 619290 621146
rect 619406 621144 619412 621146
rect 619476 621144 619482 621208
rect 619590 621144 619596 621208
rect 619660 621144 619666 621208
rect 619222 620872 619228 620936
rect 619292 620872 619298 620936
rect 252377 620798 252443 620801
rect 252377 620796 252578 620798
rect 252377 620740 252382 620796
rect 252438 620740 252578 620796
rect 252377 620738 252578 620740
rect 252377 620735 252443 620738
rect 619590 618350 619596 618352
rect 619230 618290 619596 618350
rect 619590 618288 619596 618290
rect 619660 618288 619666 618352
rect 247409 613726 247475 613729
rect 247409 613724 252578 613726
rect 247409 613668 247414 613724
rect 247470 613668 252578 613724
rect 247409 613666 252578 613668
rect 247409 613663 247475 613666
rect 208166 612984 208172 613048
rect 208236 613046 208242 613048
rect 209321 613046 209387 613049
rect 208236 613044 209387 613046
rect 208236 612988 209326 613044
rect 209382 612988 209387 613044
rect 208236 612986 209387 612988
rect 208236 612984 208242 612986
rect 209321 612983 209387 612986
rect 675301 613046 675367 613049
rect 675301 613044 676353 613046
rect 675301 612988 675306 613044
rect 675362 612988 676353 613044
rect 675301 612986 676353 612988
rect 675301 612983 675367 612986
rect 676293 612927 676353 612986
rect 676293 612861 676466 612927
rect 619089 611822 619155 611825
rect 619089 611820 619474 611822
rect 619089 611764 619094 611820
rect 619150 611764 619474 611820
rect 619089 611762 619474 611764
rect 619089 611759 619155 611762
rect 619089 611686 619155 611689
rect 619222 611686 619228 611688
rect 619089 611684 619228 611686
rect 208073 611654 208504 611655
rect 208073 611649 208559 611654
rect 208073 611611 208498 611649
rect 207946 611595 208498 611611
rect 207946 611551 208133 611595
rect 208480 611593 208498 611595
rect 208554 611593 208559 611649
rect 619089 611628 619094 611684
rect 619150 611628 619228 611684
rect 619089 611626 619228 611628
rect 619089 611623 619155 611626
rect 619222 611624 619228 611626
rect 619292 611624 619298 611688
rect 208480 611591 208559 611593
rect 208493 611588 208559 611591
rect 619414 611550 619474 611762
rect 208309 611529 208375 611532
rect 208193 611527 208375 611529
rect 208193 611479 208314 611527
rect 207946 611471 208314 611479
rect 208370 611471 208375 611527
rect 207946 611466 208375 611471
rect 619230 611490 619474 611550
rect 207946 611419 208253 611466
rect 619230 611218 619290 611490
rect 619089 610734 619155 610737
rect 619222 610734 619228 610736
rect 619089 610732 619228 610734
rect 619089 610676 619094 610732
rect 619150 610676 619228 610732
rect 619089 610674 619228 610676
rect 619089 610671 619155 610674
rect 619222 610672 619228 610674
rect 619292 610672 619298 610736
rect 208534 609176 208540 609240
rect 208604 609238 208610 609240
rect 208677 609238 208743 609241
rect 208604 609236 208743 609238
rect 208604 609180 208682 609236
rect 208738 609180 208743 609236
rect 208604 609178 208743 609180
rect 208604 609176 208610 609178
rect 208677 609175 208743 609178
rect 252009 606654 252075 606657
rect 252377 606654 252443 606657
rect 252009 606652 252578 606654
rect 252009 606596 252014 606652
rect 252070 606596 252382 606652
rect 252438 606596 252578 606652
rect 252009 606594 252578 606596
rect 252009 606591 252075 606594
rect 252377 606591 252443 606594
rect 675577 606382 675643 606385
rect 675577 606380 676453 606382
rect 675577 606324 675582 606380
rect 675638 606324 676453 606380
rect 675577 606322 676453 606324
rect 675577 606319 675643 606322
rect 208166 606184 208172 606248
rect 208236 606246 208242 606248
rect 208718 606246 208724 606248
rect 208236 606186 208724 606246
rect 208236 606184 208242 606186
rect 208718 606184 208724 606186
rect 208788 606184 208794 606248
rect 669689 606246 669755 606249
rect 669689 606244 676453 606246
rect 669689 606188 669694 606244
rect 669750 606188 676453 606244
rect 669689 606186 676453 606188
rect 669689 606183 669755 606186
rect 208033 605725 208099 605730
rect 208033 605669 208038 605725
rect 208094 605669 208099 605725
rect 208033 605664 208099 605669
rect 208036 605566 208096 605664
rect 208166 605566 208172 605568
rect 208036 605506 208172 605566
rect 208166 605504 208172 605506
rect 208236 605504 208242 605568
rect 619222 605368 619228 605432
rect 619292 605430 619298 605432
rect 619365 605430 619431 605433
rect 619292 605428 619431 605430
rect 619292 605372 619370 605428
rect 619426 605372 619431 605428
rect 619292 605370 619431 605372
rect 619292 605368 619298 605370
rect 619365 605367 619431 605370
rect 207934 604886 208138 604939
rect 208217 604886 208283 604889
rect 207934 604884 208283 604886
rect 207934 604873 208222 604884
rect 208071 604828 208222 604873
rect 208278 604828 208283 604884
rect 208071 604826 208283 604828
rect 208217 604823 208283 604826
rect 208219 604734 208283 604823
rect 208219 604729 208285 604734
rect 208219 604673 208224 604729
rect 208280 604673 208285 604729
rect 208219 604666 208285 604673
rect 619457 604206 619523 604209
rect 619230 604204 619523 604206
rect 619230 604148 619462 604204
rect 619518 604148 619523 604204
rect 619230 604146 619523 604148
rect 619457 604143 619523 604146
rect 619222 603872 619228 603936
rect 619292 603934 619298 603936
rect 619365 603934 619431 603937
rect 619292 603932 619431 603934
rect 619292 603876 619370 603932
rect 619426 603876 619431 603932
rect 619292 603874 619431 603876
rect 619292 603872 619298 603874
rect 619365 603871 619431 603874
rect 208033 603432 208099 603437
rect 208033 603376 208038 603432
rect 208094 603390 208099 603432
rect 208534 603390 208540 603392
rect 208094 603376 208540 603390
rect 208033 603371 208540 603376
rect 208036 603330 208540 603371
rect 208534 603328 208540 603330
rect 208604 603328 208610 603392
rect 208493 602166 208559 602169
rect 208036 602164 208559 602166
rect 208036 602122 208498 602164
rect 208033 602117 208498 602122
rect 208033 602061 208038 602117
rect 208094 602108 208498 602117
rect 208554 602108 208559 602164
rect 208094 602106 208559 602108
rect 208094 602061 208099 602106
rect 208493 602103 208559 602106
rect 208033 602056 208099 602061
rect 208350 600262 208356 600264
rect 208036 600230 208356 600262
rect 208033 600225 208356 600230
rect 208033 600169 208038 600225
rect 208094 600202 208356 600225
rect 208094 600169 208099 600202
rect 208350 600200 208356 600202
rect 208420 600200 208426 600264
rect 208033 600164 208099 600169
rect 244649 599582 244715 599585
rect 244649 599580 252578 599582
rect 244649 599524 244654 599580
rect 244710 599524 252578 599580
rect 244649 599522 252578 599524
rect 244649 599519 244715 599522
rect 620009 597134 620075 597137
rect 619230 597132 620075 597134
rect 619230 597076 620014 597132
rect 620070 597076 620075 597132
rect 619230 597074 620075 597076
rect 620009 597071 620075 597074
rect 208401 596456 208467 596457
rect 208350 596454 208356 596456
rect 208036 596431 208356 596454
rect 208420 596452 208467 596456
rect 208033 596426 208356 596431
rect 208033 596370 208038 596426
rect 208094 596394 208356 596426
rect 208462 596396 208467 596452
rect 208094 596370 208099 596394
rect 208350 596392 208356 596394
rect 208420 596392 208467 596396
rect 208401 596391 208467 596392
rect 208033 596365 208099 596370
rect 250077 585438 250143 585441
rect 250077 585436 252578 585438
rect 250077 585380 250082 585436
rect 250138 585380 252578 585436
rect 250077 585378 252578 585380
rect 250077 585375 250143 585378
rect 209689 584214 209755 584217
rect 207946 584212 209755 584214
rect 207946 584156 209694 584212
rect 209750 584156 209755 584212
rect 207946 584154 209755 584156
rect 209689 584151 209755 584154
rect 208309 584078 208375 584081
rect 207946 584076 208375 584078
rect 207946 584020 208314 584076
rect 208370 584020 208375 584076
rect 207946 584018 208375 584020
rect 208309 584015 208375 584018
rect 619222 583744 619228 583808
rect 619292 583806 619298 583808
rect 619365 583806 619431 583809
rect 619292 583804 619431 583806
rect 619292 583748 619370 583804
rect 619426 583748 619431 583804
rect 619292 583746 619431 583748
rect 619292 583744 619298 583746
rect 619365 583743 619431 583746
rect 619038 583472 619044 583536
rect 619108 583534 619114 583536
rect 619273 583534 619339 583537
rect 619108 583532 619339 583534
rect 619108 583476 619278 583532
rect 619334 583476 619339 583532
rect 619108 583474 619339 583476
rect 619108 583472 619114 583474
rect 619273 583471 619339 583474
rect 619038 582928 619044 582992
rect 619108 582928 619114 582992
rect 676078 581568 676084 581632
rect 676148 581630 676154 581632
rect 676681 581630 676747 581633
rect 676148 581628 676747 581630
rect 676148 581572 676686 581628
rect 676742 581572 676747 581628
rect 676148 581570 676747 581572
rect 676148 581568 676154 581570
rect 676681 581567 676747 581570
rect 676262 581432 676268 581496
rect 676332 581494 676338 581496
rect 676589 581494 676655 581497
rect 676332 581492 676655 581494
rect 676332 581436 676594 581492
rect 676650 581436 676655 581492
rect 676332 581434 676655 581436
rect 676332 581432 676338 581434
rect 676589 581431 676655 581434
rect 252142 578304 252148 578368
rect 252212 578366 252218 578368
rect 252212 578306 252578 578366
rect 252212 578304 252218 578306
rect 207934 577473 208106 577539
rect 208046 577414 208106 577473
rect 208861 577414 208927 577417
rect 208046 577412 208927 577414
rect 208046 577356 208866 577412
rect 208922 577356 208927 577412
rect 208046 577354 208927 577356
rect 208861 577351 208927 577354
rect 208493 576054 208559 576057
rect 208036 576052 208559 576054
rect 208036 576037 208498 576052
rect 208033 576032 208498 576037
rect 208033 575976 208038 576032
rect 208094 575996 208498 576032
rect 208554 575996 208559 576052
rect 208094 575994 208559 575996
rect 208094 575976 208099 575994
rect 208493 575991 208559 575994
rect 208033 575971 208099 575976
rect 619038 575856 619044 575920
rect 619108 575856 619114 575920
rect 208033 575442 208099 575445
rect 208033 575440 208234 575442
rect 208033 575384 208038 575440
rect 208094 575384 208234 575440
rect 208033 575382 208234 575384
rect 208033 575379 208099 575382
rect 208174 575374 208234 575382
rect 208309 575374 208375 575377
rect 208174 575372 208375 575374
rect 208174 575316 208314 575372
rect 208370 575316 208375 575372
rect 208174 575314 208375 575316
rect 208309 575311 208375 575314
rect 619038 575312 619044 575376
rect 619108 575374 619114 575376
rect 619273 575374 619339 575377
rect 619108 575372 619339 575374
rect 619108 575316 619278 575372
rect 619334 575316 619339 575372
rect 619108 575314 619339 575316
rect 619108 575312 619114 575314
rect 619273 575311 619339 575314
rect 676262 575040 676268 575104
rect 676332 575040 676338 575104
rect 675761 574830 675827 574833
rect 676270 574830 676330 575040
rect 675761 574828 676330 574830
rect 675761 574772 675766 574828
rect 675822 574772 676330 574828
rect 675761 574770 676330 574772
rect 675761 574767 675827 574770
rect 208861 574558 208927 574561
rect 208174 574556 208927 574558
rect 208033 574506 208099 574509
rect 208174 574506 208866 574556
rect 208033 574504 208866 574506
rect 208033 574448 208038 574504
rect 208094 574500 208866 574504
rect 208922 574500 208927 574556
rect 208094 574498 208927 574500
rect 208094 574448 208234 574498
rect 208861 574495 208927 574498
rect 208033 574446 208234 574448
rect 208033 574443 208099 574446
rect 208033 574054 208099 574057
rect 208033 574052 208234 574054
rect 208033 573996 208038 574052
rect 208094 574014 208234 574052
rect 208401 574014 208467 574017
rect 208094 574012 208467 574014
rect 208094 573996 208406 574012
rect 208033 573994 208406 573996
rect 208033 573991 208099 573994
rect 208174 573956 208406 573994
rect 208462 573956 208467 574012
rect 208174 573954 208467 573956
rect 208401 573951 208467 573954
rect 675485 574014 675551 574017
rect 676078 574014 676084 574016
rect 675485 574012 676084 574014
rect 675485 573956 675490 574012
rect 675546 573956 676084 574012
rect 675485 573954 676084 573956
rect 675485 573951 675551 573954
rect 676078 573952 676084 573954
rect 676148 573952 676154 574016
rect 675393 572246 675459 572249
rect 675853 572246 675919 572249
rect 675393 572244 676333 572246
rect 675393 572188 675398 572244
rect 675454 572188 675858 572244
rect 675914 572188 676333 572244
rect 675393 572186 676333 572188
rect 675393 572183 675459 572186
rect 675853 572183 675919 572186
rect 676273 572127 676333 572186
rect 676273 572061 676466 572127
rect 676273 572050 676333 572061
rect 619222 571912 619228 571976
rect 619292 571974 619298 571976
rect 619365 571974 619431 571977
rect 619292 571972 619431 571974
rect 619292 571916 619370 571972
rect 619426 571916 619431 571972
rect 619292 571914 619431 571916
rect 619292 571912 619298 571914
rect 619365 571911 619431 571914
rect 208033 571618 208099 571621
rect 208033 571616 208234 571618
rect 208033 571560 208038 571616
rect 208094 571566 208234 571616
rect 208861 571566 208927 571569
rect 208094 571564 208927 571566
rect 208094 571560 208866 571564
rect 208033 571558 208866 571560
rect 208033 571555 208099 571558
rect 208174 571508 208866 571558
rect 208922 571508 208927 571564
rect 208174 571506 208927 571508
rect 208861 571503 208927 571506
rect 623413 568846 623479 568849
rect 619230 568844 623479 568846
rect 619230 568788 623418 568844
rect 623474 568788 623479 568844
rect 619230 568786 623479 568788
rect 623413 568783 623479 568786
rect 676221 565582 676287 565585
rect 676221 565580 676453 565582
rect 676221 565524 676226 565580
rect 676282 565524 676453 565580
rect 676221 565522 676453 565524
rect 676221 565519 676287 565522
rect 670793 565446 670859 565449
rect 670793 565444 676453 565446
rect 670793 565388 670798 565444
rect 670854 565388 676453 565444
rect 670793 565386 676453 565388
rect 670793 565383 670859 565386
rect 251958 564160 251964 564224
rect 252028 564222 252034 564224
rect 252028 564162 252578 564222
rect 252028 564160 252034 564162
rect 622585 561774 622651 561777
rect 619230 561772 622651 561774
rect 619230 561716 622590 561772
rect 622646 561716 622651 561772
rect 619230 561714 622651 561716
rect 622585 561711 622651 561714
rect 244649 557150 244715 557153
rect 207806 557090 209982 557150
rect 207806 556811 207866 557090
rect 207806 556751 208006 556811
rect 209922 556742 209982 557090
rect 244649 557148 252578 557150
rect 244649 557092 244654 557148
rect 244710 557092 252578 557148
rect 244649 557090 252578 557092
rect 244649 557087 244715 557090
rect 211529 556742 211595 556745
rect 209922 556740 211595 556742
rect 209922 556684 211534 556740
rect 211590 556684 211595 556740
rect 209922 556682 211595 556684
rect 207933 556679 208099 556682
rect 211529 556679 211595 556682
rect 207905 556677 208099 556679
rect 207905 556621 208038 556677
rect 208094 556621 208099 556677
rect 207905 556619 208099 556621
rect 207933 556616 208099 556619
rect 208534 555592 208540 555656
rect 208604 555654 208610 555656
rect 209413 555654 209479 555657
rect 208604 555652 209479 555654
rect 208604 555596 209418 555652
rect 209474 555596 209479 555652
rect 208604 555594 209479 555596
rect 208604 555592 208610 555594
rect 209413 555591 209479 555594
rect 619089 551302 619155 551305
rect 619222 551302 619228 551304
rect 619089 551300 619228 551302
rect 619089 551244 619094 551300
rect 619150 551244 619228 551300
rect 619089 551242 619228 551244
rect 619089 551239 619155 551242
rect 619222 551240 619228 551242
rect 619292 551240 619298 551304
rect 208125 550136 208191 550139
rect 207946 550134 208191 550136
rect 207946 550078 208130 550134
rect 208186 550078 208191 550134
rect 207946 550076 208191 550078
rect 208125 550073 208191 550076
rect 248053 550078 248119 550081
rect 248053 550076 252578 550078
rect 248053 550020 248058 550076
rect 248114 550020 252578 550076
rect 248053 550018 252578 550020
rect 248053 550015 248119 550018
rect 620009 547630 620075 547633
rect 619230 547628 620075 547630
rect 619230 547572 620014 547628
rect 620070 547572 620075 547628
rect 619230 547570 620075 547572
rect 620009 547567 620075 547570
rect 208033 546812 208099 546817
rect 208033 546756 208038 546812
rect 208094 546756 208099 546812
rect 208033 546751 208099 546756
rect 208036 546545 208096 546751
rect 208033 546540 208099 546545
rect 208033 546484 208038 546540
rect 208094 546484 208099 546540
rect 208033 546479 208099 546484
rect 208534 545454 208540 545456
rect 208033 545427 208099 545430
rect 208174 545427 208540 545454
rect 208033 545425 208540 545427
rect 208033 545369 208038 545425
rect 208094 545394 208540 545425
rect 208094 545369 208234 545394
rect 208534 545392 208540 545394
rect 208604 545392 208610 545456
rect 208033 545367 208234 545369
rect 208033 545364 208099 545367
rect 208033 544230 208099 544233
rect 208769 544230 208835 544233
rect 208033 544228 208835 544230
rect 208033 544172 208038 544228
rect 208094 544172 208774 544228
rect 208830 544172 208835 544228
rect 208033 544170 208835 544172
rect 208033 544167 208099 544170
rect 208769 544167 208835 544170
rect 208585 543550 208651 543553
rect 208174 543548 208651 543550
rect 208033 543507 208099 543510
rect 208174 543507 208590 543548
rect 208033 543505 208590 543507
rect 208033 543449 208038 543505
rect 208094 543492 208590 543505
rect 208646 543492 208651 543548
rect 208094 543490 208651 543492
rect 208094 543449 208234 543490
rect 208585 543487 208651 543490
rect 208033 543447 208234 543449
rect 208033 543444 208099 543447
rect 246778 543064 246908 543074
rect 246778 542964 246793 543064
rect 246889 543042 246908 543064
rect 246889 542982 252603 543042
rect 246889 542964 246908 542982
rect 246778 542949 246908 542964
rect 619273 542054 619339 542057
rect 619406 542054 619412 542056
rect 619273 542052 619412 542054
rect 619273 541996 619278 542052
rect 619334 541996 619412 542052
rect 619273 541994 619412 541996
rect 619273 541991 619339 541994
rect 619406 541992 619412 541994
rect 619476 541992 619482 542056
rect 208493 541646 208559 541649
rect 208174 541644 208559 541646
rect 208033 541628 208099 541631
rect 208174 541628 208498 541644
rect 208033 541626 208498 541628
rect 208033 541570 208038 541626
rect 208094 541588 208498 541626
rect 208554 541588 208559 541644
rect 208094 541586 208559 541588
rect 208094 541570 208234 541586
rect 208493 541583 208559 541586
rect 208033 541568 208234 541570
rect 208033 541565 208099 541568
rect 619590 540558 619596 540560
rect 619230 540498 619596 540558
rect 619590 540496 619596 540498
rect 619660 540496 619666 540560
rect 676221 537836 676287 537841
rect 676221 537780 676226 537836
rect 676282 537780 676287 537836
rect 676221 537775 676287 537780
rect 676224 537705 676284 537775
rect 676221 537700 676287 537705
rect 676221 537644 676226 537700
rect 676282 537644 676287 537700
rect 676221 537639 676287 537644
rect 675894 536144 675900 536208
rect 675964 536206 675970 536208
rect 676221 536206 676287 536209
rect 675964 536204 676287 536206
rect 675964 536148 676226 536204
rect 676282 536148 676287 536204
rect 675964 536146 676287 536148
rect 675964 536144 675970 536146
rect 676221 536143 676287 536146
rect 676078 536008 676084 536072
rect 676148 536070 676154 536072
rect 676303 536070 676369 536073
rect 676148 536068 676369 536070
rect 676148 536012 676308 536068
rect 676364 536012 676369 536068
rect 676148 536010 676369 536012
rect 676148 536008 676154 536010
rect 676303 536007 676369 536010
rect 252009 535662 252075 535665
rect 252009 535660 252578 535662
rect 252009 535604 252014 535660
rect 252070 535604 252578 535660
rect 252009 535602 252578 535604
rect 252009 535599 252075 535602
rect 675894 534920 675900 534984
rect 675964 534982 675970 534984
rect 676221 534982 676287 534985
rect 675964 534980 676287 534982
rect 675964 534924 676226 534980
rect 676282 534924 676287 534980
rect 675964 534922 676287 534924
rect 675964 534920 675970 534922
rect 676221 534919 676287 534922
rect 675894 534104 675900 534168
rect 675964 534166 675970 534168
rect 675964 534157 676284 534166
rect 675964 534152 676287 534157
rect 675964 534106 676226 534152
rect 675964 534104 675970 534106
rect 676221 534096 676226 534106
rect 676282 534096 676287 534152
rect 676221 534091 676287 534096
rect 619406 533486 619412 533488
rect 619230 533426 619412 533486
rect 619406 533424 619412 533426
rect 619476 533424 619482 533488
rect 675761 532534 675827 532537
rect 676262 532534 676268 532536
rect 675761 532532 676268 532534
rect 675761 532476 675766 532532
rect 675822 532476 676268 532532
rect 675761 532474 676268 532476
rect 675761 532471 675827 532474
rect 676262 532472 676268 532474
rect 676332 532472 676338 532536
rect 675894 531062 675900 531126
rect 675964 531124 675970 531126
rect 675964 531064 676453 531124
rect 675964 531062 675970 531064
rect 675669 530086 675735 530089
rect 675894 530086 675900 530088
rect 675669 530084 675900 530086
rect 675669 530028 675674 530084
rect 675730 530028 675900 530084
rect 675669 530026 675900 530028
rect 675669 530023 675735 530026
rect 675894 530024 675900 530026
rect 675964 530024 675970 530088
rect 208033 529542 208099 529545
rect 208033 529540 208234 529542
rect 208033 529484 208038 529540
rect 208094 529484 208234 529540
rect 208033 529482 208234 529484
rect 208033 529479 208099 529482
rect 208174 529280 208234 529482
rect 208677 529280 208743 529283
rect 207946 529278 208743 529280
rect 207946 529222 208682 529278
rect 208738 529222 208743 529278
rect 207946 529220 208743 529222
rect 208677 529217 208743 529220
rect 208677 526958 208743 526961
rect 208036 526956 208743 526958
rect 208036 526926 208682 526956
rect 208033 526921 208682 526926
rect 208033 526865 208038 526921
rect 208094 526900 208682 526921
rect 208738 526900 208743 526956
rect 208094 526898 208743 526900
rect 208094 526865 208099 526898
rect 208677 526895 208743 526898
rect 619181 526958 619247 526961
rect 619181 526956 619290 526958
rect 619181 526900 619186 526956
rect 619242 526900 619290 526956
rect 619181 526895 619290 526900
rect 208033 526860 208099 526865
rect 619230 526354 619290 526895
rect 675761 524646 675827 524649
rect 676262 524646 676268 524648
rect 675761 524644 676268 524646
rect 675761 524588 675766 524644
rect 675822 524588 676268 524644
rect 675761 524586 676268 524588
rect 675761 524583 675827 524586
rect 676262 524584 676268 524586
rect 676332 524584 676338 524648
rect 676270 524581 676338 524584
rect 676270 524521 676453 524581
rect 675902 524389 676453 524449
rect 674197 524374 674263 524377
rect 675902 524374 675962 524389
rect 674197 524372 675962 524374
rect 674197 524316 674202 524372
rect 674258 524316 675962 524372
rect 674197 524314 675962 524316
rect 674197 524311 674263 524314
rect 676078 524040 676084 524104
rect 676148 524102 676154 524104
rect 676589 524102 676655 524105
rect 676148 524100 676655 524102
rect 676148 524044 676594 524100
rect 676650 524044 676655 524100
rect 676148 524042 676655 524044
rect 676148 524040 676154 524042
rect 676589 524039 676655 524042
rect 208086 522739 208146 522742
rect 207934 522673 208146 522739
rect 208086 522606 208146 522673
rect 208217 522606 208283 522609
rect 208493 522606 208559 522609
rect 208086 522604 208559 522606
rect 208086 522548 208222 522604
rect 208278 522548 208498 522604
rect 208554 522548 208559 522604
rect 208086 522546 208559 522548
rect 208217 522543 208283 522546
rect 208493 522543 208559 522546
rect 250997 521518 251063 521521
rect 250997 521516 252578 521518
rect 250997 521460 251002 521516
rect 251058 521460 252578 521516
rect 250997 521458 252578 521460
rect 250997 521455 251063 521458
rect 619089 519886 619155 519889
rect 619046 519884 619155 519886
rect 619046 519828 619094 519884
rect 619150 519828 619155 519884
rect 619046 519823 619155 519828
rect 208033 519478 208099 519481
rect 208677 519478 208743 519481
rect 208033 519476 208743 519478
rect 208033 519420 208038 519476
rect 208094 519420 208682 519476
rect 208738 519420 208743 519476
rect 208033 519418 208743 519420
rect 208033 519415 208099 519418
rect 208677 519415 208743 519418
rect 619046 519282 619106 519823
rect 208309 518934 208375 518937
rect 208036 518932 208375 518934
rect 208036 518876 208314 518932
rect 208370 518876 208375 518932
rect 208036 518874 208375 518876
rect 208036 518869 208099 518874
rect 208309 518871 208375 518874
rect 208033 518864 208099 518869
rect 208033 518808 208038 518864
rect 208094 518808 208099 518864
rect 208033 518803 208099 518808
rect 208033 516105 208099 516110
rect 208033 516049 208038 516105
rect 208094 516078 208099 516105
rect 208309 516078 208375 516081
rect 208094 516076 208375 516078
rect 208094 516049 208314 516076
rect 208033 516044 208314 516049
rect 208036 516020 208314 516044
rect 208370 516020 208375 516076
rect 208036 516018 208375 516020
rect 208309 516015 208375 516018
rect 250813 514446 250879 514449
rect 250813 514444 252578 514446
rect 250813 514388 250818 514444
rect 250874 514388 252578 514444
rect 250813 514386 252578 514388
rect 250813 514383 250879 514386
rect 252469 507646 252535 507649
rect 252334 507644 252535 507646
rect 252334 507588 252474 507644
rect 252530 507588 252535 507644
rect 252334 507586 252535 507588
rect 252334 507374 252394 507586
rect 252469 507583 252535 507586
rect 252334 507314 252578 507374
rect 619457 504926 619523 504929
rect 619230 504924 619523 504926
rect 619230 504868 619462 504924
rect 619518 504868 619523 504924
rect 619230 504866 619523 504868
rect 619457 504863 619523 504866
rect 207946 502006 208174 502011
rect 207946 501951 208094 502006
rect 208089 501950 208094 501951
rect 208150 501950 208174 502006
rect 208089 501946 208174 501950
rect 208089 501945 208155 501946
rect 208493 501879 208559 501882
rect 207946 501877 208559 501879
rect 207946 501821 208498 501877
rect 208554 501821 208559 501877
rect 207946 501819 208559 501821
rect 208493 501816 208559 501819
rect 246857 500302 246923 500305
rect 246857 500300 252578 500302
rect 246857 500244 246862 500300
rect 246918 500244 252578 500300
rect 246857 500242 252578 500244
rect 246857 500239 246923 500242
rect 208033 499521 208099 499526
rect 208033 499465 208038 499521
rect 208094 499486 208099 499521
rect 208677 499486 208743 499489
rect 208094 499484 208743 499486
rect 208094 499465 208682 499484
rect 208033 499460 208682 499465
rect 208036 499428 208682 499460
rect 208738 499428 208743 499484
rect 208036 499426 208743 499428
rect 208677 499423 208743 499426
rect 621389 497854 621455 497857
rect 619230 497852 621455 497854
rect 619230 497796 621394 497852
rect 621450 497796 621455 497852
rect 619230 497794 621455 497796
rect 621389 497791 621455 497794
rect 208033 496125 208099 496130
rect 208033 496069 208038 496125
rect 208094 496086 208099 496125
rect 208677 496086 208743 496089
rect 208861 496086 208927 496089
rect 208094 496084 208927 496086
rect 208094 496069 208682 496084
rect 208033 496064 208682 496069
rect 208036 496028 208682 496064
rect 208738 496028 208866 496084
rect 208922 496028 208927 496084
rect 208036 496026 208927 496028
rect 208677 496023 208743 496026
rect 208861 496023 208927 496026
rect 207934 495336 208206 495339
rect 207866 495276 208206 495336
rect 207934 495273 208206 495276
rect 208140 495134 208206 495273
rect 208401 495134 208467 495137
rect 208677 495134 208743 495137
rect 208139 495132 208743 495134
rect 208139 495076 208406 495132
rect 208462 495076 208682 495132
rect 208738 495076 208743 495132
rect 208139 495074 208743 495076
rect 208401 495071 208467 495074
rect 208677 495071 208743 495074
rect 208585 493322 208651 493325
rect 208542 493320 208651 493322
rect 208542 493264 208590 493320
rect 208646 493264 208651 493320
rect 208542 493259 208651 493264
rect 208033 493230 208099 493233
rect 208542 493230 208602 493259
rect 208033 493228 208602 493230
rect 208033 493172 208038 493228
rect 208094 493172 208602 493228
rect 208033 493170 208602 493172
rect 248973 493230 249039 493233
rect 248973 493228 252578 493230
rect 248973 493172 248978 493228
rect 249034 493172 252578 493228
rect 248973 493170 252578 493172
rect 208033 493167 208099 493170
rect 248973 493167 249039 493170
rect 208769 492550 208835 492553
rect 208174 492548 208835 492550
rect 208033 492519 208099 492522
rect 208174 492519 208774 492548
rect 208033 492517 208774 492519
rect 208033 492461 208038 492517
rect 208094 492492 208774 492517
rect 208830 492492 208835 492548
rect 208094 492490 208835 492492
rect 208094 492461 208234 492490
rect 208769 492487 208835 492490
rect 208033 492459 208234 492461
rect 208033 492456 208099 492459
rect 619046 490241 619106 490782
rect 675301 490374 675367 490377
rect 675301 490372 676146 490374
rect 675301 490316 675306 490372
rect 675362 490324 676146 490372
rect 675362 490322 676453 490324
rect 675362 490316 676042 490322
rect 675301 490314 676042 490316
rect 675301 490311 675367 490314
rect 675956 490266 676042 490314
rect 676098 490266 676453 490322
rect 675956 490264 676453 490266
rect 676037 490261 676103 490264
rect 619046 490236 619155 490241
rect 619046 490180 619094 490236
rect 619150 490180 619155 490236
rect 619046 490178 619155 490180
rect 619089 490175 619155 490178
rect 208861 486838 208927 486841
rect 208036 486836 208927 486838
rect 208036 486831 208866 486836
rect 208033 486826 208866 486831
rect 208033 486770 208038 486826
rect 208094 486780 208866 486826
rect 208922 486780 208927 486836
rect 208094 486778 208927 486780
rect 208094 486770 208099 486778
rect 208861 486775 208927 486778
rect 208033 486765 208099 486770
rect 676129 486430 676195 486433
rect 676262 486430 676268 486432
rect 676129 486428 676268 486430
rect 676129 486372 676134 486428
rect 676190 486372 676268 486428
rect 676129 486370 676268 486372
rect 676129 486367 676195 486370
rect 676262 486368 676268 486370
rect 676332 486368 676338 486432
rect 252285 486158 252351 486161
rect 252285 486156 252578 486158
rect 252285 486100 252290 486156
rect 252346 486100 252578 486156
rect 252285 486098 252578 486100
rect 252285 486095 252351 486098
rect 676262 483719 676268 483783
rect 676332 483781 676338 483783
rect 676332 483721 676453 483781
rect 676332 483719 676338 483721
rect 676393 483589 676514 483649
rect 676129 483438 676195 483441
rect 676454 483438 676514 483589
rect 676129 483436 676514 483438
rect 676129 483380 676134 483436
rect 676190 483380 676514 483436
rect 676129 483378 676514 483380
rect 676129 483375 676195 483378
rect 250813 479086 250879 479089
rect 250813 479084 252578 479086
rect 250813 479028 250818 479084
rect 250874 479028 252578 479084
rect 250813 479026 252578 479028
rect 250813 479023 250879 479026
rect 211161 474598 211227 474601
rect 207946 474596 211227 474598
rect 207946 474540 211166 474596
rect 211222 474540 211227 474596
rect 207946 474538 211227 474540
rect 207946 474351 208006 474538
rect 211161 474535 211227 474538
rect 207934 474279 208150 474282
rect 207934 474216 208156 474279
rect 208096 474190 208156 474216
rect 208585 474190 208651 474193
rect 208861 474190 208927 474193
rect 208096 474188 208927 474190
rect 208096 474132 208590 474188
rect 208646 474132 208866 474188
rect 208922 474132 208927 474188
rect 208096 474130 208927 474132
rect 208585 474127 208651 474130
rect 208861 474127 208927 474130
rect 252193 472014 252259 472017
rect 252193 472012 252578 472014
rect 252193 471956 252198 472012
rect 252254 471956 252578 472012
rect 252193 471954 252578 471956
rect 252193 471951 252259 471954
rect 620101 469566 620167 469569
rect 619230 469564 620167 469566
rect 619230 469508 620106 469564
rect 620162 469508 620167 469564
rect 619230 469506 620167 469508
rect 620101 469503 620167 469506
rect 209045 467934 209111 467937
rect 208096 467932 209111 467934
rect 208096 467876 209050 467932
rect 209106 467876 209111 467932
rect 208096 467874 209111 467876
rect 208096 467739 208156 467874
rect 209045 467871 209111 467874
rect 207934 467673 208156 467739
rect 251089 464942 251155 464945
rect 251089 464940 252578 464942
rect 251089 464884 251094 464940
rect 251150 464884 252578 464940
rect 251089 464882 252578 464884
rect 251089 464879 251155 464882
rect 622401 462494 622467 462497
rect 619230 462492 622467 462494
rect 619230 462436 622406 462492
rect 622462 462436 622467 462492
rect 619230 462434 622467 462436
rect 622401 462431 622467 462434
rect 208033 461814 208099 461817
rect 208861 461814 208927 461817
rect 208033 461812 208927 461814
rect 208033 461756 208038 461812
rect 208094 461756 208866 461812
rect 208922 461756 208927 461812
rect 208033 461754 208927 461756
rect 208033 461751 208099 461754
rect 208861 461751 208927 461754
rect 208033 459782 208099 459785
rect 208033 459780 208234 459782
rect 208033 459724 208038 459780
rect 208094 459724 208234 459780
rect 208033 459722 208234 459724
rect 208033 459719 208099 459722
rect 208033 459638 208099 459641
rect 208174 459638 208234 459722
rect 208585 459638 208651 459641
rect 208861 459638 208927 459641
rect 208033 459636 208927 459638
rect 208033 459580 208038 459636
rect 208094 459580 208590 459636
rect 208646 459580 208866 459636
rect 208922 459580 208927 459636
rect 208033 459578 208927 459580
rect 208033 459575 208099 459578
rect 208585 459575 208651 459578
rect 208861 459575 208927 459578
rect 208677 459366 208743 459369
rect 208174 459364 208743 459366
rect 208174 459308 208682 459364
rect 208738 459308 208743 459364
rect 208174 459306 208743 459308
rect 208174 459101 208234 459306
rect 208677 459303 208743 459306
rect 208125 459096 208234 459101
rect 208125 459040 208130 459096
rect 208186 459040 208234 459096
rect 208125 459038 208234 459040
rect 208125 459035 208191 459038
rect 641874 458408 676910 458600
rect 209070 457870 209146 457876
rect 209070 457866 252602 457870
rect 209070 457810 209080 457866
rect 209136 457810 252602 457866
rect 209070 457806 252602 457810
rect 209070 457801 209146 457806
rect 623321 455422 623387 455425
rect 619230 455420 623387 455422
rect 619230 455364 623326 455420
rect 623382 455364 623387 455420
rect 619230 455362 623387 455364
rect 623321 455359 623387 455362
rect 641874 454112 642378 458408
rect 648850 454112 676910 458408
rect 641874 453800 676910 454112
rect 642378 452696 648850 452862
rect 641794 448278 676910 448549
rect 210425 447126 210491 447129
rect 207946 447124 210491 447126
rect 207946 447068 210430 447124
rect 210486 447068 210491 447124
rect 207946 447066 210491 447068
rect 207946 446948 208006 447066
rect 210425 447063 210491 447066
rect 207946 446854 208234 446888
rect 208585 446854 208651 446857
rect 207946 446852 208651 446854
rect 207946 446828 208590 446852
rect 208174 446796 208590 446828
rect 208646 446796 208651 446852
rect 208174 446794 208651 446796
rect 208585 446791 208651 446794
rect 641794 443982 642404 448278
rect 648876 443982 676910 448278
rect 641794 443760 676910 443982
rect 252377 443726 252443 443729
rect 252377 443724 252578 443726
rect 252377 443668 252382 443724
rect 252438 443668 252578 443724
rect 252377 443666 252578 443668
rect 252377 443663 252443 443666
rect 620193 441278 620259 441281
rect 619230 441276 620259 441278
rect 619230 441220 620198 441276
rect 620254 441220 620259 441276
rect 619230 441218 620259 441220
rect 620193 441215 620259 441218
rect 208585 441142 208651 441145
rect 208036 441140 208651 441142
rect 208036 441130 208590 441140
rect 208033 441125 208590 441130
rect 208033 441069 208038 441125
rect 208094 441084 208590 441125
rect 208646 441084 208651 441140
rect 208094 441082 208651 441084
rect 208094 441069 208099 441082
rect 208585 441079 208651 441082
rect 208033 441064 208099 441069
rect 208217 440336 208283 440339
rect 208769 440336 208835 440339
rect 207946 440334 208835 440336
rect 207946 440278 208222 440334
rect 208278 440278 208774 440334
rect 208830 440278 208835 440334
rect 207946 440276 208835 440278
rect 208217 440273 208283 440276
rect 208769 440273 208835 440276
rect 208033 438832 208099 438837
rect 208033 438776 208038 438832
rect 208094 438830 208099 438832
rect 208401 438830 208467 438833
rect 208094 438828 208467 438830
rect 208094 438776 208406 438828
rect 208033 438772 208406 438776
rect 208462 438772 208467 438828
rect 208033 438771 208467 438772
rect 208036 438770 208467 438771
rect 208401 438767 208467 438770
rect 247317 436654 247383 436657
rect 247317 436652 252578 436654
rect 247317 436596 247322 436652
rect 247378 436596 252578 436652
rect 247317 436594 252578 436596
rect 247317 436591 247383 436594
rect 623229 434206 623295 434209
rect 619230 434204 623295 434206
rect 619230 434148 623234 434204
rect 623290 434148 623295 434204
rect 619230 434146 623295 434148
rect 623229 434143 623295 434146
rect 208033 431826 208099 431829
rect 208033 431824 208234 431826
rect 208033 431768 208038 431824
rect 208094 431768 208234 431824
rect 208033 431766 208234 431768
rect 208033 431763 208099 431766
rect 208174 431758 208234 431766
rect 208677 431758 208743 431761
rect 208861 431758 208927 431761
rect 208174 431756 208927 431758
rect 208174 431700 208682 431756
rect 208738 431700 208866 431756
rect 208922 431700 208927 431756
rect 208174 431698 208927 431700
rect 208677 431695 208743 431698
rect 208861 431695 208927 431698
rect 252101 429582 252167 429585
rect 252101 429580 252578 429582
rect 252101 429524 252106 429580
rect 252162 429524 252578 429580
rect 252101 429522 252578 429524
rect 252101 429519 252167 429522
rect 621205 427134 621271 427137
rect 619230 427132 621271 427134
rect 619230 427076 621210 427132
rect 621266 427076 621271 427132
rect 619230 427074 621271 427076
rect 621205 427071 621271 427074
rect 250813 422510 250879 422513
rect 250813 422508 252578 422510
rect 250813 422452 250818 422508
rect 250874 422452 252578 422508
rect 250813 422450 252578 422452
rect 250813 422447 250879 422450
rect 620193 420062 620259 420065
rect 619230 420060 620259 420062
rect 619230 420004 620198 420060
rect 620254 420004 620259 420060
rect 619230 420002 620259 420004
rect 620193 419999 620259 420002
rect 641678 418576 676548 418801
rect 249249 415438 249315 415441
rect 249249 415436 252578 415438
rect 249249 415380 249254 415436
rect 249310 415380 252578 415436
rect 249249 415378 252578 415380
rect 249249 415375 249315 415378
rect 641678 414218 642392 418576
rect 648886 414218 676548 418576
rect 641678 414021 676548 414218
rect 622309 412990 622375 412993
rect 619230 412988 622375 412990
rect 619230 412932 622314 412988
rect 622370 412932 622375 412988
rect 619230 412930 622375 412932
rect 622309 412927 622375 412930
rect 641678 408620 676548 408822
rect 207990 406380 208144 406484
rect 619181 406462 619247 406465
rect 619181 406460 619290 406462
rect 619181 406404 619186 406460
rect 619242 406404 619290 406460
rect 619181 406399 619290 406404
rect 619230 405858 619290 406399
rect 641678 404262 642392 408620
rect 648886 404262 676548 408620
rect 641678 404042 676548 404262
rect 250261 401022 250327 401025
rect 250261 401020 252578 401022
rect 250261 400964 250266 401020
rect 250322 400964 252578 401020
rect 250261 400962 252578 400964
rect 250261 400959 250327 400962
rect 623137 398846 623203 398849
rect 619230 398844 623203 398846
rect 619230 398788 623142 398844
rect 623198 398788 623203 398844
rect 619230 398786 623203 398788
rect 623137 398783 623203 398786
rect 251273 393950 251339 393953
rect 251273 393948 252578 393950
rect 251273 393892 251278 393948
rect 251334 393892 252578 393948
rect 251273 393890 252578 393892
rect 251273 393887 251339 393890
rect 208861 393134 208927 393137
rect 208174 393132 208927 393134
rect 208174 393079 208866 393132
rect 207946 393076 208866 393079
rect 208922 393076 208927 393132
rect 207946 393074 208927 393076
rect 207946 393019 208234 393074
rect 208861 393071 208927 393074
rect 250077 386878 250143 386881
rect 250077 386876 252578 386878
rect 250077 386820 250082 386876
rect 250138 386820 252578 386876
rect 250077 386818 252578 386820
rect 250077 386815 250143 386818
rect 208125 386536 208191 386539
rect 207946 386534 208191 386536
rect 207946 386478 208130 386534
rect 208186 386478 208191 386534
rect 207946 386476 208191 386478
rect 208125 386473 208191 386476
rect 621021 384430 621087 384433
rect 619230 384428 621087 384430
rect 619230 384372 621026 384428
rect 621082 384372 621087 384428
rect 619230 384370 621087 384372
rect 621021 384367 621087 384370
rect 208493 383750 208559 383753
rect 208174 383748 208559 383750
rect 208033 383719 208099 383722
rect 208174 383719 208498 383748
rect 208033 383717 208498 383719
rect 208033 383661 208038 383717
rect 208094 383692 208498 383717
rect 208554 383692 208559 383748
rect 208094 383690 208559 383692
rect 208094 383661 208234 383690
rect 208493 383687 208559 383690
rect 208033 383659 208234 383661
rect 208033 383656 208099 383659
rect 627548 378694 676460 378801
rect 627548 374174 629506 378694
rect 636022 374174 676460 378694
rect 627548 374021 676460 374174
rect 620193 370286 620259 370289
rect 619230 370284 620259 370286
rect 619230 370228 620198 370284
rect 620254 370228 620259 370284
rect 619230 370226 620259 370228
rect 620193 370223 620259 370226
rect 627548 368714 676548 368822
rect 207824 365470 244070 365758
rect 250353 365662 250419 365665
rect 250353 365660 252578 365662
rect 250353 365604 250358 365660
rect 250414 365604 252578 365660
rect 250353 365602 252578 365604
rect 250353 365599 250419 365602
rect 207824 361160 236392 365470
rect 242928 361160 244070 365470
rect 627548 364194 629506 368714
rect 636022 364194 676548 368714
rect 627548 364042 676548 364194
rect 619222 363152 619228 363216
rect 619292 363152 619298 363216
rect 207824 360978 244070 361160
rect 236392 359874 242928 360978
rect 249341 358590 249407 358593
rect 249341 358588 252578 358590
rect 249341 358532 249346 358588
rect 249402 358532 252578 358588
rect 249341 358530 252578 358532
rect 249341 358527 249407 358530
rect 207824 355508 244128 355779
rect 207824 351198 236506 355508
rect 243042 351198 244128 355508
rect 252101 351518 252167 351521
rect 252101 351516 252578 351518
rect 252101 351460 252106 351516
rect 252162 351460 252578 351516
rect 252101 351458 252578 351460
rect 252101 351455 252167 351458
rect 207824 350999 244128 351198
rect 622217 349070 622283 349073
rect 619230 349068 622283 349070
rect 619230 349012 622222 349068
rect 622278 349012 622283 349068
rect 619230 349010 622283 349012
rect 622217 349007 622283 349010
rect 252653 344718 252719 344721
rect 252380 344716 252719 344718
rect 252380 344660 252658 344716
rect 252714 344660 252719 344716
rect 252380 344658 252719 344660
rect 252380 344446 252440 344658
rect 252653 344655 252719 344658
rect 252380 344386 252578 344446
rect 620929 341998 620995 342001
rect 619230 341996 620995 341998
rect 619230 341940 620934 341996
rect 620990 341940 620995 341996
rect 619230 341938 620995 341940
rect 620929 341935 620995 341938
rect 207438 339360 223360 339440
rect 207438 334842 215366 339360
rect 222020 334842 223360 339360
rect 665308 339000 670089 339052
rect 251917 337374 251983 337377
rect 251917 337372 252578 337374
rect 251917 337316 251922 337372
rect 251978 337316 252578 337372
rect 251917 337314 252578 337316
rect 251917 337311 251983 337314
rect 620837 334926 620903 334929
rect 619230 334924 620903 334926
rect 619230 334868 620842 334924
rect 620898 334868 620903 334924
rect 619230 334866 620903 334868
rect 620837 334863 620903 334866
rect 207438 334651 223360 334842
rect 665308 334200 676940 339000
rect 252285 330302 252351 330305
rect 252285 330300 252578 330302
rect 252285 330244 252290 330300
rect 252346 330244 252578 330300
rect 252285 330242 252578 330244
rect 252285 330239 252351 330242
rect 207438 329222 223360 329400
rect 207438 324704 215346 329222
rect 222000 324704 223360 329222
rect 665308 328949 670089 334200
rect 620694 327854 620700 327856
rect 619230 327794 620700 327854
rect 620694 327792 620700 327794
rect 620764 327792 620770 327856
rect 207438 324600 223360 324704
rect 665308 324160 676940 328949
rect 252193 323230 252259 323233
rect 252193 323228 252578 323230
rect 252193 323172 252198 323228
rect 252254 323172 252578 323228
rect 252193 323170 252578 323172
rect 252193 323167 252259 323170
rect 622125 320782 622191 320785
rect 619230 320780 622191 320782
rect 619230 320724 622130 320780
rect 622186 320724 622191 320780
rect 619230 320722 622191 320724
rect 622125 320719 622191 320722
rect 246305 316158 246371 316161
rect 246305 316156 252578 316158
rect 246305 316100 246310 316156
rect 246366 316100 252578 316156
rect 246305 316098 252578 316100
rect 246305 316095 246371 316098
rect 620101 313710 620167 313713
rect 619230 313708 620167 313710
rect 619230 313652 620106 313708
rect 620162 313652 620167 313708
rect 619230 313650 620167 313652
rect 620101 313647 620167 313650
rect 252193 309086 252259 309089
rect 252193 309084 252578 309086
rect 252193 309028 252198 309084
rect 252254 309028 252578 309084
rect 252193 309026 252578 309028
rect 252193 309023 252259 309026
rect 619406 306638 619412 306640
rect 619230 306578 619412 306638
rect 619406 306576 619412 306578
rect 619476 306576 619482 306640
rect 251774 301952 251780 302016
rect 251844 302014 251850 302016
rect 251844 301954 252578 302014
rect 251844 301952 251850 301954
rect 619038 299504 619044 299568
rect 619108 299504 619114 299568
rect 665308 299201 670089 324160
rect 252377 294942 252443 294945
rect 252377 294940 252578 294942
rect 252377 294884 252382 294940
rect 252438 294884 252578 294940
rect 252377 294882 252578 294884
rect 252377 294879 252443 294882
rect 665252 294421 676500 299201
rect 619917 292494 619983 292497
rect 619230 292492 619983 292494
rect 619230 292436 619922 292492
rect 619978 292436 619983 292492
rect 619230 292434 619983 292436
rect 619917 292431 619983 292434
rect 665308 289222 670089 294421
rect 231217 284742 231283 284745
rect 233609 284742 233675 284745
rect 231217 284740 233675 284742
rect 231217 284684 231222 284740
rect 231278 284684 233614 284740
rect 233670 284684 233675 284740
rect 231217 284682 233675 284684
rect 231217 284679 231283 284682
rect 233609 284679 233675 284682
rect 665308 284442 676500 289222
rect 232229 283790 232295 283793
rect 232229 283788 232338 283790
rect 232229 283732 232234 283788
rect 232290 283732 232338 283788
rect 232229 283727 232338 283732
rect 232278 283186 232338 283727
rect 228222 283116 228228 283180
rect 228292 283116 228298 283180
rect 634912 281126 636294 281152
rect 634912 280890 634944 281126
rect 636264 280890 636294 281126
rect 634912 280868 636294 280890
rect 642298 280916 643130 280936
rect 642298 280712 642326 280916
rect 643110 280712 643130 280916
rect 642298 280692 643130 280712
rect 226985 280526 227051 280529
rect 230205 280526 230271 280529
rect 226985 280524 230271 280526
rect 226985 280468 226990 280524
rect 227046 280468 230210 280524
rect 230266 280468 230271 280524
rect 226985 280466 230271 280468
rect 226985 280463 227051 280466
rect 230205 280463 230271 280466
rect 252285 280526 252351 280529
rect 674105 280526 674171 280529
rect 252285 280524 674171 280526
rect 252285 280468 252290 280524
rect 252346 280468 674110 280524
rect 674166 280468 674171 280524
rect 252285 280466 674171 280468
rect 252285 280463 252351 280466
rect 674105 280463 674171 280466
rect 240233 280118 240299 280121
rect 619406 280118 619412 280120
rect 240233 280116 619412 280118
rect 240233 280060 240238 280116
rect 240294 280060 619412 280116
rect 240233 280058 619412 280060
rect 240233 280055 240299 280058
rect 619406 280056 619412 280058
rect 619476 280056 619482 280120
rect 228222 279920 228228 279984
rect 228292 279982 228298 279984
rect 232321 279982 232387 279985
rect 228292 279980 232387 279982
rect 228292 279924 232326 279980
rect 232382 279924 232387 279980
rect 228292 279922 232387 279924
rect 228292 279920 228298 279922
rect 232321 279919 232387 279922
rect 244649 279982 244715 279985
rect 619222 279982 619228 279984
rect 244649 279980 619228 279982
rect 244649 279924 244654 279980
rect 244710 279924 619228 279980
rect 244649 279922 619228 279924
rect 244649 279919 244715 279922
rect 619222 279920 619228 279922
rect 619292 279920 619298 279984
rect 252510 279784 252516 279848
rect 252580 279846 252586 279848
rect 396633 279846 396699 279849
rect 252580 279844 396699 279846
rect 252580 279788 396638 279844
rect 396694 279788 396699 279844
rect 252580 279786 396699 279788
rect 252580 279784 252586 279786
rect 396633 279783 396699 279786
rect 252694 279648 252700 279712
rect 252764 279710 252770 279712
rect 276849 279710 276915 279713
rect 252764 279708 276915 279710
rect 252764 279652 276854 279708
rect 276910 279652 276915 279708
rect 252764 279650 276915 279652
rect 252764 279648 252770 279650
rect 276849 279647 276915 279650
rect 252326 278968 252332 279032
rect 252396 279030 252402 279032
rect 478145 279030 478211 279033
rect 252396 279028 478211 279030
rect 252396 278972 478150 279028
rect 478206 278972 478211 279028
rect 252396 278970 478211 278972
rect 252396 278968 252402 278970
rect 478145 278967 478211 278970
rect 236098 276276 365740 276332
rect 236098 273804 236380 276276
rect 243110 273804 365740 276276
rect 236098 273678 365740 273804
rect 286556 271806 292449 272236
rect 286556 265298 288684 271806
rect 292340 265298 292449 271806
rect 287660 258886 292449 265298
rect 297700 271730 302500 272310
rect 297700 265280 297852 271730
rect 301846 265280 302500 271730
rect 297700 258886 302500 265280
rect 350900 259010 355700 273678
rect 360951 259010 365740 273678
rect 609705 259990 609771 259993
rect 609705 259988 610549 259990
rect 609705 259932 609710 259988
rect 609766 259932 610549 259988
rect 609705 259930 610549 259932
rect 609705 259927 609771 259930
rect 384305 259738 384371 259741
rect 384489 259738 384555 259741
rect 516141 259738 516207 259741
rect 384305 259736 384555 259738
rect 384305 259680 384310 259736
rect 384366 259680 384494 259736
rect 384550 259680 384555 259736
rect 515388 259736 516207 259738
rect 384305 259678 384555 259680
rect 384305 259675 384371 259678
rect 384489 259675 384555 259678
rect 388370 259718 388436 259721
rect 392191 259718 392257 259721
rect 392631 259718 392697 259721
rect 393021 259718 393087 259721
rect 393870 259718 393936 259721
rect 395069 259718 395135 259721
rect 388370 259716 395135 259718
rect 384308 259612 384368 259675
rect 388370 259660 388375 259716
rect 388431 259660 392196 259716
rect 392252 259660 392636 259716
rect 392692 259660 393026 259716
rect 393082 259660 393875 259716
rect 393931 259660 395074 259716
rect 395130 259660 395135 259716
rect 388370 259658 395135 259660
rect 388370 259655 388436 259658
rect 383967 259592 384368 259612
rect 382618 259552 384368 259592
rect 382618 259532 384041 259552
rect 382618 259434 382684 259532
rect 389164 259446 389224 259658
rect 392191 259655 392257 259658
rect 392631 259655 392697 259658
rect 393021 259655 393087 259658
rect 393870 259655 393936 259658
rect 395069 259655 395135 259658
rect 414849 259718 414915 259721
rect 415419 259718 415485 259721
rect 417574 259718 417640 259721
rect 420967 259718 421033 259721
rect 424785 259718 424851 259721
rect 425243 259718 425309 259721
rect 425613 259718 425679 259721
rect 426441 259718 426507 259721
rect 414849 259716 415281 259718
rect 414849 259660 414854 259716
rect 414910 259660 415281 259716
rect 414849 259658 415281 259660
rect 414849 259655 414915 259658
rect 415221 259446 415281 259658
rect 415419 259716 426507 259718
rect 415419 259660 415424 259716
rect 415480 259660 417579 259716
rect 417635 259660 420972 259716
rect 421028 259660 424790 259716
rect 424846 259660 425248 259716
rect 425304 259660 425618 259716
rect 425674 259660 426446 259716
rect 426502 259660 426507 259716
rect 415419 259658 426507 259660
rect 415419 259655 415485 259658
rect 417574 259655 417640 259658
rect 420967 259655 421033 259658
rect 421764 259446 421824 259658
rect 424785 259655 424851 259658
rect 425243 259655 425309 259658
rect 425613 259655 425679 259658
rect 426441 259655 426507 259658
rect 446313 259718 446379 259721
rect 451005 259718 451071 259721
rect 480261 259718 480327 259721
rect 446313 259716 451071 259718
rect 446313 259660 446318 259716
rect 446374 259660 451010 259716
rect 451066 259660 451071 259716
rect 446313 259658 451071 259660
rect 446313 259655 446379 259658
rect 447621 259446 447681 259658
rect 451005 259655 451071 259658
rect 480221 259716 480327 259718
rect 480221 259660 480266 259716
rect 480322 259660 480327 259716
rect 480221 259655 480327 259660
rect 482574 259718 482640 259721
rect 485965 259718 486031 259721
rect 489783 259718 489849 259721
rect 490243 259718 490309 259721
rect 490611 259718 490677 259721
rect 491470 259718 491536 259721
rect 492679 259718 492745 259721
rect 494705 259718 494771 259721
rect 512829 259718 512895 259721
rect 515388 259718 516146 259736
rect 482574 259716 494771 259718
rect 482574 259660 482579 259716
rect 482635 259660 485970 259716
rect 486026 259660 489788 259716
rect 489844 259660 490248 259716
rect 490304 259660 490616 259716
rect 490672 259660 491475 259716
rect 491531 259660 492684 259716
rect 492740 259660 494710 259716
rect 494766 259660 494771 259716
rect 482574 259658 494771 259660
rect 512702 259716 516146 259718
rect 512702 259660 512834 259716
rect 512890 259680 516146 259716
rect 516202 259680 516207 259736
rect 512890 259678 516207 259680
rect 512890 259660 515465 259678
rect 516141 259675 516207 259678
rect 518533 259718 518599 259721
rect 522397 259718 522463 259721
rect 518533 259716 522463 259718
rect 512702 259658 515465 259660
rect 518533 259660 518538 259716
rect 518594 259660 522402 259716
rect 522458 259660 522463 259716
rect 518533 259658 522463 259660
rect 482574 259655 482640 259658
rect 485965 259655 486031 259658
rect 454409 259642 454475 259645
rect 454162 259640 454475 259642
rect 454162 259584 454414 259640
rect 454470 259584 454475 259640
rect 454162 259582 454475 259584
rect 454162 259446 454222 259582
rect 454409 259579 454475 259582
rect 480221 259446 480281 259655
rect 486761 259434 486827 259658
rect 489783 259655 489849 259658
rect 490243 259655 490309 259658
rect 490611 259655 490677 259658
rect 491470 259655 491536 259658
rect 492679 259655 492745 259658
rect 494705 259655 494771 259658
rect 512821 259655 512895 259658
rect 518533 259655 518599 259658
rect 512821 259446 512881 259655
rect 519361 259434 519427 259658
rect 522397 259655 522463 259658
rect 551170 259718 551236 259721
rect 554991 259718 555057 259721
rect 551170 259716 555057 259718
rect 551170 259660 551175 259716
rect 551231 259660 554996 259716
rect 555052 259660 555057 259716
rect 578057 259716 578123 259721
rect 578057 259691 578062 259716
rect 551170 259658 555057 259660
rect 551170 259655 551236 259658
rect 545029 259646 545095 259649
rect 545029 259644 545484 259646
rect 545029 259588 545034 259644
rect 545090 259588 545484 259644
rect 545029 259586 545484 259588
rect 545029 259583 545095 259586
rect 545418 259434 545484 259586
rect 551964 259446 552024 259658
rect 554991 259655 555057 259658
rect 578018 259660 578062 259691
rect 578118 259660 578123 259716
rect 578018 259655 578123 259660
rect 580817 259718 580883 259721
rect 583770 259718 583836 259721
rect 580817 259716 583836 259718
rect 580817 259660 580822 259716
rect 580878 259660 583775 259716
rect 583831 259660 583836 259716
rect 580817 259658 583836 259660
rect 580817 259655 580883 259658
rect 583770 259655 583836 259658
rect 584497 259718 584563 259721
rect 587579 259718 587645 259721
rect 588039 259718 588105 259721
rect 588421 259718 588487 259721
rect 590477 259718 590543 259721
rect 584497 259716 590543 259718
rect 584497 259660 584502 259716
rect 584558 259660 587584 259716
rect 587640 259660 588044 259716
rect 588100 259660 588426 259716
rect 588482 259660 590482 259716
rect 590538 259660 590543 259716
rect 584497 259658 590543 259660
rect 584497 259655 584624 259658
rect 587579 259655 587645 259658
rect 588039 259655 588105 259658
rect 588421 259655 588487 259658
rect 590477 259655 590543 259658
rect 578018 259622 578120 259655
rect 577597 259506 577663 259509
rect 577597 259504 577949 259506
rect 577597 259448 577602 259504
rect 577658 259448 577949 259504
rect 577597 259446 577949 259448
rect 577597 259443 577663 259446
rect 578018 259434 578084 259622
rect 584564 259446 584624 259655
rect 610489 259446 610549 259930
rect 610625 259854 610691 259857
rect 610621 259852 610691 259854
rect 610621 259796 610630 259852
rect 610686 259796 610691 259852
rect 610621 259791 610691 259796
rect 610621 259446 610681 259791
rect 615593 259718 615659 259721
rect 620193 259718 620259 259721
rect 621021 259718 621087 259721
rect 623079 259718 623145 259721
rect 625115 259718 625181 259721
rect 615593 259716 625181 259718
rect 615593 259660 615598 259716
rect 615654 259660 620198 259716
rect 620254 259660 621026 259716
rect 621082 259660 623084 259716
rect 623140 259660 625120 259716
rect 625176 259660 625181 259716
rect 615593 259658 625181 259660
rect 615593 259655 615659 259658
rect 617164 259446 617224 259658
rect 620193 259655 620259 259658
rect 621021 259655 621087 259658
rect 623079 259655 623145 259658
rect 625115 259655 625181 259658
rect 632521 259718 632587 259721
rect 651849 259718 651915 259721
rect 656395 259718 656461 259721
rect 660857 259718 660923 259721
rect 632521 259716 643281 259718
rect 632521 259660 632526 259716
rect 632582 259660 643281 259716
rect 632521 259658 643281 259660
rect 632521 259655 632587 259658
rect 640249 259582 640315 259585
rect 640249 259580 643149 259582
rect 640249 259524 640254 259580
rect 640310 259524 643149 259580
rect 640249 259522 643149 259524
rect 640249 259519 640315 259522
rect 643086 259462 643149 259522
rect 643089 259446 643149 259462
rect 643221 259446 643281 259658
rect 651849 259716 660923 259718
rect 651849 259660 651854 259716
rect 651910 259660 656400 259716
rect 656456 259660 660862 259716
rect 660918 259660 660923 259716
rect 651849 259658 660923 259660
rect 651849 259655 651915 259658
rect 656395 259655 656461 259658
rect 660857 259655 660923 259658
rect 649633 259614 649699 259619
rect 649633 259558 649638 259614
rect 649694 259609 649699 259614
rect 649694 259558 649827 259609
rect 649633 259553 649827 259558
rect 649636 259546 649827 259553
rect 649637 259543 649827 259546
rect 649761 259434 649827 259543
<< via3 >>
rect 210592 735934 215276 736476
rect 210598 732568 215282 733110
rect 272398 708222 276856 714638
rect 298404 718358 302880 724720
rect 308406 718386 312882 724748
rect 324690 718358 328652 724586
rect 335230 718386 339192 724614
rect 282478 708246 286936 714662
rect 252700 706184 252764 706248
rect 583517 729341 583581 729405
rect 583532 728720 583596 728784
rect 290420 699208 290484 699272
rect 252516 698800 252580 698864
rect 364572 694448 364636 694512
rect 382236 694448 382300 694512
rect 320780 688396 320844 688460
rect 320964 681800 321028 681864
rect 320780 675000 320844 675064
rect 321148 675000 321212 675064
rect 324036 669868 326786 670324
rect 359258 669812 362026 670284
rect 220076 667552 222120 667728
rect 290420 667248 290484 667312
rect 236536 665954 242984 667020
rect 320596 667112 320660 667176
rect 320964 667112 321028 667176
rect 364572 666976 364636 667040
rect 382236 666704 382300 666768
rect 251780 666024 251844 666088
rect 364572 664936 364636 665000
rect 215274 658184 216250 658662
rect 210476 656586 211618 657478
rect 619412 651880 619476 651944
rect 619044 651744 619108 651808
rect 620700 651608 620764 651672
rect 619228 651472 619292 651536
rect 619596 650792 619660 650856
rect 320596 650520 320660 650584
rect 252332 648480 252396 648544
rect 320780 648344 320844 648408
rect 252148 647392 252212 647456
rect 208172 647120 208236 647184
rect 251964 646984 252028 647048
rect 619412 644672 619476 644736
rect 619780 644400 619844 644464
rect 619228 637464 619292 637528
rect 619044 632432 619108 632496
rect 619044 632160 619108 632224
rect 619044 632024 619108 632088
rect 619044 628624 619108 628688
rect 619228 628352 619292 628416
rect 208172 628216 208236 628280
rect 619090 624468 619154 624472
rect 619090 624412 619094 624468
rect 619094 624412 619150 624468
rect 619150 624412 619154 624468
rect 619090 624408 619154 624412
rect 619412 621144 619476 621208
rect 619596 621144 619660 621208
rect 619228 620872 619292 620936
rect 619596 618288 619660 618352
rect 208172 612984 208236 613048
rect 619228 611624 619292 611688
rect 619228 610672 619292 610736
rect 208540 609176 208604 609240
rect 208172 606184 208236 606248
rect 208724 606184 208788 606248
rect 208172 605504 208236 605568
rect 619228 605368 619292 605432
rect 619228 603872 619292 603936
rect 208540 603328 208604 603392
rect 208356 600200 208420 600264
rect 208356 596452 208420 596456
rect 208356 596396 208406 596452
rect 208406 596396 208420 596452
rect 208356 596392 208420 596396
rect 619228 583744 619292 583808
rect 619044 583472 619108 583536
rect 619044 582928 619108 582992
rect 676084 581568 676148 581632
rect 676268 581432 676332 581496
rect 252148 578304 252212 578368
rect 619044 575856 619108 575920
rect 619044 575312 619108 575376
rect 676268 575040 676332 575104
rect 676084 573952 676148 574016
rect 619228 571912 619292 571976
rect 251964 564160 252028 564224
rect 208540 555592 208604 555656
rect 619228 551240 619292 551304
rect 208540 545392 208604 545456
rect 619412 541992 619476 542056
rect 619596 540496 619660 540560
rect 675900 536144 675964 536208
rect 676084 536008 676148 536072
rect 675900 534920 675964 534984
rect 675900 534104 675964 534168
rect 619412 533424 619476 533488
rect 676268 532472 676332 532536
rect 675900 531062 675964 531126
rect 675900 530024 675964 530088
rect 676268 524584 676332 524648
rect 676084 524040 676148 524104
rect 676268 486368 676332 486432
rect 676268 483719 676332 483783
rect 642378 454112 648850 458408
rect 642404 443982 648876 448278
rect 642392 414218 648886 418576
rect 642392 404262 648886 408620
rect 629506 374174 636022 378694
rect 236392 361160 242928 365470
rect 629506 364194 636022 368714
rect 619228 363152 619292 363216
rect 236506 351198 243042 355508
rect 215366 334842 222020 339360
rect 215346 324704 222000 329222
rect 620700 327792 620764 327856
rect 619412 306576 619476 306640
rect 251780 301952 251844 302016
rect 619044 299504 619108 299568
rect 228228 283116 228292 283180
rect 634944 280890 636264 281126
rect 642326 280712 643110 280916
rect 619412 280056 619476 280120
rect 228228 279920 228292 279984
rect 619228 279920 619292 279984
rect 252516 279784 252580 279848
rect 252700 279648 252764 279712
rect 252332 278968 252396 279032
rect 236380 273804 243110 276276
rect 288684 265298 292340 271806
rect 297852 265280 301846 271730
<< metal4 >>
rect 210544 735934 210592 736476
rect 215276 735934 215334 736476
rect 210562 732568 210598 733110
rect 215282 732568 215338 733110
rect 583516 729405 583582 729406
rect 583516 729341 583517 729405
rect 583581 729341 583582 729405
rect 583516 729340 583582 729341
rect 583519 729267 583579 729340
rect 583519 729202 583594 729267
rect 583534 728785 583594 729202
rect 583531 728784 583597 728785
rect 583531 728720 583532 728784
rect 583596 728720 583597 728784
rect 583531 728719 583597 728720
rect 236260 724588 243260 726448
rect 236260 718282 236496 724588
rect 242950 718282 243260 724588
rect 215178 714742 222178 716572
rect 215178 708210 215294 714742
rect 221958 708210 222178 714742
rect 215178 667728 222178 708210
rect 215178 667552 220076 667728
rect 222120 667552 222178 667728
rect 215178 658662 222178 667552
rect 215178 658184 215274 658662
rect 216250 658184 222178 658662
rect 210342 657478 211698 657548
rect 210342 656586 210476 657478
rect 211618 656586 211698 657478
rect 210342 656482 211698 656586
rect 208171 647184 208237 647185
rect 208171 647120 208172 647184
rect 208236 647120 208237 647184
rect 208171 647119 208237 647120
rect 208174 644570 208234 647119
rect 208174 644510 208418 644570
rect 208358 636842 208418 644510
rect 208174 636782 208418 636842
rect 208174 628281 208234 636782
rect 208171 628280 208237 628281
rect 208171 628216 208172 628280
rect 208236 628216 208237 628280
rect 208171 628215 208237 628216
rect 215178 621236 222178 658184
rect 215178 620726 215334 621236
rect 222024 620726 222178 621236
rect 208171 613048 208237 613049
rect 208171 612984 208172 613048
rect 208236 612984 208237 613048
rect 208171 612983 208237 612984
rect 208174 606249 208234 612983
rect 208539 609240 208605 609241
rect 208539 609176 208540 609240
rect 208604 609176 208605 609240
rect 208539 609175 208605 609176
rect 208171 606248 208237 606249
rect 208171 606184 208172 606248
rect 208236 606184 208237 606248
rect 208171 606183 208237 606184
rect 208171 605568 208237 605569
rect 208171 605504 208172 605568
rect 208236 605504 208237 605568
rect 208171 605503 208237 605504
rect 208174 598202 208234 605503
rect 208542 603393 208602 609175
rect 208723 606248 208789 606249
rect 208723 606184 208724 606248
rect 208788 606184 208789 606248
rect 208723 606183 208789 606184
rect 208539 603392 208605 603393
rect 208539 603328 208540 603392
rect 208604 603328 208605 603392
rect 208539 603327 208605 603328
rect 208726 601514 208786 606183
rect 208358 601454 208786 601514
rect 208358 600265 208418 601454
rect 208355 600264 208421 600265
rect 208355 600200 208356 600264
rect 208420 600200 208421 600264
rect 208355 600199 208421 600200
rect 208174 598142 208418 598202
rect 208358 596457 208418 598142
rect 208355 596456 208421 596457
rect 208355 596392 208356 596456
rect 208420 596392 208421 596456
rect 208355 596391 208421 596392
rect 215178 590600 222178 620726
rect 215178 590090 215334 590600
rect 222024 590090 222178 590600
rect 215178 559964 222178 590090
rect 215178 559454 215334 559964
rect 222024 559454 222178 559964
rect 208539 555656 208605 555657
rect 208539 555592 208540 555656
rect 208604 555592 208605 555656
rect 208539 555591 208605 555592
rect 208542 545457 208602 555591
rect 208539 545456 208605 545457
rect 208539 545392 208540 545456
rect 208604 545392 208605 545456
rect 208539 545391 208605 545392
rect 215178 529328 222178 559454
rect 215178 528818 215334 529328
rect 222024 528818 222178 529328
rect 215178 498692 222178 528818
rect 215178 498182 215334 498692
rect 222024 498182 222178 498692
rect 215178 468056 222178 498182
rect 215178 467546 215334 468056
rect 222024 467546 222178 468056
rect 215178 437420 222178 467546
rect 215178 436910 215334 437420
rect 222024 436910 222178 437420
rect 215178 406784 222178 436910
rect 215178 406274 215334 406784
rect 222024 406274 222178 406784
rect 215178 376148 222178 406274
rect 215178 375638 215334 376148
rect 222024 375638 222178 376148
rect 215178 345512 222178 375638
rect 215178 345002 215334 345512
rect 222024 345002 222178 345512
rect 215178 339360 222178 345002
rect 215178 334842 215366 339360
rect 222020 334842 222178 339360
rect 215178 329222 222178 334842
rect 215178 324704 215346 329222
rect 222000 324704 222178 329222
rect 215178 314876 222178 324704
rect 215178 314366 215334 314876
rect 222024 314366 222178 314876
rect 215178 284240 222178 314366
rect 215178 283730 215334 284240
rect 222024 283730 222178 284240
rect 215178 281764 222178 283730
rect 236260 667020 243260 718282
rect 298108 724748 339760 724882
rect 298108 724720 308406 724748
rect 298108 718358 298404 724720
rect 312882 724640 339760 724748
rect 312882 724586 328086 724640
rect 335662 724614 339760 724640
rect 302880 718386 308406 718412
rect 312882 718386 324690 724586
rect 302880 718358 324690 718386
rect 339192 718386 339760 724614
rect 298108 718332 328086 718358
rect 335662 718332 339760 718386
rect 298108 718196 339760 718332
rect 271852 714662 287358 714884
rect 271852 708272 272100 714662
rect 287134 708272 287358 714662
rect 271852 708222 272398 708272
rect 276856 708246 282478 708272
rect 286936 708246 287358 708272
rect 276856 708222 287358 708246
rect 271852 708048 287358 708222
rect 323992 714582 326872 715042
rect 323992 708230 324296 714582
rect 326628 708230 326872 714582
rect 252702 706249 252762 706270
rect 252699 706248 252765 706249
rect 252699 706184 252700 706248
rect 252764 706184 252765 706248
rect 252699 706183 252765 706184
rect 252515 698864 252581 698865
rect 252515 698800 252516 698864
rect 252580 698800 252581 698864
rect 252515 698799 252581 698800
rect 236260 665954 236536 667020
rect 242984 665954 243260 667020
rect 251779 666088 251845 666089
rect 251779 666024 251780 666088
rect 251844 666024 251845 666088
rect 251779 666023 251845 666024
rect 236260 657484 243260 665954
rect 236260 650864 236480 657484
rect 243016 650864 243260 657484
rect 236260 606090 243260 650864
rect 236260 605286 236480 606090
rect 243084 605286 243260 606090
rect 236260 575454 243260 605286
rect 236260 574650 236480 575454
rect 243084 574650 243260 575454
rect 236260 544818 243260 574650
rect 236260 544014 236480 544818
rect 243084 544014 243260 544818
rect 236260 514182 243260 544014
rect 236260 513378 236480 514182
rect 243084 513378 243260 514182
rect 236260 483546 243260 513378
rect 236260 482742 236480 483546
rect 243084 482742 243260 483546
rect 236260 452910 243260 482742
rect 236260 452106 236480 452910
rect 243084 452106 243260 452910
rect 236260 422274 243260 452106
rect 236260 421470 236480 422274
rect 243084 421470 243260 422274
rect 236260 391638 243260 421470
rect 236260 390834 236480 391638
rect 243084 390834 243260 391638
rect 236260 365470 243260 390834
rect 236260 361160 236392 365470
rect 242928 361160 243260 365470
rect 236260 361002 243260 361160
rect 236260 360198 236480 361002
rect 243084 360198 243260 361002
rect 236260 355508 243260 360198
rect 236260 351198 236506 355508
rect 243042 351198 243260 355508
rect 236260 330366 243260 351198
rect 236260 329562 236480 330366
rect 243084 329562 243260 330366
rect 236260 299730 243260 329562
rect 251782 302017 251842 666023
rect 252331 648544 252397 648545
rect 252331 648480 252332 648544
rect 252396 648480 252397 648544
rect 252331 648479 252397 648480
rect 252147 647456 252213 647457
rect 252147 647392 252148 647456
rect 252212 647392 252213 647456
rect 252147 647391 252213 647392
rect 251963 647048 252029 647049
rect 251963 646984 251964 647048
rect 252028 646984 252029 647048
rect 251963 646983 252029 646984
rect 251966 564225 252026 646983
rect 252150 578369 252210 647391
rect 252147 578368 252213 578369
rect 252147 578304 252148 578368
rect 252212 578304 252213 578368
rect 252147 578303 252213 578304
rect 251963 564224 252029 564225
rect 251963 564160 251964 564224
rect 252028 564160 252029 564224
rect 251963 564159 252029 564160
rect 251779 302016 251845 302017
rect 251779 301952 251780 302016
rect 251844 301952 251845 302016
rect 251779 301951 251845 301952
rect 236260 298926 236480 299730
rect 243084 298926 243260 299730
rect 236260 283224 243260 298926
rect 228227 283180 228293 283181
rect 228227 283116 228228 283180
rect 228292 283116 228293 283180
rect 228227 283115 228293 283116
rect 215178 281280 220364 281764
rect 221902 281280 222178 281764
rect 215178 271514 222178 281280
rect 228230 279985 228290 283115
rect 236260 282740 236796 283224
rect 238334 282740 243260 283224
rect 228227 279984 228293 279985
rect 228227 279920 228228 279984
rect 228292 279920 228293 279984
rect 228227 279919 228293 279920
rect 215178 265590 215702 271514
rect 221700 265590 222178 271514
rect 215178 264092 222178 265590
rect 236260 276276 243260 282740
rect 252334 279033 252394 648479
rect 252518 279849 252578 698799
rect 252515 279848 252581 279849
rect 252515 279784 252516 279848
rect 252580 279784 252581 279848
rect 252515 279783 252581 279784
rect 252702 279713 252762 706183
rect 281084 686494 283964 700450
rect 290419 699272 290485 699273
rect 290419 699208 290420 699272
rect 290484 699208 290485 699272
rect 290419 699207 290485 699208
rect 281084 685816 281194 686494
rect 283826 685816 283964 686494
rect 256047 645904 256367 657936
rect 271407 657592 271727 657936
rect 271244 650806 271254 657592
rect 271868 650806 271878 657592
rect 281084 657408 283964 685816
rect 290422 667313 290482 699207
rect 320779 688460 320845 688461
rect 320779 688396 320780 688460
rect 320844 688396 320845 688460
rect 320779 688395 320845 688396
rect 320782 675065 320842 688395
rect 320963 681864 321029 681865
rect 320963 681800 320964 681864
rect 321028 681800 321029 681864
rect 320963 681799 321029 681800
rect 320779 675064 320845 675065
rect 320779 675000 320780 675064
rect 320844 675000 320845 675064
rect 320779 674999 320845 675000
rect 320966 674790 321026 681799
rect 321147 675064 321213 675065
rect 321147 675000 321148 675064
rect 321212 675000 321213 675064
rect 321147 674999 321213 675000
rect 320782 674730 321026 674790
rect 290419 667312 290485 667313
rect 290419 667248 290420 667312
rect 290484 667248 290485 667312
rect 290419 667247 290485 667248
rect 320595 667176 320661 667177
rect 320595 667112 320596 667176
rect 320660 667112 320661 667176
rect 320595 667111 320661 667112
rect 281084 651056 281274 657408
rect 283606 651056 283964 657408
rect 271407 645904 271727 650806
rect 281084 650778 283964 651056
rect 286767 645904 287087 657936
rect 302127 657592 302447 657936
rect 301964 650806 301974 657592
rect 302588 650806 302598 657592
rect 302127 645904 302447 650806
rect 317487 645904 317807 657936
rect 320598 650585 320658 667111
rect 320595 650584 320661 650585
rect 320595 650520 320596 650584
rect 320660 650520 320661 650584
rect 320595 650519 320661 650520
rect 320782 648409 320842 674730
rect 321150 671066 321210 674999
rect 320966 671006 321210 671066
rect 323992 671124 326872 708230
rect 395620 714662 398500 715510
rect 395620 708310 395782 714662
rect 398114 708310 398500 714662
rect 320966 667177 321026 671006
rect 323992 670496 324082 671124
rect 326756 670496 326872 671124
rect 323992 670324 326872 670496
rect 323992 669868 324036 670324
rect 326786 669868 326872 670324
rect 320963 667176 321029 667177
rect 320963 667112 320964 667176
rect 321028 667112 321029 667176
rect 320963 667111 321029 667112
rect 323992 665370 326872 669868
rect 359204 686432 362084 700182
rect 364571 694512 364637 694513
rect 364571 694448 364572 694512
rect 364636 694448 364637 694512
rect 364571 694447 364637 694448
rect 382235 694512 382301 694513
rect 382235 694448 382236 694512
rect 382300 694448 382301 694512
rect 382235 694447 382301 694448
rect 359204 686356 362086 686432
rect 359204 685884 359270 686356
rect 361980 685884 362086 686356
rect 359204 685818 362086 685884
rect 359204 670284 362084 685818
rect 359204 669812 359258 670284
rect 362026 669812 362084 670284
rect 332847 657592 333167 657936
rect 332684 650806 332694 657592
rect 333308 650806 333318 657592
rect 320779 648408 320845 648409
rect 320779 648344 320780 648408
rect 320844 648344 320845 648408
rect 320779 648343 320845 648344
rect 332847 645904 333167 650806
rect 348207 645904 348527 657936
rect 359204 657328 362084 669812
rect 364574 667041 364634 694447
rect 364571 667040 364637 667041
rect 364571 666976 364572 667040
rect 364636 666976 364637 667040
rect 364571 666975 364637 666976
rect 364574 665001 364634 666975
rect 382238 666769 382298 694447
rect 395620 671074 398500 708310
rect 395620 670572 395734 671074
rect 398428 670572 398500 671074
rect 395620 669254 398500 670572
rect 629314 714720 636314 715798
rect 629314 708100 629592 714720
rect 636128 708100 636314 714720
rect 382235 666768 382301 666769
rect 382235 666704 382236 666768
rect 382300 666704 382301 666768
rect 382235 666703 382301 666704
rect 364571 665000 364637 665001
rect 364571 664936 364572 665000
rect 364636 664936 364637 665000
rect 364571 664935 364637 664936
rect 363567 657592 363887 657936
rect 359204 650976 359354 657328
rect 361686 650976 362084 657328
rect 359204 650510 362084 650976
rect 363404 650806 363414 657592
rect 364028 650806 364038 657592
rect 363567 645904 363887 650806
rect 378927 645904 379247 657936
rect 394287 657592 394607 657936
rect 394124 650806 394134 657592
rect 394748 650806 394758 657592
rect 394287 645904 394607 650806
rect 409647 645904 409967 657936
rect 425007 657592 425327 657936
rect 424844 650806 424854 657592
rect 425468 650806 425478 657592
rect 425007 645904 425327 650806
rect 440367 645904 440687 657936
rect 455727 657592 456047 657936
rect 455564 650806 455574 657592
rect 456188 650806 456198 657592
rect 455727 645904 456047 650806
rect 471087 645904 471407 657936
rect 486447 657592 486767 657936
rect 486284 650806 486294 657592
rect 486908 650806 486918 657592
rect 486447 645904 486767 650806
rect 501807 645904 502127 657936
rect 517167 657592 517487 657936
rect 517004 650806 517014 657592
rect 517628 650806 517638 657592
rect 517167 645904 517487 650806
rect 532527 645904 532847 657936
rect 547887 657592 548207 657936
rect 547724 650806 547734 657592
rect 548348 650806 548358 657592
rect 547887 645904 548207 650806
rect 563247 645904 563567 657936
rect 578607 657592 578927 657936
rect 578444 650806 578454 657592
rect 579068 650806 579078 657592
rect 578607 645904 578927 650806
rect 593967 645904 594287 657936
rect 609327 657592 609647 657936
rect 609164 650806 609174 657592
rect 609788 650806 609798 657592
rect 619411 651944 619477 651945
rect 619411 651880 619412 651944
rect 619476 651880 619477 651944
rect 619411 651879 619477 651880
rect 619043 651808 619109 651809
rect 619043 651744 619044 651808
rect 619108 651744 619109 651808
rect 619043 651743 619109 651744
rect 609327 645904 609647 650806
rect 619046 633038 619106 651743
rect 619227 651536 619293 651537
rect 619227 651472 619228 651536
rect 619292 651472 619293 651536
rect 619227 651471 619293 651472
rect 619230 637529 619290 651471
rect 619414 644737 619474 651879
rect 620699 651672 620765 651673
rect 620699 651608 620700 651672
rect 620764 651608 620765 651672
rect 620699 651607 620765 651608
rect 619595 650856 619661 650857
rect 619595 650792 619596 650856
rect 619660 650792 619661 650856
rect 619595 650791 619661 650792
rect 619411 644736 619477 644737
rect 619411 644672 619412 644736
rect 619476 644672 619477 644736
rect 619411 644671 619477 644672
rect 619598 644570 619658 650791
rect 619414 644510 619658 644570
rect 619227 637528 619293 637529
rect 619227 637464 619228 637528
rect 619292 637464 619293 637528
rect 619227 637463 619293 637464
rect 619414 637390 619474 644510
rect 619779 644464 619845 644465
rect 619779 644400 619780 644464
rect 619844 644400 619845 644464
rect 619779 644399 619845 644400
rect 619230 637330 619474 637390
rect 619230 636842 619290 637330
rect 619230 636782 619658 636842
rect 619046 632978 619290 633038
rect 619043 632496 619109 632497
rect 619043 632432 619044 632496
rect 619108 632432 619109 632496
rect 619043 632431 619109 632432
rect 619046 632225 619106 632431
rect 619043 632224 619109 632225
rect 619043 632160 619044 632224
rect 619108 632160 619109 632224
rect 619043 632159 619109 632160
rect 619043 632088 619109 632089
rect 619043 632024 619044 632088
rect 619108 632024 619109 632088
rect 619043 632023 619109 632024
rect 619046 628689 619106 632023
rect 619043 628688 619109 628689
rect 619043 628624 619044 628688
rect 619108 628624 619109 628688
rect 619043 628623 619109 628624
rect 619230 628550 619290 632978
rect 619598 629114 619658 636782
rect 619046 628490 619290 628550
rect 619414 629054 619658 629114
rect 619046 624473 619106 628490
rect 619227 628416 619293 628417
rect 619227 628352 619228 628416
rect 619292 628352 619293 628416
rect 619227 628351 619293 628352
rect 619046 624472 619155 624473
rect 619046 624410 619090 624472
rect 619089 624408 619090 624410
rect 619154 624408 619155 624472
rect 619089 624407 619155 624408
rect 619230 622430 619290 628351
rect 619046 622370 619290 622430
rect 619046 611550 619106 622370
rect 619414 621750 619474 629054
rect 619782 624698 619842 644399
rect 619230 621690 619474 621750
rect 619598 624638 619842 624698
rect 619230 621070 619290 621690
rect 619598 621386 619658 624638
rect 619414 621326 619658 621386
rect 619414 621209 619474 621326
rect 619411 621208 619477 621209
rect 619411 621144 619412 621208
rect 619476 621144 619477 621208
rect 619411 621143 619477 621144
rect 619595 621208 619661 621209
rect 619595 621144 619596 621208
rect 619660 621144 619661 621208
rect 619595 621143 619661 621144
rect 619230 621010 619474 621070
rect 619227 620936 619293 620937
rect 619227 620872 619228 620936
rect 619292 620872 619293 620936
rect 619227 620871 619293 620872
rect 619230 611689 619290 620871
rect 619227 611688 619293 611689
rect 619227 611624 619228 611688
rect 619292 611624 619293 611688
rect 619227 611623 619293 611624
rect 619046 611490 619290 611550
rect 619230 610870 619290 611490
rect 619046 610810 619290 610870
rect 619046 604750 619106 610810
rect 619227 610736 619293 610737
rect 619227 610672 619228 610736
rect 619292 610672 619293 610736
rect 619227 610671 619293 610672
rect 619230 605433 619290 610671
rect 619227 605432 619293 605433
rect 619227 605368 619228 605432
rect 619292 605368 619293 605432
rect 619227 605367 619293 605368
rect 619046 604690 619290 604750
rect 619230 604070 619290 604690
rect 619046 604010 619290 604070
rect 619046 583670 619106 604010
rect 619227 603936 619293 603937
rect 619227 603872 619228 603936
rect 619292 603872 619293 603936
rect 619227 603871 619293 603872
rect 619230 583809 619290 603871
rect 619227 583808 619293 583809
rect 619227 583744 619228 583808
rect 619292 583744 619293 583808
rect 619227 583743 619293 583744
rect 619046 583610 619290 583670
rect 619043 583536 619109 583537
rect 619043 583472 619044 583536
rect 619108 583472 619109 583536
rect 619043 583471 619109 583472
rect 619046 582993 619106 583471
rect 619043 582992 619109 582993
rect 619043 582928 619044 582992
rect 619108 582928 619109 582992
rect 619043 582927 619109 582928
rect 619230 578330 619290 583610
rect 619046 578270 619290 578330
rect 619046 576190 619106 578270
rect 619046 576130 619290 576190
rect 619043 575920 619109 575921
rect 619043 575856 619044 575920
rect 619108 575856 619109 575920
rect 619043 575855 619109 575856
rect 619046 575377 619106 575855
rect 619043 575376 619109 575377
rect 619043 575312 619044 575376
rect 619108 575312 619109 575376
rect 619043 575311 619109 575312
rect 619230 574150 619290 576130
rect 619046 574090 619290 574150
rect 619046 547418 619106 574090
rect 619227 571976 619293 571977
rect 619227 571912 619228 571976
rect 619292 571912 619293 571976
rect 619227 571911 619293 571912
rect 619230 551305 619290 571911
rect 619227 551304 619293 551305
rect 619227 551240 619228 551304
rect 619292 551240 619293 551304
rect 619227 551239 619293 551240
rect 619046 547358 619290 547418
rect 619230 377402 619290 547358
rect 619414 542190 619474 621010
rect 619598 618353 619658 621143
rect 619595 618352 619661 618353
rect 619595 618288 619596 618352
rect 619660 618288 619661 618352
rect 619595 618287 619661 618288
rect 619414 542130 619658 542190
rect 619411 542056 619477 542057
rect 619411 541992 619412 542056
rect 619476 541992 619477 542056
rect 619411 541991 619477 541992
rect 619414 533489 619474 541991
rect 619598 540561 619658 542130
rect 619595 540560 619661 540561
rect 619595 540496 619596 540560
rect 619660 540496 619661 540560
rect 619595 540495 619661 540496
rect 619411 533488 619477 533489
rect 619411 533424 619412 533488
rect 619476 533424 619477 533488
rect 619411 533423 619477 533424
rect 619046 377342 619290 377402
rect 619046 299569 619106 377342
rect 619227 363216 619293 363217
rect 619227 363152 619228 363216
rect 619292 363152 619293 363216
rect 619227 363151 619293 363152
rect 619043 299568 619109 299569
rect 619043 299504 619044 299568
rect 619108 299504 619109 299568
rect 619043 299503 619109 299504
rect 252699 279712 252765 279713
rect 252699 279648 252700 279712
rect 252764 279648 252765 279712
rect 252699 279647 252765 279648
rect 252331 279032 252397 279033
rect 252331 278968 252332 279032
rect 252396 278968 252397 279032
rect 252331 278967 252397 278968
rect 236260 273804 236380 276276
rect 243110 273804 243260 276276
rect 236260 263944 243260 273804
rect 256047 271840 256367 281104
rect 255796 271794 256490 271840
rect 255796 265110 255878 271794
rect 256414 265110 256490 271794
rect 255796 265018 256490 265110
rect 256047 264280 256367 265018
rect 271407 264280 271727 281104
rect 286767 271840 287087 281104
rect 286516 271794 287210 271840
rect 286516 265110 286598 271794
rect 287134 265110 287210 271794
rect 286516 265018 287210 265110
rect 288608 271806 302016 271880
rect 288608 265298 288684 271806
rect 292340 271730 302016 271806
rect 292340 271598 297852 271730
rect 292340 265298 297852 265318
rect 288608 265280 297852 265298
rect 301846 265280 302016 271730
rect 288608 265074 302016 265280
rect 286767 264280 287087 265018
rect 302127 264280 302447 281104
rect 317487 271840 317807 281104
rect 317236 271794 317930 271840
rect 317236 265110 317318 271794
rect 317854 265110 317930 271794
rect 317236 265018 317930 265110
rect 317487 264280 317807 265018
rect 332847 264280 333167 281104
rect 348207 271840 348527 281104
rect 347956 271794 348650 271840
rect 347956 265110 348038 271794
rect 348574 265110 348650 271794
rect 347956 265018 348650 265110
rect 348207 264280 348527 265018
rect 363567 264280 363887 281104
rect 378927 271840 379247 281104
rect 378676 271794 379370 271840
rect 378676 265110 378758 271794
rect 379294 265110 379370 271794
rect 378676 265018 379370 265110
rect 378927 264280 379247 265018
rect 394287 264280 394607 281104
rect 409647 271840 409967 281104
rect 409396 271794 410090 271840
rect 409396 265110 409478 271794
rect 410014 265110 410090 271794
rect 409396 265018 410090 265110
rect 409647 264280 409967 265018
rect 425007 264280 425327 281104
rect 440367 271840 440687 281104
rect 440116 271794 440810 271840
rect 440116 265110 440198 271794
rect 440734 265110 440810 271794
rect 440116 265018 440810 265110
rect 440367 264280 440687 265018
rect 455727 264280 456047 281104
rect 471087 271840 471407 281104
rect 470836 271794 471530 271840
rect 470836 265110 470918 271794
rect 471454 265110 471530 271794
rect 470836 265018 471530 265110
rect 471087 264280 471407 265018
rect 486447 264280 486767 281104
rect 501807 271840 502127 281104
rect 501656 271794 502350 271840
rect 501656 265110 501738 271794
rect 502274 265110 502350 271794
rect 501656 265018 502350 265110
rect 501807 264280 502127 265018
rect 517167 264280 517487 281104
rect 532527 271840 532847 281104
rect 532276 271794 532970 271840
rect 532276 265110 532358 271794
rect 532894 265110 532970 271794
rect 532276 265018 532970 265110
rect 532527 264280 532847 265018
rect 547887 264280 548207 281104
rect 563247 271840 563567 281104
rect 562996 271794 563690 271840
rect 562996 265110 563078 271794
rect 563614 265110 563690 271794
rect 562996 265018 563690 265110
rect 563247 264280 563567 265018
rect 578607 264280 578927 281104
rect 593967 271840 594287 281104
rect 593716 271794 594410 271840
rect 593716 265110 593798 271794
rect 594334 265110 594410 271794
rect 593716 265018 594410 265110
rect 593967 264280 594287 265018
rect 609327 264280 609647 281104
rect 619230 279985 619290 363151
rect 620702 327857 620762 651607
rect 629314 621302 636314 708100
rect 629314 620772 629388 621302
rect 636238 620772 636314 621302
rect 629314 590666 636314 620772
rect 629314 590136 629388 590666
rect 636238 590136 636314 590666
rect 629314 560030 636314 590136
rect 629314 559500 629388 560030
rect 636238 559500 636314 560030
rect 629314 529394 636314 559500
rect 629314 528864 629388 529394
rect 636238 528864 636314 529394
rect 629314 498758 636314 528864
rect 629314 498228 629388 498758
rect 636238 498228 636314 498758
rect 629314 468122 636314 498228
rect 629314 467592 629388 468122
rect 636238 467592 636314 468122
rect 629314 437486 636314 467592
rect 629314 436956 629388 437486
rect 636238 436956 636314 437486
rect 629314 406850 636314 436956
rect 629314 406320 629388 406850
rect 636238 406320 636314 406850
rect 629314 378694 636314 406320
rect 629314 376214 629506 378694
rect 636022 376214 636314 378694
rect 629314 375684 629388 376214
rect 636238 375684 636314 376214
rect 629314 374174 629506 375684
rect 636022 374174 636314 375684
rect 629314 368714 636314 374174
rect 629314 364194 629506 368714
rect 636022 364194 636314 368714
rect 629314 345578 636314 364194
rect 629314 345048 629388 345578
rect 636238 345048 636314 345578
rect 620699 327856 620765 327857
rect 620699 327792 620700 327856
rect 620764 327792 620765 327856
rect 620699 327791 620765 327792
rect 629314 314942 636314 345048
rect 629314 314412 629388 314942
rect 636238 314412 636314 314942
rect 619411 306640 619477 306641
rect 619411 306576 619412 306640
rect 619476 306576 619477 306640
rect 619411 306575 619477 306576
rect 619414 280121 619474 306575
rect 629314 284306 636314 314412
rect 629314 283776 629388 284306
rect 636238 283776 636314 284306
rect 629314 281126 636314 283776
rect 629314 280890 634944 281126
rect 636264 280890 636314 281126
rect 619411 280120 619477 280121
rect 619411 280056 619412 280120
rect 619476 280056 619477 280120
rect 619411 280055 619477 280056
rect 619227 279984 619293 279985
rect 619227 279920 619228 279984
rect 619292 279920 619293 279984
rect 619227 279919 619293 279920
rect 629314 271568 636314 280890
rect 642172 657556 649172 705258
rect 642172 650882 642350 657556
rect 648922 650882 649172 657556
rect 642172 636546 649172 650882
rect 642172 636112 642360 636546
rect 648994 636112 649172 636546
rect 642172 605910 649172 636112
rect 642172 605476 642360 605910
rect 648994 605476 649172 605910
rect 642172 575274 649172 605476
rect 676083 581632 676149 581633
rect 676083 581568 676084 581632
rect 676148 581568 676149 581632
rect 676083 581567 676149 581568
rect 642172 574840 642360 575274
rect 648994 574840 649172 575274
rect 642172 544638 649172 574840
rect 676086 574017 676146 581567
rect 676267 581496 676333 581497
rect 676267 581432 676268 581496
rect 676332 581432 676333 581496
rect 676267 581431 676333 581432
rect 676270 575105 676330 581431
rect 676267 575104 676333 575105
rect 676267 575040 676268 575104
rect 676332 575040 676333 575104
rect 676267 575039 676333 575040
rect 676083 574016 676149 574017
rect 676083 573952 676084 574016
rect 676148 573952 676149 574016
rect 676083 573951 676149 573952
rect 642172 544204 642360 544638
rect 648994 544204 649172 544638
rect 642172 514002 649172 544204
rect 675899 536208 675965 536209
rect 675899 536144 675900 536208
rect 675964 536144 675965 536208
rect 675899 536143 675965 536144
rect 675902 534985 675962 536143
rect 676083 536072 676149 536073
rect 676083 536008 676084 536072
rect 676148 536008 676149 536072
rect 676083 536007 676149 536008
rect 675899 534984 675965 534985
rect 675899 534920 675900 534984
rect 675964 534920 675965 534984
rect 675899 534919 675965 534920
rect 675902 534169 675962 534919
rect 675899 534168 675965 534169
rect 675899 534104 675900 534168
rect 675964 534104 675965 534168
rect 675899 534103 675965 534104
rect 675902 531127 675962 534103
rect 675899 531126 675965 531127
rect 675899 531062 675900 531126
rect 675964 531062 675965 531126
rect 675899 531061 675965 531062
rect 675902 530089 675962 531061
rect 675899 530088 675965 530089
rect 675899 530024 675900 530088
rect 675964 530024 675965 530088
rect 675899 530023 675965 530024
rect 676086 524105 676146 536007
rect 676267 532536 676333 532537
rect 676267 532472 676268 532536
rect 676332 532472 676333 532536
rect 676267 532471 676333 532472
rect 676270 524649 676330 532471
rect 676267 524648 676333 524649
rect 676267 524584 676268 524648
rect 676332 524584 676333 524648
rect 676267 524583 676333 524584
rect 676083 524104 676149 524105
rect 676083 524040 676084 524104
rect 676148 524040 676149 524104
rect 676083 524039 676149 524040
rect 642172 513568 642360 514002
rect 648994 513568 649172 514002
rect 642172 483366 649172 513568
rect 676267 486432 676333 486433
rect 676267 486368 676268 486432
rect 676332 486368 676333 486432
rect 676267 486367 676333 486368
rect 676270 483784 676330 486367
rect 676267 483783 676333 483784
rect 676267 483719 676268 483783
rect 676332 483719 676333 483783
rect 676267 483718 676333 483719
rect 642172 482932 642360 483366
rect 648994 482932 649172 483366
rect 642172 458408 649172 482932
rect 642172 454112 642378 458408
rect 648850 454112 649172 458408
rect 642172 452730 649172 454112
rect 642172 452296 642360 452730
rect 648994 452296 649172 452730
rect 642172 448278 649172 452296
rect 642172 443982 642404 448278
rect 648876 443982 649172 448278
rect 642172 422094 649172 443982
rect 642172 421660 642360 422094
rect 648994 421660 649172 422094
rect 642172 418576 649172 421660
rect 642172 414218 642392 418576
rect 648886 414218 649172 418576
rect 642172 408620 649172 414218
rect 642172 404262 642392 408620
rect 648886 404262 649172 408620
rect 642172 391458 649172 404262
rect 642172 391024 642360 391458
rect 648994 391024 649172 391458
rect 642172 360822 649172 391024
rect 642172 360388 642360 360822
rect 648994 360388 649172 360822
rect 642172 330186 649172 360388
rect 642172 329752 642360 330186
rect 648994 329752 649172 330186
rect 642172 299550 649172 329752
rect 642172 299116 642360 299550
rect 648994 299116 649172 299550
rect 642172 280916 649172 299116
rect 642172 280712 642326 280916
rect 643110 280712 649172 280916
rect 642172 276316 649172 280712
rect 629314 265302 629662 271568
rect 635970 265302 636314 271568
rect 629314 264404 636314 265302
<< via4 >>
rect 236496 718282 242950 724588
rect 215294 708210 221958 714742
rect 210476 656586 211618 657478
rect 215334 620726 222024 621236
rect 215334 590090 222024 590600
rect 215334 559454 222024 559964
rect 215334 528818 222024 529328
rect 215334 498182 222024 498692
rect 215334 467546 222024 468056
rect 215334 436910 222024 437420
rect 215334 406274 222024 406784
rect 215334 375638 222024 376148
rect 215334 345002 222024 345512
rect 215334 314366 222024 314876
rect 215334 283730 222024 284240
rect 301344 718412 302880 724720
rect 302880 718412 308406 724720
rect 308406 718412 308920 724720
rect 328086 724614 335662 724640
rect 328086 724586 335230 724614
rect 328086 718358 328652 724586
rect 328652 718386 335230 724586
rect 335230 718386 335662 724614
rect 328652 718358 335662 718386
rect 328086 718332 335662 718358
rect 272100 714638 282478 714662
rect 272100 708272 272398 714638
rect 272398 708272 276856 714638
rect 276856 708272 282478 714638
rect 282478 708272 286936 714662
rect 286936 708272 287134 714662
rect 324296 708230 326628 714582
rect 236480 650864 243016 657484
rect 236480 605286 243084 606090
rect 236480 574650 243084 575454
rect 236480 544014 243084 544818
rect 236480 513378 243084 514182
rect 236480 482742 243084 483546
rect 236480 452106 243084 452910
rect 236480 421470 243084 422274
rect 236480 390834 243084 391638
rect 236480 360198 243084 361002
rect 236480 329562 243084 330366
rect 236480 298926 243084 299730
rect 220364 281280 221902 281764
rect 236796 282740 238334 283224
rect 215702 265590 221700 271514
rect 281194 685816 283826 686494
rect 271254 650806 271868 657592
rect 281274 651056 283606 657408
rect 301974 650806 302588 657592
rect 395782 708310 398114 714662
rect 324082 670496 326756 671124
rect 359270 685884 361980 686356
rect 332694 650806 333308 657592
rect 395734 670572 398428 671074
rect 629592 708100 636128 714720
rect 359354 650976 361686 657328
rect 363414 650806 364028 657592
rect 394134 650806 394748 657592
rect 424854 650806 425468 657592
rect 455574 650806 456188 657592
rect 486294 650806 486908 657592
rect 517014 650806 517628 657592
rect 547734 650806 548348 657592
rect 578454 650806 579068 657592
rect 609174 650806 609788 657592
rect 255878 265110 256414 271794
rect 286598 265110 287134 271794
rect 289058 265318 292340 271598
rect 292340 265318 297852 271598
rect 297852 265318 301660 271598
rect 317318 265110 317854 271794
rect 348038 265110 348574 271794
rect 378758 265110 379294 271794
rect 409478 265110 410014 271794
rect 440198 265110 440734 271794
rect 470918 265110 471454 271794
rect 501738 265110 502274 271794
rect 532358 265110 532894 271794
rect 563078 265110 563614 271794
rect 593798 265110 594334 271794
rect 629388 620772 636238 621302
rect 629388 590136 636238 590666
rect 629388 559500 636238 560030
rect 629388 528864 636238 529394
rect 629388 498228 636238 498758
rect 629388 467592 636238 468122
rect 629388 436956 636238 437486
rect 629388 406320 636238 406850
rect 629388 375684 629506 376214
rect 629506 375684 636022 376214
rect 636022 375684 636238 376214
rect 629388 345048 636238 345578
rect 629388 314412 636238 314942
rect 629388 283776 636238 284306
rect 642350 650882 648922 657556
rect 642360 636112 648994 636546
rect 642360 605476 648994 605910
rect 642360 574840 648994 575274
rect 642360 544204 648994 544638
rect 642360 513568 648994 514002
rect 642360 482932 648994 483366
rect 642360 452296 648994 452730
rect 642360 421660 648994 422094
rect 642360 391024 648994 391458
rect 642360 360388 648994 360822
rect 642360 329752 648994 330186
rect 642360 299116 648994 299550
rect 629662 265302 635970 271568
<< metal5 >>
rect 209798 730450 215828 731626
rect 235552 724720 341316 725034
rect 235552 724588 301344 724720
rect 235552 718282 236496 724588
rect 242950 718412 301344 724588
rect 308920 724640 341316 724720
rect 308920 718412 328086 724640
rect 242950 718332 328086 718412
rect 335662 718332 341316 724640
rect 242950 718282 341316 718332
rect 235552 718034 341316 718282
rect 214554 714742 656140 714960
rect 214554 708210 215294 714742
rect 221958 714720 656140 714742
rect 221958 714662 629592 714720
rect 221958 708272 272100 714662
rect 287134 714582 395782 714662
rect 287134 708272 324296 714582
rect 221958 708230 324296 708272
rect 326628 708310 395782 714582
rect 398114 708310 629592 714662
rect 326628 708230 629592 708310
rect 221958 708210 629592 708230
rect 214554 708100 629592 708210
rect 636128 708100 656140 714720
rect 214554 707960 656140 708100
rect 281094 686494 283948 686572
rect 281094 686293 281194 686494
rect 281066 685973 281194 686293
rect 281094 685816 281194 685973
rect 283826 686293 283948 686494
rect 359212 686356 362086 686432
rect 283826 685973 289570 686293
rect 283826 685816 283948 685973
rect 359212 685884 359270 686356
rect 361980 686293 362086 686356
rect 361980 685973 363322 686293
rect 361980 685884 362086 685973
rect 359212 685818 362086 685884
rect 281094 685728 283948 685816
rect 324004 671124 326844 671190
rect 324004 670975 324082 671124
rect 320188 670655 324082 670975
rect 324004 670496 324082 670655
rect 326756 670975 326844 671124
rect 395638 671074 398514 671132
rect 395638 670975 395734 671074
rect 326756 670655 326876 670975
rect 389994 670655 395734 670975
rect 326756 670496 326844 670655
rect 324004 670446 326844 670496
rect 395638 670572 395734 670655
rect 398428 670572 398514 671074
rect 395638 670486 398514 670572
rect 210232 657592 654534 657716
rect 210232 657484 271254 657592
rect 210232 657478 236480 657484
rect 210232 656586 210476 657478
rect 211618 656586 236480 657478
rect 210232 650864 236480 656586
rect 243016 650864 271254 657484
rect 210232 650806 271254 650864
rect 271868 657408 301974 657592
rect 271868 651056 281274 657408
rect 283606 651056 301974 657408
rect 271868 650806 301974 651056
rect 302588 650806 332694 657592
rect 333308 657328 363414 657592
rect 333308 650976 359354 657328
rect 361686 650976 363414 657328
rect 333308 650806 363414 650976
rect 364028 650806 394134 657592
rect 394748 650806 424854 657592
rect 425468 650806 455574 657592
rect 456188 650806 486294 657592
rect 486908 650806 517014 657592
rect 517628 650806 547734 657592
rect 548348 650806 578454 657592
rect 579068 650806 609174 657592
rect 609788 657556 654534 657592
rect 609788 650882 642350 657556
rect 648922 650882 654534 657556
rect 609788 650806 654534 650882
rect 210232 650716 654534 650806
rect 642242 636546 649094 636638
rect 642242 636504 642360 636546
rect 618438 636184 642360 636504
rect 642242 636112 642360 636184
rect 648994 636504 649094 636546
rect 648994 636184 649574 636504
rect 648994 636112 649094 636184
rect 642242 636008 649094 636112
rect 215266 621236 222110 621304
rect 215266 621186 215334 621236
rect 214996 620866 215334 621186
rect 215266 620726 215334 620866
rect 222024 621186 222110 621236
rect 629304 621302 636306 621374
rect 629304 621186 629388 621302
rect 222024 620866 253382 621186
rect 618438 620866 629388 621186
rect 222024 620726 222110 620866
rect 215266 620650 222110 620726
rect 629304 620772 629388 620866
rect 636238 621186 636306 621302
rect 636238 620866 636706 621186
rect 636238 620772 636306 620866
rect 629304 620690 636306 620772
rect 236328 606090 243170 606176
rect 236328 605868 236480 606090
rect 236204 605548 236480 605868
rect 236328 605286 236480 605548
rect 243084 605868 243170 606090
rect 642242 605910 649094 606002
rect 642242 605868 642360 605910
rect 243084 605548 253382 605868
rect 618438 605548 642360 605868
rect 243084 605286 243170 605548
rect 642242 605476 642360 605548
rect 648994 605868 649094 605910
rect 648994 605548 649588 605868
rect 648994 605476 649094 605548
rect 642242 605372 649094 605476
rect 236328 605200 243170 605286
rect 215266 590600 222110 590668
rect 215266 590550 215334 590600
rect 214466 590230 215334 590550
rect 215266 590090 215334 590230
rect 222024 590550 222110 590600
rect 629304 590666 636306 590738
rect 629304 590550 629388 590666
rect 222024 590230 253382 590550
rect 618438 590230 629388 590550
rect 222024 590090 222110 590230
rect 215266 590014 222110 590090
rect 629304 590136 629388 590230
rect 636238 590550 636306 590666
rect 636238 590230 636706 590550
rect 636238 590136 636306 590230
rect 629304 590054 636306 590136
rect 236328 575454 243170 575540
rect 236328 575232 236480 575454
rect 236204 574912 236480 575232
rect 236328 574650 236480 574912
rect 243084 575232 243170 575454
rect 642242 575274 649094 575366
rect 642242 575232 642360 575274
rect 243084 574912 253382 575232
rect 618438 574912 642360 575232
rect 243084 574650 243170 574912
rect 642242 574840 642360 574912
rect 648994 575232 649094 575274
rect 648994 574912 649588 575232
rect 648994 574840 649094 574912
rect 642242 574736 649094 574840
rect 236328 574564 243170 574650
rect 215266 559964 222110 560032
rect 215266 559914 215334 559964
rect 214728 559594 215334 559914
rect 215266 559454 215334 559594
rect 222024 559914 222110 559964
rect 629304 560030 636306 560102
rect 629304 559914 629388 560030
rect 222024 559594 253382 559914
rect 618438 559594 629388 559914
rect 222024 559454 222110 559594
rect 215266 559378 222110 559454
rect 629304 559500 629388 559594
rect 636238 559914 636306 560030
rect 636238 559594 636706 559914
rect 636238 559500 636306 559594
rect 629304 559418 636306 559500
rect 236328 544818 243170 544904
rect 236328 544596 236480 544818
rect 236204 544276 236480 544596
rect 236328 544014 236480 544276
rect 243084 544596 243170 544818
rect 642242 544638 649094 544730
rect 642242 544596 642360 544638
rect 243084 544276 253382 544596
rect 618438 544276 642360 544596
rect 243084 544014 243170 544276
rect 642242 544204 642360 544276
rect 648994 544596 649094 544638
rect 648994 544276 649588 544596
rect 648994 544204 649094 544276
rect 642242 544100 649094 544204
rect 236328 543928 243170 544014
rect 215266 529328 222110 529396
rect 215266 529278 215334 529328
rect 214466 528958 215334 529278
rect 215266 528818 215334 528958
rect 222024 529278 222110 529328
rect 629304 529394 636306 529466
rect 629304 529278 629388 529394
rect 222024 528958 253382 529278
rect 618438 528958 629388 529278
rect 222024 528818 222110 528958
rect 215266 528742 222110 528818
rect 629304 528864 629388 528958
rect 636238 529278 636306 529394
rect 636238 528958 636706 529278
rect 636238 528864 636306 528958
rect 629304 528782 636306 528864
rect 236328 514182 243170 514268
rect 236328 513960 236480 514182
rect 236204 513640 236480 513960
rect 236328 513378 236480 513640
rect 243084 513960 243170 514182
rect 642242 514002 649094 514094
rect 642242 513960 642360 514002
rect 243084 513640 253382 513960
rect 618438 513640 642360 513960
rect 243084 513378 243170 513640
rect 642242 513568 642360 513640
rect 648994 513960 649094 514002
rect 648994 513640 649720 513960
rect 648994 513568 649094 513640
rect 642242 513464 649094 513568
rect 236328 513292 243170 513378
rect 215266 498692 222110 498760
rect 215266 498642 215334 498692
rect 214596 498322 215334 498642
rect 215266 498182 215334 498322
rect 222024 498642 222110 498692
rect 629304 498758 636306 498830
rect 629304 498642 629388 498758
rect 222024 498322 253382 498642
rect 618438 498322 629388 498642
rect 222024 498182 222110 498322
rect 215266 498106 222110 498182
rect 629304 498228 629388 498322
rect 636238 498642 636306 498758
rect 636238 498322 636706 498642
rect 636238 498228 636306 498322
rect 629304 498146 636306 498228
rect 236328 483546 243170 483632
rect 236328 483324 236480 483546
rect 236204 483004 236480 483324
rect 236328 482742 236480 483004
rect 243084 483324 243170 483546
rect 642242 483366 649094 483458
rect 642242 483324 642360 483366
rect 243084 483004 253382 483324
rect 618438 483004 642360 483324
rect 243084 482742 243170 483004
rect 642242 482932 642360 483004
rect 648994 483324 649094 483366
rect 648994 483004 649720 483324
rect 648994 482932 649094 483004
rect 642242 482828 649094 482932
rect 236328 482656 243170 482742
rect 215266 468056 222110 468124
rect 215266 468006 215334 468056
rect 214596 467686 215334 468006
rect 215266 467546 215334 467686
rect 222024 468006 222110 468056
rect 629304 468122 636306 468194
rect 629304 468006 629388 468122
rect 222024 467686 253382 468006
rect 618438 467686 629388 468006
rect 222024 467546 222110 467686
rect 215266 467470 222110 467546
rect 629304 467592 629388 467686
rect 636238 468006 636306 468122
rect 636238 467686 636706 468006
rect 636238 467592 636306 467686
rect 629304 467510 636306 467592
rect 236328 452910 243170 452996
rect 236328 452688 236480 452910
rect 236204 452368 236480 452688
rect 236328 452106 236480 452368
rect 243084 452688 243170 452910
rect 642242 452730 649094 452822
rect 642242 452688 642360 452730
rect 243084 452368 253382 452688
rect 618438 452368 642360 452688
rect 243084 452106 243170 452368
rect 642242 452296 642360 452368
rect 648994 452688 649094 452730
rect 648994 452368 649720 452688
rect 648994 452296 649094 452368
rect 642242 452192 649094 452296
rect 236328 452020 243170 452106
rect 215266 437420 222110 437488
rect 215266 437370 215334 437420
rect 214728 437050 215334 437370
rect 215266 436910 215334 437050
rect 222024 437370 222110 437420
rect 629304 437486 636306 437558
rect 629304 437370 629388 437486
rect 222024 437050 253382 437370
rect 618438 437050 629388 437370
rect 222024 436910 222110 437050
rect 215266 436834 222110 436910
rect 629304 436956 629388 437050
rect 636238 437370 636306 437486
rect 636238 437050 636706 437370
rect 636238 436956 636306 437050
rect 629304 436874 636306 436956
rect 236328 422274 243170 422360
rect 236328 422052 236480 422274
rect 236204 421732 236480 422052
rect 236328 421470 236480 421732
rect 243084 422052 243170 422274
rect 642242 422094 649094 422186
rect 642242 422052 642360 422094
rect 243084 421732 253382 422052
rect 618438 421732 642360 422052
rect 243084 421470 243170 421732
rect 642242 421660 642360 421732
rect 648994 422052 649094 422094
rect 648994 421732 649720 422052
rect 648994 421660 649094 421732
rect 642242 421556 649094 421660
rect 236328 421384 243170 421470
rect 215266 406784 222110 406852
rect 215266 406734 215334 406784
rect 214596 406414 215334 406734
rect 215266 406274 215334 406414
rect 222024 406734 222110 406784
rect 629304 406850 636306 406922
rect 629304 406734 629388 406850
rect 222024 406414 253382 406734
rect 618438 406414 629388 406734
rect 222024 406274 222110 406414
rect 215266 406198 222110 406274
rect 629304 406320 629388 406414
rect 636238 406734 636306 406850
rect 636238 406414 636706 406734
rect 636238 406320 636306 406414
rect 629304 406238 636306 406320
rect 236328 391638 243170 391724
rect 236328 391416 236480 391638
rect 236204 391096 236480 391416
rect 236328 390834 236480 391096
rect 243084 391416 243170 391638
rect 642242 391458 649094 391550
rect 642242 391416 642360 391458
rect 243084 391096 253382 391416
rect 618438 391096 642360 391416
rect 243084 390834 243170 391096
rect 642242 391024 642360 391096
rect 648994 391416 649094 391458
rect 648994 391096 649588 391416
rect 648994 391024 649094 391096
rect 642242 390920 649094 391024
rect 236328 390748 243170 390834
rect 215266 376148 222110 376216
rect 215266 376098 215334 376148
rect 214596 375778 215334 376098
rect 215266 375638 215334 375778
rect 222024 376098 222110 376148
rect 629304 376214 636306 376286
rect 629304 376098 629388 376214
rect 222024 375778 253382 376098
rect 618438 375778 629388 376098
rect 222024 375638 222110 375778
rect 215266 375562 222110 375638
rect 629304 375684 629388 375778
rect 636238 376098 636306 376214
rect 636238 375778 636706 376098
rect 636238 375684 636306 375778
rect 629304 375602 636306 375684
rect 236328 361002 243170 361088
rect 236328 360780 236480 361002
rect 236204 360460 236480 360780
rect 236328 360198 236480 360460
rect 243084 360780 243170 361002
rect 642242 360822 649094 360914
rect 642242 360780 642360 360822
rect 243084 360460 253382 360780
rect 618438 360460 642360 360780
rect 243084 360198 243170 360460
rect 642242 360388 642360 360460
rect 648994 360780 649094 360822
rect 648994 360460 649328 360780
rect 648994 360388 649094 360460
rect 642242 360284 649094 360388
rect 236328 360112 243170 360198
rect 215266 345512 222110 345580
rect 215266 345462 215334 345512
rect 214728 345142 215334 345462
rect 215266 345002 215334 345142
rect 222024 345462 222110 345512
rect 629304 345578 636306 345650
rect 629304 345462 629388 345578
rect 222024 345142 253382 345462
rect 618438 345142 629388 345462
rect 222024 345002 222110 345142
rect 215266 344926 222110 345002
rect 629304 345048 629388 345142
rect 636238 345462 636306 345578
rect 636238 345142 636706 345462
rect 636238 345048 636306 345142
rect 629304 344966 636306 345048
rect 236328 330366 243170 330452
rect 236328 330144 236480 330366
rect 236204 329824 236480 330144
rect 236328 329562 236480 329824
rect 243084 330144 243170 330366
rect 642242 330186 649094 330278
rect 642242 330144 642360 330186
rect 243084 329824 253382 330144
rect 618438 329824 642360 330144
rect 243084 329562 243170 329824
rect 642242 329752 642360 329824
rect 648994 330144 649094 330186
rect 648994 329824 649146 330144
rect 648994 329752 649094 329824
rect 642242 329648 649094 329752
rect 236328 329476 243170 329562
rect 215266 314876 222110 314944
rect 215266 314826 215334 314876
rect 214596 314506 215334 314826
rect 215266 314366 215334 314506
rect 222024 314826 222110 314876
rect 629304 314942 636306 315014
rect 629304 314826 629388 314942
rect 222024 314506 253382 314826
rect 618438 314506 629388 314826
rect 222024 314366 222110 314506
rect 215266 314290 222110 314366
rect 629304 314412 629388 314506
rect 636238 314826 636306 314942
rect 636238 314506 636706 314826
rect 636238 314412 636306 314506
rect 629304 314330 636306 314412
rect 236328 299730 243170 299816
rect 236328 299508 236480 299730
rect 236204 299188 236480 299508
rect 236328 298926 236480 299188
rect 243084 299508 243170 299730
rect 642242 299550 649094 299642
rect 642242 299508 642360 299550
rect 243084 299188 253382 299508
rect 618438 299188 642360 299508
rect 243084 298926 243170 299188
rect 642242 299116 642360 299188
rect 648994 299508 649094 299550
rect 648994 299188 649588 299508
rect 648994 299116 649094 299188
rect 642242 299012 649094 299116
rect 236328 298840 243170 298926
rect 215266 284240 222110 284308
rect 215266 284190 215334 284240
rect 214596 283870 215334 284190
rect 215266 283730 215334 283870
rect 222024 284190 222110 284240
rect 629304 284306 636306 284378
rect 629304 284190 629388 284306
rect 222024 283870 253382 284190
rect 618438 283870 629388 284190
rect 222024 283730 222110 283870
rect 215266 283654 222110 283730
rect 629304 283776 629388 283870
rect 636238 284190 636306 284306
rect 636238 283870 636706 284190
rect 636238 283776 636306 283870
rect 629304 283694 636306 283776
rect 236688 283224 238436 283278
rect 236688 283160 236796 283224
rect 232080 282840 236796 283160
rect 236688 282740 236796 282840
rect 238334 283160 238436 283224
rect 238334 282840 238440 283160
rect 238334 282740 238436 282840
rect 236688 282666 238436 282740
rect 220234 281764 222052 281824
rect 220234 281280 220364 281764
rect 221902 281660 222052 281764
rect 221902 281340 228400 281660
rect 221902 281280 222052 281340
rect 220234 281210 222052 281280
rect 212802 271794 655872 271942
rect 212802 271514 255878 271794
rect 212802 265590 215702 271514
rect 221700 265590 255878 271514
rect 212802 265110 255878 265590
rect 256414 265110 286598 271794
rect 287134 271598 317318 271794
rect 287134 265318 289058 271598
rect 301660 265318 317318 271598
rect 287134 265110 317318 265318
rect 317854 265110 348038 271794
rect 348574 265110 378758 271794
rect 379294 265110 409478 271794
rect 410014 265110 440198 271794
rect 440734 265110 470918 271794
rect 471454 265110 501738 271794
rect 502274 265110 532358 271794
rect 532894 265110 563078 271794
rect 563614 265110 593798 271794
rect 594334 271568 655872 271794
rect 594334 265302 629662 271568
rect 635970 265302 655872 271568
rect 594334 265110 655872 265302
rect 212802 264942 655872 265110
use sky130_ef_io__corner_pad  corner[1] /usr/share/pdk/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1587416550
transform -1 0 208000 0 -1 260300
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_1um  FILLER_1025 /usr/share/pdk/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1587416550
transform -1 0 208200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1026
timestamp 1587416550
transform -1 0 208400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1027
timestamp 1587416550
transform -1 0 208600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1028
timestamp 1587416550
transform -1 0 208800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1029
timestamp 1587416550
transform -1 0 209000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1030
timestamp 1587416550
transform -1 0 209200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1031
timestamp 1587416550
transform -1 0 209400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1032
timestamp 1587416550
transform -1 0 209600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1033
timestamp 1587416550
transform -1 0 209800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1034
timestamp 1587416550
transform -1 0 210000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1035
timestamp 1587416550
transform -1 0 210200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1036
timestamp 1587416550
transform -1 0 210400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1037
timestamp 1587416550
transform -1 0 210600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1038
timestamp 1587416550
transform -1 0 210800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1039
timestamp 1587416550
transform -1 0 211000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1040
timestamp 1587416550
transform -1 0 211200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1041
timestamp 1587416550
transform -1 0 211400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1042
timestamp 1587416550
transform -1 0 211600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1043
timestamp 1587416550
transform -1 0 211800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1044
timestamp 1587416550
transform -1 0 212000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1045
timestamp 1587416550
transform -1 0 212200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1046
timestamp 1587416550
transform -1 0 212400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1047
timestamp 1587416550
transform -1 0 212600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1048
timestamp 1587416550
transform -1 0 212800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1049
timestamp 1587416550
transform -1 0 213000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1050
timestamp 1587416550
transform -1 0 213200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1051
timestamp 1587416550
transform -1 0 213400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1052
timestamp 1587416550
transform -1 0 213600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1053
timestamp 1587416550
transform -1 0 213800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1054
timestamp 1587416550
transform -1 0 214000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1055
timestamp 1587416550
transform -1 0 214200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1056
timestamp 1587416550
transform -1 0 214400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1057
timestamp 1587416550
transform -1 0 214600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1058
timestamp 1587416550
transform -1 0 214800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1059
timestamp 1587416550
transform -1 0 215000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1060
timestamp 1587416550
transform -1 0 215200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1061
timestamp 1587416550
transform -1 0 215400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1062
timestamp 1587416550
transform -1 0 215600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1063
timestamp 1587416550
transform -1 0 215800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1064
timestamp 1587416550
transform -1 0 216000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1065
timestamp 1587416550
transform -1 0 216200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1066
timestamp 1587416550
transform -1 0 216400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1067
timestamp 1587416550
transform -1 0 216600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1068
timestamp 1587416550
transform -1 0 216800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1069
timestamp 1587416550
transform -1 0 217000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1070
timestamp 1587416550
transform -1 0 217200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1071
timestamp 1587416550
transform -1 0 217400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1072
timestamp 1587416550
transform -1 0 217600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1073
timestamp 1587416550
transform -1 0 217800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1074
timestamp 1587416550
transform -1 0 218000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1075
timestamp 1587416550
transform -1 0 218200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1076
timestamp 1587416550
transform -1 0 218400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1077
timestamp 1587416550
transform -1 0 218600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1078
timestamp 1587416550
transform -1 0 218800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1079
timestamp 1587416550
transform -1 0 219000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1080
timestamp 1587416550
transform -1 0 219200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1081
timestamp 1587416550
transform -1 0 219400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1082
timestamp 1587416550
transform -1 0 219600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1083
timestamp 1587416550
transform -1 0 219800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1084
timestamp 1587416550
transform -1 0 220000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1085
timestamp 1587416550
transform -1 0 220200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1086
timestamp 1587416550
transform -1 0 220400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1087
timestamp 1587416550
transform -1 0 220600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1088
timestamp 1587416550
transform -1 0 220800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1089
timestamp 1587416550
transform -1 0 221000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1090
timestamp 1587416550
transform -1 0 221200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1091
timestamp 1587416550
transform -1 0 221400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1092
timestamp 1587416550
transform -1 0 221600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1093
timestamp 1587416550
transform -1 0 221800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1094
timestamp 1587416550
transform -1 0 222000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1095
timestamp 1587416550
transform -1 0 222200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1096
timestamp 1587416550
transform -1 0 222400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1097
timestamp 1587416550
transform -1 0 222600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1098
timestamp 1587416550
transform -1 0 222800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1099
timestamp 1587416550
transform -1 0 223000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1106
timestamp 1587416550
transform -1 0 224400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1105
timestamp 1587416550
transform -1 0 224200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1104
timestamp 1587416550
transform -1 0 224000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1103
timestamp 1587416550
transform -1 0 223800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1102
timestamp 1587416550
transform -1 0 223600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1101
timestamp 1587416550
transform -1 0 223400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1100
timestamp 1587416550
transform -1 0 223200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__vddio_hvc_pad  sky130_ef_io__vddio_hvc_pad_0 /usr/share/pdk/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1587416550
transform -1 0 239400 0 -1 259093
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1109
timestamp 1587416550
transform -1 0 239800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1108
timestamp 1587416550
transform -1 0 239600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1111
timestamp 1587416550
transform -1 0 240200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1110
timestamp 1587416550
transform -1 0 240000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1112
timestamp 1587416550
transform -1 0 240400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1113
timestamp 1587416550
transform -1 0 240600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1114
timestamp 1587416550
transform -1 0 240800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1115
timestamp 1587416550
transform -1 0 241000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1116
timestamp 1587416550
transform -1 0 241200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1117
timestamp 1587416550
transform -1 0 241400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1118
timestamp 1587416550
transform -1 0 241600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1119
timestamp 1587416550
transform -1 0 241800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1120
timestamp 1587416550
transform -1 0 242000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1121
timestamp 1587416550
transform -1 0 242200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1122
timestamp 1587416550
transform -1 0 242400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1123
timestamp 1587416550
transform -1 0 242600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1124
timestamp 1587416550
transform -1 0 242800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1125
timestamp 1587416550
transform -1 0 243000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1126
timestamp 1587416550
transform -1 0 243200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1127
timestamp 1587416550
transform -1 0 243400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1128
timestamp 1587416550
transform -1 0 243600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1129
timestamp 1587416550
transform -1 0 243800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1130
timestamp 1587416550
transform -1 0 244000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1131
timestamp 1587416550
transform -1 0 244200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1132
timestamp 1587416550
transform -1 0 244400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1133
timestamp 1587416550
transform -1 0 244600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1134
timestamp 1587416550
transform -1 0 244800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1135
timestamp 1587416550
transform -1 0 245000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1136
timestamp 1587416550
transform -1 0 245200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1137
timestamp 1587416550
transform -1 0 245400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1138
timestamp 1587416550
transform -1 0 245600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1139
timestamp 1587416550
transform -1 0 245800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1140
timestamp 1587416550
transform -1 0 246000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1141
timestamp 1587416550
transform -1 0 246200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1142
timestamp 1587416550
transform -1 0 246400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1143
timestamp 1587416550
transform -1 0 246600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1144
timestamp 1587416550
transform -1 0 246800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1145
timestamp 1587416550
transform -1 0 247000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1146
timestamp 1587416550
transform -1 0 247200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1147
timestamp 1587416550
transform -1 0 247400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1148
timestamp 1587416550
transform -1 0 247600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1149
timestamp 1587416550
transform -1 0 247800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1150
timestamp 1587416550
transform -1 0 248000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1151
timestamp 1587416550
transform -1 0 248200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1152
timestamp 1587416550
transform -1 0 248400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1153
timestamp 1587416550
transform -1 0 248600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1154
timestamp 1587416550
transform -1 0 248800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1155
timestamp 1587416550
transform -1 0 249000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1156
timestamp 1587416550
transform -1 0 249200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1157
timestamp 1587416550
transform -1 0 249400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1158
timestamp 1587416550
transform -1 0 249600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1159
timestamp 1587416550
transform -1 0 249800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1160
timestamp 1587416550
transform -1 0 250000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1161
timestamp 1587416550
transform -1 0 250200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1162
timestamp 1587416550
transform -1 0 250400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1163
timestamp 1587416550
transform -1 0 250600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1164
timestamp 1587416550
transform -1 0 250800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1165
timestamp 1587416550
transform -1 0 251000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1166
timestamp 1587416550
transform -1 0 251200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1167
timestamp 1587416550
transform -1 0 251400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1168
timestamp 1587416550
transform -1 0 251600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1169
timestamp 1587416550
transform -1 0 251800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1170
timestamp 1587416550
transform -1 0 252000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1171
timestamp 1587416550
transform -1 0 252200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1172
timestamp 1587416550
transform -1 0 252400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1173
timestamp 1587416550
transform -1 0 252600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1174
timestamp 1587416550
transform -1 0 252800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1175
timestamp 1587416550
transform -1 0 253000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1176
timestamp 1587416550
transform -1 0 253200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1177
timestamp 1587416550
transform -1 0 253400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1178
timestamp 1587416550
transform -1 0 253600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1179
timestamp 1587416550
transform -1 0 253800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1180
timestamp 1587416550
transform -1 0 254000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1181
timestamp 1587416550
transform -1 0 254200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1182
timestamp 1587416550
transform -1 0 254400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1183
timestamp 1587416550
transform -1 0 254600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1184
timestamp 1587416550
transform -1 0 254800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1185
timestamp 1587416550
transform -1 0 255000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1186
timestamp 1587416550
transform -1 0 255200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1187
timestamp 1587416550
transform -1 0 255400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1188
timestamp 1587416550
transform -1 0 255600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1189
timestamp 1587416550
transform -1 0 255800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1190
timestamp 1587416550
transform -1 0 256000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__vdda_lvc_pad  vdd3v3lclamp[2] /usr/share/pdk/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1587416550
transform -1 0 271000 0 -1 259093
box 0 -7 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1192
timestamp 1587416550
transform -1 0 271200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1193
timestamp 1587416550
transform -1 0 271400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1194
timestamp 1587416550
transform -1 0 271600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1195
timestamp 1587416550
transform -1 0 271800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1196
timestamp 1587416550
transform -1 0 272000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1197
timestamp 1587416550
transform -1 0 272200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1198
timestamp 1587416550
transform -1 0 272400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1199
timestamp 1587416550
transform -1 0 272600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1200
timestamp 1587416550
transform -1 0 272800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1201
timestamp 1587416550
transform -1 0 273000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1202
timestamp 1587416550
transform -1 0 273200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1203
timestamp 1587416550
transform -1 0 273400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1204
timestamp 1587416550
transform -1 0 273600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1206
timestamp 1587416550
transform -1 0 274000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1205
timestamp 1587416550
transform -1 0 273800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1208
timestamp 1587416550
transform -1 0 274400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1207
timestamp 1587416550
transform -1 0 274200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1209
timestamp 1587416550
transform -1 0 274600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1210
timestamp 1587416550
transform -1 0 274800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1211
timestamp 1587416550
transform -1 0 275000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1212
timestamp 1587416550
transform -1 0 275200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1213
timestamp 1587416550
transform -1 0 275400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1214
timestamp 1587416550
transform -1 0 275600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1216
timestamp 1587416550
transform -1 0 276000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1215
timestamp 1587416550
transform -1 0 275800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1218
timestamp 1587416550
transform -1 0 276400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1217
timestamp 1587416550
transform -1 0 276200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1219
timestamp 1587416550
transform -1 0 276600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1220
timestamp 1587416550
transform -1 0 276800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1221
timestamp 1587416550
transform -1 0 277000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1222
timestamp 1587416550
transform -1 0 277200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1223
timestamp 1587416550
transform -1 0 277400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1224
timestamp 1587416550
transform -1 0 277600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1225
timestamp 1587416550
transform -1 0 277800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1226
timestamp 1587416550
transform -1 0 278000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1227
timestamp 1587416550
transform -1 0 278200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1229
timestamp 1587416550
transform -1 0 278600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1228
timestamp 1587416550
transform -1 0 278400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1230
timestamp 1587416550
transform -1 0 278800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1231
timestamp 1587416550
transform -1 0 279000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1232
timestamp 1587416550
transform -1 0 279200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1233
timestamp 1587416550
transform -1 0 279400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1234
timestamp 1587416550
transform -1 0 279600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1235
timestamp 1587416550
transform -1 0 279800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1236
timestamp 1587416550
transform -1 0 280000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1237
timestamp 1587416550
transform -1 0 280200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1238
timestamp 1587416550
transform -1 0 280400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1239
timestamp 1587416550
transform -1 0 280600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1240
timestamp 1587416550
transform -1 0 280800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1241
timestamp 1587416550
transform -1 0 281000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1242
timestamp 1587416550
transform -1 0 281200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1243
timestamp 1587416550
transform -1 0 281400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1244
timestamp 1587416550
transform -1 0 281600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1245
timestamp 1587416550
transform -1 0 281800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1246
timestamp 1587416550
transform -1 0 282000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1247
timestamp 1587416550
transform -1 0 282200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1248
timestamp 1587416550
transform -1 0 282400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1249
timestamp 1587416550
transform -1 0 282600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1250
timestamp 1587416550
transform -1 0 282800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1251
timestamp 1587416550
transform -1 0 283000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1252
timestamp 1587416550
transform -1 0 283200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1253
timestamp 1587416550
transform -1 0 283400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1254
timestamp 1587416550
transform -1 0 283600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1255
timestamp 1587416550
transform -1 0 283800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1256
timestamp 1587416550
transform -1 0 284000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1257
timestamp 1587416550
transform -1 0 284200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1258
timestamp 1587416550
transform -1 0 284400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1259
timestamp 1587416550
transform -1 0 284600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1260
timestamp 1587416550
transform -1 0 284800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1261
timestamp 1587416550
transform -1 0 285000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1262
timestamp 1587416550
transform -1 0 285200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1263
timestamp 1587416550
transform -1 0 285400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1264
timestamp 1587416550
transform -1 0 285600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1265
timestamp 1587416550
transform -1 0 285800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1266
timestamp 1587416550
transform -1 0 286000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1267
timestamp 1587416550
transform -1 0 286200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1268
timestamp 1587416550
transform -1 0 286400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1269
timestamp 1587416550
transform -1 0 286600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1270
timestamp 1587416550
transform -1 0 286800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1271
timestamp 1587416550
transform -1 0 287000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1272
timestamp 1587416550
transform -1 0 287200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1273
timestamp 1587416550
transform -1 0 287400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1274
timestamp 1587416550
transform -1 0 287600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__vccd_lvc_pad  vdd1v8lclamp[0] /usr/share/pdk/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1587416550
transform -1 0 302600 0 -1 259093
box 0 -7 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1276
timestamp 1587416550
transform -1 0 302800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1277
timestamp 1587416550
transform -1 0 303000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1278
timestamp 1587416550
transform -1 0 303200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1279
timestamp 1587416550
transform -1 0 303400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1280
timestamp 1587416550
transform -1 0 303600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1281
timestamp 1587416550
transform -1 0 303800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1282
timestamp 1587416550
transform -1 0 304000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1283
timestamp 1587416550
transform -1 0 304200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1285
timestamp 1587416550
transform -1 0 304600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1284
timestamp 1587416550
transform -1 0 304400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1286
timestamp 1587416550
transform -1 0 304800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1287
timestamp 1587416550
transform -1 0 305000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1288
timestamp 1587416550
transform -1 0 305200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1289
timestamp 1587416550
transform -1 0 305400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1290
timestamp 1587416550
transform -1 0 305600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1291
timestamp 1587416550
transform -1 0 305800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1292
timestamp 1587416550
transform -1 0 306000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1293
timestamp 1587416550
transform -1 0 306200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1294
timestamp 1587416550
transform -1 0 306400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1295
timestamp 1587416550
transform -1 0 306600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1296
timestamp 1587416550
transform -1 0 306800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1297
timestamp 1587416550
transform -1 0 307000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1298
timestamp 1587416550
transform -1 0 307200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1299
timestamp 1587416550
transform -1 0 307400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1300
timestamp 1587416550
transform -1 0 307600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1301
timestamp 1587416550
transform -1 0 307800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1302
timestamp 1587416550
transform -1 0 308000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1303
timestamp 1587416550
transform -1 0 308200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1304
timestamp 1587416550
transform -1 0 308400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1305
timestamp 1587416550
transform -1 0 308600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1306
timestamp 1587416550
transform -1 0 308800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1307
timestamp 1587416550
transform -1 0 309000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1308
timestamp 1587416550
transform -1 0 309200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1309
timestamp 1587416550
transform -1 0 309400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1310
timestamp 1587416550
transform -1 0 309600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1311
timestamp 1587416550
transform -1 0 309800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1312
timestamp 1587416550
transform -1 0 310000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1313
timestamp 1587416550
transform -1 0 310200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1314
timestamp 1587416550
transform -1 0 310400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1315
timestamp 1587416550
transform -1 0 310600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1316
timestamp 1587416550
transform -1 0 310800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1317
timestamp 1587416550
transform -1 0 311000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1318
timestamp 1587416550
transform -1 0 311200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1319
timestamp 1587416550
transform -1 0 311400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1320
timestamp 1587416550
transform -1 0 311600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1321
timestamp 1587416550
transform -1 0 311800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1322
timestamp 1587416550
transform -1 0 312000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1323
timestamp 1587416550
transform -1 0 312200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1324
timestamp 1587416550
transform -1 0 312400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1325
timestamp 1587416550
transform -1 0 312600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1326
timestamp 1587416550
transform -1 0 312800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1327
timestamp 1587416550
transform -1 0 313000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1328
timestamp 1587416550
transform -1 0 313200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1329
timestamp 1587416550
transform -1 0 313400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1330
timestamp 1587416550
transform -1 0 313600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1331
timestamp 1587416550
transform -1 0 313800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1332
timestamp 1587416550
transform -1 0 314000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1333
timestamp 1587416550
transform -1 0 314200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1334
timestamp 1587416550
transform -1 0 314400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1335
timestamp 1587416550
transform -1 0 314600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1336
timestamp 1587416550
transform -1 0 314800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1337
timestamp 1587416550
transform -1 0 315000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1338
timestamp 1587416550
transform -1 0 315200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1339
timestamp 1587416550
transform -1 0 315400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1340
timestamp 1587416550
transform -1 0 315600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1341
timestamp 1587416550
transform -1 0 315800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1342
timestamp 1587416550
transform -1 0 316000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1343
timestamp 1587416550
transform -1 0 316200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1344
timestamp 1587416550
transform -1 0 316400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1345
timestamp 1587416550
transform -1 0 316600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1346
timestamp 1587416550
transform -1 0 316800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1347
timestamp 1587416550
transform -1 0 317000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1348
timestamp 1587416550
transform -1 0 317200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1349
timestamp 1587416550
transform -1 0 317400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1350
timestamp 1587416550
transform -1 0 317600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1351
timestamp 1587416550
transform -1 0 317800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1352
timestamp 1587416550
transform -1 0 318000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1353
timestamp 1587416550
transform -1 0 318200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1354
timestamp 1587416550
transform -1 0 318400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1355
timestamp 1587416550
transform -1 0 318600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1356
timestamp 1587416550
transform -1 0 318800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1357
timestamp 1587416550
transform -1 0 319000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1358
timestamp 1587416550
transform -1 0 319200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__vssa_hvc_pad  vsshclamp[1] /usr/share/pdk/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1587416550
transform -1 0 334200 0 -1 259093
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1360
timestamp 1587416550
transform -1 0 334400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1361
timestamp 1587416550
transform -1 0 334600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1362
timestamp 1587416550
transform -1 0 334800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1364
timestamp 1587416550
transform -1 0 335200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1363
timestamp 1587416550
transform -1 0 335000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1365
timestamp 1587416550
transform -1 0 335400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1366
timestamp 1587416550
transform -1 0 335600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1367
timestamp 1587416550
transform -1 0 335800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1368
timestamp 1587416550
transform -1 0 336000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1369
timestamp 1587416550
transform -1 0 336200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1370
timestamp 1587416550
transform -1 0 336400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1371
timestamp 1587416550
transform -1 0 336600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1372
timestamp 1587416550
transform -1 0 336800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1373
timestamp 1587416550
transform -1 0 337000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1374
timestamp 1587416550
transform -1 0 337200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1375
timestamp 1587416550
transform -1 0 337400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1376
timestamp 1587416550
transform -1 0 337600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1377
timestamp 1587416550
transform -1 0 337800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1378
timestamp 1587416550
transform -1 0 338000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1379
timestamp 1587416550
transform -1 0 338200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1380
timestamp 1587416550
transform -1 0 338400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1381
timestamp 1587416550
transform -1 0 338600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1382
timestamp 1587416550
transform -1 0 338800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1383
timestamp 1587416550
transform -1 0 339000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1384
timestamp 1587416550
transform -1 0 339200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1385
timestamp 1587416550
transform -1 0 339400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1386
timestamp 1587416550
transform -1 0 339600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1387
timestamp 1587416550
transform -1 0 339800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1388
timestamp 1587416550
transform -1 0 340000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1389
timestamp 1587416550
transform -1 0 340200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1390
timestamp 1587416550
transform -1 0 340400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1391
timestamp 1587416550
transform -1 0 340600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1392
timestamp 1587416550
transform -1 0 340800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1393
timestamp 1587416550
transform -1 0 341000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1394
timestamp 1587416550
transform -1 0 341200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1395
timestamp 1587416550
transform -1 0 341400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1396
timestamp 1587416550
transform -1 0 341600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1397
timestamp 1587416550
transform -1 0 341800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1398
timestamp 1587416550
transform -1 0 342000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1399
timestamp 1587416550
transform -1 0 342200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1400
timestamp 1587416550
transform -1 0 342400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1401
timestamp 1587416550
transform -1 0 342600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1402
timestamp 1587416550
transform -1 0 342800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1403
timestamp 1587416550
transform -1 0 343000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1404
timestamp 1587416550
transform -1 0 343200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1405
timestamp 1587416550
transform -1 0 343400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1406
timestamp 1587416550
transform -1 0 343600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1407
timestamp 1587416550
transform -1 0 343800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1408
timestamp 1587416550
transform -1 0 344000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1409
timestamp 1587416550
transform -1 0 344200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1410
timestamp 1587416550
transform -1 0 344400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1411
timestamp 1587416550
transform -1 0 344600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1412
timestamp 1587416550
transform -1 0 344800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1413
timestamp 1587416550
transform -1 0 345000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1414
timestamp 1587416550
transform -1 0 345200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1415
timestamp 1587416550
transform -1 0 345400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1416
timestamp 1587416550
transform -1 0 345600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1417
timestamp 1587416550
transform -1 0 345800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1418
timestamp 1587416550
transform -1 0 346000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1419
timestamp 1587416550
transform -1 0 346200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1420
timestamp 1587416550
transform -1 0 346400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1421
timestamp 1587416550
transform -1 0 346600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1422
timestamp 1587416550
transform -1 0 346800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1423
timestamp 1587416550
transform -1 0 347000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1424
timestamp 1587416550
transform -1 0 347200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1425
timestamp 1587416550
transform -1 0 347400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1426
timestamp 1587416550
transform -1 0 347600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1427
timestamp 1587416550
transform -1 0 347800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1428
timestamp 1587416550
transform -1 0 348000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1429
timestamp 1587416550
transform -1 0 348200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1430
timestamp 1587416550
transform -1 0 348400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1431
timestamp 1587416550
transform -1 0 348600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1432
timestamp 1587416550
transform -1 0 348800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1433
timestamp 1587416550
transform -1 0 349000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1434
timestamp 1587416550
transform -1 0 349200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1435
timestamp 1587416550
transform -1 0 349400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1436
timestamp 1587416550
transform -1 0 349600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1437
timestamp 1587416550
transform -1 0 349800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1438
timestamp 1587416550
transform -1 0 350000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1439
timestamp 1587416550
transform -1 0 350200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1440
timestamp 1587416550
transform -1 0 350400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1441
timestamp 1587416550
transform -1 0 350600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1442
timestamp 1587416550
transform -1 0 350800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__vssio_lvc_pad  vssiolclamp /usr/share/pdk/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1587416550
transform -1 0 365800 0 -1 259093
box 0 -7 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1444
timestamp 1587416550
transform -1 0 366000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1445
timestamp 1587416550
transform -1 0 366200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1446
timestamp 1587416550
transform -1 0 366400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1447
timestamp 1587416550
transform -1 0 366600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1448
timestamp 1587416550
transform -1 0 366800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2282
timestamp 1587416550
transform 0 -1 207593 1 0 260300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2283
timestamp 1587416550
transform 0 -1 207593 1 0 260500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2284
timestamp 1587416550
transform 0 -1 207593 1 0 260700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2285
timestamp 1587416550
transform 0 -1 207593 1 0 260900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2286
timestamp 1587416550
transform 0 -1 207593 1 0 261100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2287
timestamp 1587416550
transform 0 -1 207593 1 0 261300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2288
timestamp 1587416550
transform 0 -1 207593 1 0 261500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2289
timestamp 1587416550
transform 0 -1 207593 1 0 261700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2290
timestamp 1587416550
transform 0 -1 207593 1 0 261900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2291
timestamp 1587416550
transform 0 -1 207593 1 0 262100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2292
timestamp 1587416550
transform 0 -1 207593 1 0 262300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2293
timestamp 1587416550
transform 0 -1 207593 1 0 262500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2294
timestamp 1587416550
transform 0 -1 207593 1 0 262700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2295
timestamp 1587416550
transform 0 -1 207593 1 0 262900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2296
timestamp 1587416550
transform 0 -1 207593 1 0 263100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2297
timestamp 1587416550
transform 0 -1 207593 1 0 263300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2298
timestamp 1587416550
transform 0 -1 207593 1 0 263500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2299
timestamp 1587416550
transform 0 -1 207593 1 0 263700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2300
timestamp 1587416550
transform 0 -1 207593 1 0 263900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2301
timestamp 1587416550
transform 0 -1 207593 1 0 264100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2302
timestamp 1587416550
transform 0 -1 207593 1 0 264300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2303
timestamp 1587416550
transform 0 -1 207593 1 0 264500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2304
timestamp 1587416550
transform 0 -1 207593 1 0 264700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2305
timestamp 1587416550
transform 0 -1 207593 1 0 264900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2306
timestamp 1587416550
transform 0 -1 207593 1 0 265100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2307
timestamp 1587416550
transform 0 -1 207593 1 0 265300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2308
timestamp 1587416550
transform 0 -1 207593 1 0 265500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2309
timestamp 1587416550
transform 0 -1 207593 1 0 265700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2310
timestamp 1587416550
transform 0 -1 207593 1 0 265900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2311
timestamp 1587416550
transform 0 -1 207593 1 0 266100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2312
timestamp 1587416550
transform 0 -1 207593 1 0 266300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2313
timestamp 1587416550
transform 0 -1 207593 1 0 266500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2314
timestamp 1587416550
transform 0 -1 207593 1 0 266700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2315
timestamp 1587416550
transform 0 -1 207593 1 0 266900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2316
timestamp 1587416550
transform 0 -1 207593 1 0 267100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2317
timestamp 1587416550
transform 0 -1 207593 1 0 267300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2318
timestamp 1587416550
transform 0 -1 207593 1 0 267500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2319
timestamp 1587416550
transform 0 -1 207593 1 0 267700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2320
timestamp 1587416550
transform 0 -1 207593 1 0 267900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2321
timestamp 1587416550
transform 0 -1 207593 1 0 268100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2322
timestamp 1587416550
transform 0 -1 207593 1 0 268300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2323
timestamp 1587416550
transform 0 -1 207593 1 0 268500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2324
timestamp 1587416550
transform 0 -1 207593 1 0 268700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2325
timestamp 1587416550
transform 0 -1 207593 1 0 268900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2326
timestamp 1587416550
transform 0 -1 207593 1 0 269100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2327
timestamp 1587416550
transform 0 -1 207593 1 0 269300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2328
timestamp 1587416550
transform 0 -1 207593 1 0 269500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2329
timestamp 1587416550
transform 0 -1 207593 1 0 269700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2330
timestamp 1587416550
transform 0 -1 207593 1 0 269900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2331
timestamp 1587416550
transform 0 -1 207593 1 0 270100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2332
timestamp 1587416550
transform 0 -1 207593 1 0 270300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2333
timestamp 1587416550
transform 0 -1 207593 1 0 270500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2334
timestamp 1587416550
transform 0 -1 207593 1 0 270700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2335
timestamp 1587416550
transform 0 -1 207593 1 0 270900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2336
timestamp 1587416550
transform 0 -1 207593 1 0 271100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2337
timestamp 1587416550
transform 0 -1 207593 1 0 271300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2338
timestamp 1587416550
transform 0 -1 207593 1 0 271500
box 0 0 200 39593
use sky130_ef_io__vdda_hvc_pad  vddiohclamp[1] /usr/share/pdk/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1587416550
transform 0 -1 207593 1 0 271700
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2341
timestamp 1587416550
transform 0 -1 207593 1 0 286900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2340
timestamp 1587416550
transform 0 -1 207593 1 0 286700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2342
timestamp 1587416550
transform 0 -1 207593 1 0 287100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2343
timestamp 1587416550
transform 0 -1 207593 1 0 287300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2345
timestamp 1587416550
transform 0 -1 207593 1 0 287700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2344
timestamp 1587416550
transform 0 -1 207593 1 0 287500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2347
timestamp 1587416550
transform 0 -1 207593 1 0 288100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2346
timestamp 1587416550
transform 0 -1 207593 1 0 287900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2349
timestamp 1587416550
transform 0 -1 207593 1 0 288500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2348
timestamp 1587416550
transform 0 -1 207593 1 0 288300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2350
timestamp 1587416550
transform 0 -1 207593 1 0 288700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2352
timestamp 1587416550
transform 0 -1 207593 1 0 289100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2351
timestamp 1587416550
transform 0 -1 207593 1 0 288900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2353
timestamp 1587416550
transform 0 -1 207593 1 0 289300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2354
timestamp 1587416550
transform 0 -1 207593 1 0 289500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2355
timestamp 1587416550
transform 0 -1 207593 1 0 289700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2356
timestamp 1587416550
transform 0 -1 207593 1 0 289900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2357
timestamp 1587416550
transform 0 -1 207593 1 0 290100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2358
timestamp 1587416550
transform 0 -1 207593 1 0 290300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2359
timestamp 1587416550
transform 0 -1 207593 1 0 290500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2360
timestamp 1587416550
transform 0 -1 207593 1 0 290700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2361
timestamp 1587416550
transform 0 -1 207593 1 0 290900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2362
timestamp 1587416550
transform 0 -1 207593 1 0 291100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2363
timestamp 1587416550
transform 0 -1 207593 1 0 291300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2364
timestamp 1587416550
transform 0 -1 207593 1 0 291500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2365
timestamp 1587416550
transform 0 -1 207593 1 0 291700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2366
timestamp 1587416550
transform 0 -1 207593 1 0 291900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2367
timestamp 1587416550
transform 0 -1 207593 1 0 292100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2368
timestamp 1587416550
transform 0 -1 207593 1 0 292300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2369
timestamp 1587416550
transform 0 -1 207593 1 0 292500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2370
timestamp 1587416550
transform 0 -1 207593 1 0 292700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2371
timestamp 1587416550
transform 0 -1 207593 1 0 292900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2372
timestamp 1587416550
transform 0 -1 207593 1 0 293100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2373
timestamp 1587416550
transform 0 -1 207593 1 0 293300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2374
timestamp 1587416550
transform 0 -1 207593 1 0 293500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2375
timestamp 1587416550
transform 0 -1 207593 1 0 293700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2376
timestamp 1587416550
transform 0 -1 207593 1 0 293900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2377
timestamp 1587416550
transform 0 -1 207593 1 0 294100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2378
timestamp 1587416550
transform 0 -1 207593 1 0 294300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2379
timestamp 1587416550
transform 0 -1 207593 1 0 294500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2380
timestamp 1587416550
transform 0 -1 207593 1 0 294700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2381
timestamp 1587416550
transform 0 -1 207593 1 0 294900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2382
timestamp 1587416550
transform 0 -1 207593 1 0 295100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2383
timestamp 1587416550
transform 0 -1 207593 1 0 295300
box 0 0 200 39593
use striVe_clkrst  clkrst
timestamp 1587660775
transform 1 0 228000 0 1 280300
box 0 0 4543 4543
use sky130_ef_io__com_bus_slice_1um  FILLER_2384
timestamp 1587416550
transform 0 -1 207593 1 0 295500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2385
timestamp 1587416550
transform 0 -1 207593 1 0 295700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2386
timestamp 1587416550
transform 0 -1 207593 1 0 295900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2387
timestamp 1587416550
transform 0 -1 207593 1 0 296100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2388
timestamp 1587416550
transform 0 -1 207593 1 0 296300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2389
timestamp 1587416550
transform 0 -1 207593 1 0 296500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2390
timestamp 1587416550
transform 0 -1 207593 1 0 296700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2391
timestamp 1587416550
transform 0 -1 207593 1 0 296900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2392
timestamp 1587416550
transform 0 -1 207593 1 0 297100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2393
timestamp 1587416550
transform 0 -1 207593 1 0 297300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2394
timestamp 1587416550
transform 0 -1 207593 1 0 297500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2395
timestamp 1587416550
transform 0 -1 207593 1 0 297700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2396
timestamp 1587416550
transform 0 -1 207593 1 0 297900
box 0 0 200 39593
use sky130_ef_io__vdda_lvc_pad  vdd3v3lclamp[3]
timestamp 1587416550
transform 0 -1 207593 1 0 298100
box 0 -7 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2398
timestamp 1587416550
transform 0 -1 207593 1 0 313100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2399
timestamp 1587416550
transform 0 -1 207593 1 0 313300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2400
timestamp 1587416550
transform 0 -1 207593 1 0 313500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2401
timestamp 1587416550
transform 0 -1 207593 1 0 313700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2402
timestamp 1587416550
transform 0 -1 207593 1 0 313900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2403
timestamp 1587416550
transform 0 -1 207593 1 0 314100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2404
timestamp 1587416550
transform 0 -1 207593 1 0 314300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2405
timestamp 1587416550
transform 0 -1 207593 1 0 314500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2407
timestamp 1587416550
transform 0 -1 207593 1 0 314900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2406
timestamp 1587416550
transform 0 -1 207593 1 0 314700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2408
timestamp 1587416550
transform 0 -1 207593 1 0 315100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2409
timestamp 1587416550
transform 0 -1 207593 1 0 315300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2410
timestamp 1587416550
transform 0 -1 207593 1 0 315500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2411
timestamp 1587416550
transform 0 -1 207593 1 0 315700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2412
timestamp 1587416550
transform 0 -1 207593 1 0 315900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2413
timestamp 1587416550
transform 0 -1 207593 1 0 316100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2414
timestamp 1587416550
transform 0 -1 207593 1 0 316300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2415
timestamp 1587416550
transform 0 -1 207593 1 0 316500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2416
timestamp 1587416550
transform 0 -1 207593 1 0 316700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2417
timestamp 1587416550
transform 0 -1 207593 1 0 316900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2418
timestamp 1587416550
transform 0 -1 207593 1 0 317100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2419
timestamp 1587416550
transform 0 -1 207593 1 0 317300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2420
timestamp 1587416550
transform 0 -1 207593 1 0 317500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2421
timestamp 1587416550
transform 0 -1 207593 1 0 317700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2422
timestamp 1587416550
transform 0 -1 207593 1 0 317900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2423
timestamp 1587416550
transform 0 -1 207593 1 0 318100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2424
timestamp 1587416550
transform 0 -1 207593 1 0 318300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2425
timestamp 1587416550
transform 0 -1 207593 1 0 318500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2426
timestamp 1587416550
transform 0 -1 207593 1 0 318700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2427
timestamp 1587416550
transform 0 -1 207593 1 0 318900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2428
timestamp 1587416550
transform 0 -1 207593 1 0 319100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2429
timestamp 1587416550
transform 0 -1 207593 1 0 319300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2430
timestamp 1587416550
transform 0 -1 207593 1 0 319500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2431
timestamp 1587416550
transform 0 -1 207593 1 0 319700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2432
timestamp 1587416550
transform 0 -1 207593 1 0 319900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2433
timestamp 1587416550
transform 0 -1 207593 1 0 320100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2434
timestamp 1587416550
transform 0 -1 207593 1 0 320300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2435
timestamp 1587416550
transform 0 -1 207593 1 0 320500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2436
timestamp 1587416550
transform 0 -1 207593 1 0 320700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2437
timestamp 1587416550
transform 0 -1 207593 1 0 320900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2438
timestamp 1587416550
transform 0 -1 207593 1 0 321100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2439
timestamp 1587416550
transform 0 -1 207593 1 0 321300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2440
timestamp 1587416550
transform 0 -1 207593 1 0 321500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2441
timestamp 1587416550
transform 0 -1 207593 1 0 321700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2442
timestamp 1587416550
transform 0 -1 207593 1 0 321900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2443
timestamp 1587416550
transform 0 -1 207593 1 0 322100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2444
timestamp 1587416550
transform 0 -1 207593 1 0 322300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2445
timestamp 1587416550
transform 0 -1 207593 1 0 322500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2446
timestamp 1587416550
transform 0 -1 207593 1 0 322700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2447
timestamp 1587416550
transform 0 -1 207593 1 0 322900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2448
timestamp 1587416550
transform 0 -1 207593 1 0 323100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2449
timestamp 1587416550
transform 0 -1 207593 1 0 323300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2450
timestamp 1587416550
transform 0 -1 207593 1 0 323500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2451
timestamp 1587416550
transform 0 -1 207593 1 0 323700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2453
timestamp 1587416550
transform 0 -1 207593 1 0 324100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2452
timestamp 1587416550
transform 0 -1 207593 1 0 323900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2454
timestamp 1587416550
transform 0 -1 207593 1 0 324300
box 0 0 200 39593
use sky130_ef_io__vccd_lvc_pad  vdd1v8lclamp[1]
timestamp 1587416550
transform 0 -1 207593 1 0 324500
box 0 -7 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2456
timestamp 1587416550
transform 0 -1 207593 1 0 339500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2457
timestamp 1587416550
transform 0 -1 207593 1 0 339700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2461
timestamp 1587416550
transform 0 -1 207593 1 0 340500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2458
timestamp 1587416550
transform 0 -1 207593 1 0 339900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2459
timestamp 1587416550
transform 0 -1 207593 1 0 340100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2460
timestamp 1587416550
transform 0 -1 207593 1 0 340300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2462
timestamp 1587416550
transform 0 -1 207593 1 0 340700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2463
timestamp 1587416550
transform 0 -1 207593 1 0 340900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2464
timestamp 1587416550
transform 0 -1 207593 1 0 341100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2465
timestamp 1587416550
transform 0 -1 207593 1 0 341300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2466
timestamp 1587416550
transform 0 -1 207593 1 0 341500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2467
timestamp 1587416550
transform 0 -1 207593 1 0 341700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2468
timestamp 1587416550
transform 0 -1 207593 1 0 341900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2469
timestamp 1587416550
transform 0 -1 207593 1 0 342100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2470
timestamp 1587416550
transform 0 -1 207593 1 0 342300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2471
timestamp 1587416550
transform 0 -1 207593 1 0 342500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2472
timestamp 1587416550
transform 0 -1 207593 1 0 342700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2473
timestamp 1587416550
transform 0 -1 207593 1 0 342900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2474
timestamp 1587416550
transform 0 -1 207593 1 0 343100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2475
timestamp 1587416550
transform 0 -1 207593 1 0 343300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2476
timestamp 1587416550
transform 0 -1 207593 1 0 343500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2477
timestamp 1587416550
transform 0 -1 207593 1 0 343700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2478
timestamp 1587416550
transform 0 -1 207593 1 0 343900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2479
timestamp 1587416550
transform 0 -1 207593 1 0 344100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2480
timestamp 1587416550
transform 0 -1 207593 1 0 344300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2481
timestamp 1587416550
transform 0 -1 207593 1 0 344500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2482
timestamp 1587416550
transform 0 -1 207593 1 0 344700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2483
timestamp 1587416550
transform 0 -1 207593 1 0 344900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2484
timestamp 1587416550
transform 0 -1 207593 1 0 345100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2485
timestamp 1587416550
transform 0 -1 207593 1 0 345300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2486
timestamp 1587416550
transform 0 -1 207593 1 0 345500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2487
timestamp 1587416550
transform 0 -1 207593 1 0 345700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2488
timestamp 1587416550
transform 0 -1 207593 1 0 345900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2489
timestamp 1587416550
transform 0 -1 207593 1 0 346100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2490
timestamp 1587416550
transform 0 -1 207593 1 0 346300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2491
timestamp 1587416550
transform 0 -1 207593 1 0 346500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2492
timestamp 1587416550
transform 0 -1 207593 1 0 346700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2493
timestamp 1587416550
transform 0 -1 207593 1 0 346900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2494
timestamp 1587416550
transform 0 -1 207593 1 0 347100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2495
timestamp 1587416550
transform 0 -1 207593 1 0 347300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2496
timestamp 1587416550
transform 0 -1 207593 1 0 347500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2497
timestamp 1587416550
transform 0 -1 207593 1 0 347700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2498
timestamp 1587416550
transform 0 -1 207593 1 0 347900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2499
timestamp 1587416550
transform 0 -1 207593 1 0 348100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2500
timestamp 1587416550
transform 0 -1 207593 1 0 348300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2501
timestamp 1587416550
transform 0 -1 207593 1 0 348500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2502
timestamp 1587416550
transform 0 -1 207593 1 0 348700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2503
timestamp 1587416550
transform 0 -1 207593 1 0 348900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2504
timestamp 1587416550
transform 0 -1 207593 1 0 349100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2505
timestamp 1587416550
transform 0 -1 207593 1 0 349300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2506
timestamp 1587416550
transform 0 -1 207593 1 0 349500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2507
timestamp 1587416550
transform 0 -1 207593 1 0 349700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2508
timestamp 1587416550
transform 0 -1 207593 1 0 349900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2509
timestamp 1587416550
transform 0 -1 207593 1 0 350100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2510
timestamp 1587416550
transform 0 -1 207593 1 0 350300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2511
timestamp 1587416550
transform 0 -1 207593 1 0 350500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2512
timestamp 1587416550
transform 0 -1 207593 1 0 350700
box 0 0 200 39593
use sky130_ef_io__vssa_hvc_pad  vsshclamp[2]
timestamp 1587416550
transform 0 -1 207593 1 0 350900
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2515
timestamp 1587416550
transform 0 -1 207593 1 0 366100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2514
timestamp 1587416550
transform 0 -1 207593 1 0 365900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2516
timestamp 1587416550
transform 0 -1 207593 1 0 366300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2518
timestamp 1587416550
transform 0 -1 207593 1 0 366700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2517
timestamp 1587416550
transform 0 -1 207593 1 0 366500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2519
timestamp 1587416550
transform 0 -1 207593 1 0 366900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2520
timestamp 1587416550
transform 0 -1 207593 1 0 367100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2521
timestamp 1587416550
transform 0 -1 207593 1 0 367300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2522
timestamp 1587416550
transform 0 -1 207593 1 0 367500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2523
timestamp 1587416550
transform 0 -1 207593 1 0 367700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2524
timestamp 1587416550
transform 0 -1 207593 1 0 367900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2525
timestamp 1587416550
transform 0 -1 207593 1 0 368100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2526
timestamp 1587416550
transform 0 -1 207593 1 0 368300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2527
timestamp 1587416550
transform 0 -1 207593 1 0 368500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2529
timestamp 1587416550
transform 0 -1 207593 1 0 368900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2528
timestamp 1587416550
transform 0 -1 207593 1 0 368700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2531
timestamp 1587416550
transform 0 -1 207593 1 0 369300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2530
timestamp 1587416550
transform 0 -1 207593 1 0 369100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2532
timestamp 1587416550
transform 0 -1 207593 1 0 369500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2534
timestamp 1587416550
transform 0 -1 207593 1 0 369900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2533
timestamp 1587416550
transform 0 -1 207593 1 0 369700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2535
timestamp 1587416550
transform 0 -1 207593 1 0 370100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2536
timestamp 1587416550
transform 0 -1 207593 1 0 370300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2537
timestamp 1587416550
transform 0 -1 207593 1 0 370500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2538
timestamp 1587416550
transform 0 -1 207593 1 0 370700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2539
timestamp 1587416550
transform 0 -1 207593 1 0 370900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2540
timestamp 1587416550
transform 0 -1 207593 1 0 371100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2542
timestamp 1587416550
transform 0 -1 207593 1 0 371500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2541
timestamp 1587416550
transform 0 -1 207593 1 0 371300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2544
timestamp 1587416550
transform 0 -1 207593 1 0 371900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2543
timestamp 1587416550
transform 0 -1 207593 1 0 371700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2545
timestamp 1587416550
transform 0 -1 207593 1 0 372100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2547
timestamp 1587416550
transform 0 -1 207593 1 0 372500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2546
timestamp 1587416550
transform 0 -1 207593 1 0 372300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2548
timestamp 1587416550
transform 0 -1 207593 1 0 372700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2549
timestamp 1587416550
transform 0 -1 207593 1 0 372900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2550
timestamp 1587416550
transform 0 -1 207593 1 0 373100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2551
timestamp 1587416550
transform 0 -1 207593 1 0 373300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2552
timestamp 1587416550
transform 0 -1 207593 1 0 373500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2553
timestamp 1587416550
transform 0 -1 207593 1 0 373700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2554
timestamp 1587416550
transform 0 -1 207593 1 0 373900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2555
timestamp 1587416550
transform 0 -1 207593 1 0 374100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2556
timestamp 1587416550
transform 0 -1 207593 1 0 374300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2557
timestamp 1587416550
transform 0 -1 207593 1 0 374500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2558
timestamp 1587416550
transform 0 -1 207593 1 0 374700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2559
timestamp 1587416550
transform 0 -1 207593 1 0 374900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2560
timestamp 1587416550
transform 0 -1 207593 1 0 375100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2561
timestamp 1587416550
transform 0 -1 207593 1 0 375300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2562
timestamp 1587416550
transform 0 -1 207593 1 0 375500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2563
timestamp 1587416550
transform 0 -1 207593 1 0 375700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2564
timestamp 1587416550
transform 0 -1 207593 1 0 375900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2565
timestamp 1587416550
transform 0 -1 207593 1 0 376100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2566
timestamp 1587416550
transform 0 -1 207593 1 0 376300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2567
timestamp 1587416550
transform 0 -1 207593 1 0 376500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2568
timestamp 1587416550
transform 0 -1 207593 1 0 376700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2570
timestamp 1587416550
transform 0 -1 207593 1 0 377100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2569
timestamp 1587416550
transform 0 -1 207593 1 0 376900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2572
timestamp 1587416550
transform 0 -1 207593 1 0 393300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2573
timestamp 1587416550
transform 0 -1 207593 1 0 393500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2574
timestamp 1587416550
transform 0 -1 207593 1 0 393700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2575
timestamp 1587416550
transform 0 -1 207593 1 0 393900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2576
timestamp 1587416550
transform 0 -1 207593 1 0 394100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2577
timestamp 1587416550
transform 0 -1 207593 1 0 394300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2578
timestamp 1587416550
transform 0 -1 207593 1 0 394500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2579
timestamp 1587416550
transform 0 -1 207593 1 0 394700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2580
timestamp 1587416550
transform 0 -1 207593 1 0 394900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2581
timestamp 1587416550
transform 0 -1 207593 1 0 395100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2582
timestamp 1587416550
transform 0 -1 207593 1 0 395300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2584
timestamp 1587416550
transform 0 -1 207593 1 0 395700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2583
timestamp 1587416550
transform 0 -1 207593 1 0 395500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2585
timestamp 1587416550
transform 0 -1 207593 1 0 395900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2586
timestamp 1587416550
transform 0 -1 207593 1 0 396100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2587
timestamp 1587416550
transform 0 -1 207593 1 0 396300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2588
timestamp 1587416550
transform 0 -1 207593 1 0 396500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2589
timestamp 1587416550
transform 0 -1 207593 1 0 396700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2590
timestamp 1587416550
transform 0 -1 207593 1 0 396900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2591
timestamp 1587416550
transform 0 -1 207593 1 0 397100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2592
timestamp 1587416550
transform 0 -1 207593 1 0 397300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2593
timestamp 1587416550
transform 0 -1 207593 1 0 397500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2594
timestamp 1587416550
transform 0 -1 207593 1 0 397700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2595
timestamp 1587416550
transform 0 -1 207593 1 0 397900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2596
timestamp 1587416550
transform 0 -1 207593 1 0 398100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2597
timestamp 1587416550
transform 0 -1 207593 1 0 398300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2598
timestamp 1587416550
transform 0 -1 207593 1 0 398500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2599
timestamp 1587416550
transform 0 -1 207593 1 0 398700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2600
timestamp 1587416550
transform 0 -1 207593 1 0 398900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2601
timestamp 1587416550
transform 0 -1 207593 1 0 399100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2602
timestamp 1587416550
transform 0 -1 207593 1 0 399300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2603
timestamp 1587416550
transform 0 -1 207593 1 0 399500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2604
timestamp 1587416550
transform 0 -1 207593 1 0 399700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2605
timestamp 1587416550
transform 0 -1 207593 1 0 399900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2606
timestamp 1587416550
transform 0 -1 207593 1 0 400100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2607
timestamp 1587416550
transform 0 -1 207593 1 0 400300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2608
timestamp 1587416550
transform 0 -1 207593 1 0 400500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2609
timestamp 1587416550
transform 0 -1 207593 1 0 400700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2610
timestamp 1587416550
transform 0 -1 207593 1 0 400900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2611
timestamp 1587416550
transform 0 -1 207593 1 0 401100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2612
timestamp 1587416550
transform 0 -1 207593 1 0 401300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2613
timestamp 1587416550
transform 0 -1 207593 1 0 401500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2614
timestamp 1587416550
transform 0 -1 207593 1 0 401700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2615
timestamp 1587416550
transform 0 -1 207593 1 0 401900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2616
timestamp 1587416550
transform 0 -1 207593 1 0 402100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2617
timestamp 1587416550
transform 0 -1 207593 1 0 402300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2618
timestamp 1587416550
transform 0 -1 207593 1 0 402500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2619
timestamp 1587416550
transform 0 -1 207593 1 0 402700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2620
timestamp 1587416550
transform 0 -1 207593 1 0 402900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2621
timestamp 1587416550
transform 0 -1 207593 1 0 403100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2622
timestamp 1587416550
transform 0 -1 207593 1 0 403300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2623
timestamp 1587416550
transform 0 -1 207593 1 0 403500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2624
timestamp 1587416550
transform 0 -1 207593 1 0 403700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2625
timestamp 1587416550
transform 0 -1 207593 1 0 403900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2626
timestamp 1587416550
transform 0 -1 207593 1 0 404100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2627
timestamp 1587416550
transform 0 -1 207593 1 0 404300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2628
timestamp 1587416550
transform 0 -1 207593 1 0 404500
box 0 0 200 39593
use sky130_fd_io__top_xres4v2  RSTB_pad /usr/share/pdk/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1587416550
transform 0 -1 208000 1 0 404700
box -103 0 15124 40000
use sky130_ef_io__com_bus_slice_1um  FILLER_2631
timestamp 1587416550
transform 0 -1 207593 1 0 419900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2630
timestamp 1587416550
transform 0 -1 207593 1 0 419700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2633
timestamp 1587416550
transform 0 -1 207593 1 0 420300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2632
timestamp 1587416550
transform 0 -1 207593 1 0 420100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2636
timestamp 1587416550
transform 0 -1 207593 1 0 420900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2635
timestamp 1587416550
transform 0 -1 207593 1 0 420700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2634
timestamp 1587416550
transform 0 -1 207593 1 0 420500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2640
timestamp 1587416550
transform 0 -1 207593 1 0 421700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2639
timestamp 1587416550
transform 0 -1 207593 1 0 421500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2637
timestamp 1587416550
transform 0 -1 207593 1 0 421100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2638
timestamp 1587416550
transform 0 -1 207593 1 0 421300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2641
timestamp 1587416550
transform 0 -1 207593 1 0 421900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2644
timestamp 1587416550
transform 0 -1 207593 1 0 422500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2643
timestamp 1587416550
transform 0 -1 207593 1 0 422300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2642
timestamp 1587416550
transform 0 -1 207593 1 0 422100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2645
timestamp 1587416550
transform 0 -1 207593 1 0 422700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2646
timestamp 1587416550
transform 0 -1 207593 1 0 422900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2647
timestamp 1587416550
transform 0 -1 207593 1 0 423100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2648
timestamp 1587416550
transform 0 -1 207593 1 0 423300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2649
timestamp 1587416550
transform 0 -1 207593 1 0 423500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2650
timestamp 1587416550
transform 0 -1 207593 1 0 423700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2651
timestamp 1587416550
transform 0 -1 207593 1 0 423900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2652
timestamp 1587416550
transform 0 -1 207593 1 0 424100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2653
timestamp 1587416550
transform 0 -1 207593 1 0 424300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2654
timestamp 1587416550
transform 0 -1 207593 1 0 424500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2655
timestamp 1587416550
transform 0 -1 207593 1 0 424700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2656
timestamp 1587416550
transform 0 -1 207593 1 0 424900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2657
timestamp 1587416550
transform 0 -1 207593 1 0 425100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2658
timestamp 1587416550
transform 0 -1 207593 1 0 425300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2659
timestamp 1587416550
transform 0 -1 207593 1 0 425500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2660
timestamp 1587416550
transform 0 -1 207593 1 0 425700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2661
timestamp 1587416550
transform 0 -1 207593 1 0 425900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2662
timestamp 1587416550
transform 0 -1 207593 1 0 426100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2663
timestamp 1587416550
transform 0 -1 207593 1 0 426300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2664
timestamp 1587416550
transform 0 -1 207593 1 0 426500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2665
timestamp 1587416550
transform 0 -1 207593 1 0 426700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2666
timestamp 1587416550
transform 0 -1 207593 1 0 426900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2667
timestamp 1587416550
transform 0 -1 207593 1 0 427100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2668
timestamp 1587416550
transform 0 -1 207593 1 0 427300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2669
timestamp 1587416550
transform 0 -1 207593 1 0 427500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2670
timestamp 1587416550
transform 0 -1 207593 1 0 427700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2671
timestamp 1587416550
transform 0 -1 207593 1 0 427900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2672
timestamp 1587416550
transform 0 -1 207593 1 0 428100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2673
timestamp 1587416550
transform 0 -1 207593 1 0 428300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2674
timestamp 1587416550
transform 0 -1 207593 1 0 428500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2675
timestamp 1587416550
transform 0 -1 207593 1 0 428700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2676
timestamp 1587416550
transform 0 -1 207593 1 0 428900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2677
timestamp 1587416550
transform 0 -1 207593 1 0 429100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2678
timestamp 1587416550
transform 0 -1 207593 1 0 429300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2679
timestamp 1587416550
transform 0 -1 207593 1 0 429500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2680
timestamp 1587416550
transform 0 -1 207593 1 0 429700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2681
timestamp 1587416550
transform 0 -1 207593 1 0 429900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2682
timestamp 1587416550
transform 0 -1 207593 1 0 430100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2683
timestamp 1587416550
transform 0 -1 207593 1 0 430300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2684
timestamp 1587416550
transform 0 -1 207593 1 0 430500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2685
timestamp 1587416550
transform 0 -1 207593 1 0 430700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2686
timestamp 1587416550
transform 0 -1 207593 1 0 430900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2688
timestamp 1587416550
transform 0 -1 207593 1 0 447100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2689
timestamp 1587416550
transform 0 -1 207593 1 0 447300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2690
timestamp 1587416550
transform 0 -1 207593 1 0 447500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2691
timestamp 1587416550
transform 0 -1 207593 1 0 447700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2693
timestamp 1587416550
transform 0 -1 207593 1 0 448100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2692
timestamp 1587416550
transform 0 -1 207593 1 0 447900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2695
timestamp 1587416550
transform 0 -1 207593 1 0 448500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2694
timestamp 1587416550
transform 0 -1 207593 1 0 448300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2697
timestamp 1587416550
transform 0 -1 207593 1 0 448900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2696
timestamp 1587416550
transform 0 -1 207593 1 0 448700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2698
timestamp 1587416550
transform 0 -1 207593 1 0 449100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2699
timestamp 1587416550
transform 0 -1 207593 1 0 449300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2700
timestamp 1587416550
transform 0 -1 207593 1 0 449500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2702
timestamp 1587416550
transform 0 -1 207593 1 0 449900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2701
timestamp 1587416550
transform 0 -1 207593 1 0 449700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2703
timestamp 1587416550
transform 0 -1 207593 1 0 450100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2704
timestamp 1587416550
transform 0 -1 207593 1 0 450300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2706
timestamp 1587416550
transform 0 -1 207593 1 0 450700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2705
timestamp 1587416550
transform 0 -1 207593 1 0 450500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2707
timestamp 1587416550
transform 0 -1 207593 1 0 450900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2708
timestamp 1587416550
transform 0 -1 207593 1 0 451100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2709
timestamp 1587416550
transform 0 -1 207593 1 0 451300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2710
timestamp 1587416550
transform 0 -1 207593 1 0 451500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2711
timestamp 1587416550
transform 0 -1 207593 1 0 451700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2712
timestamp 1587416550
transform 0 -1 207593 1 0 451900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2713
timestamp 1587416550
transform 0 -1 207593 1 0 452100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2714
timestamp 1587416550
transform 0 -1 207593 1 0 452300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2715
timestamp 1587416550
transform 0 -1 207593 1 0 452500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2716
timestamp 1587416550
transform 0 -1 207593 1 0 452700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2717
timestamp 1587416550
transform 0 -1 207593 1 0 452900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2718
timestamp 1587416550
transform 0 -1 207593 1 0 453100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2719
timestamp 1587416550
transform 0 -1 207593 1 0 453300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2720
timestamp 1587416550
transform 0 -1 207593 1 0 453500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2721
timestamp 1587416550
transform 0 -1 207593 1 0 453700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2722
timestamp 1587416550
transform 0 -1 207593 1 0 453900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2723
timestamp 1587416550
transform 0 -1 207593 1 0 454100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2724
timestamp 1587416550
transform 0 -1 207593 1 0 454300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2725
timestamp 1587416550
transform 0 -1 207593 1 0 454500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2726
timestamp 1587416550
transform 0 -1 207593 1 0 454700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2727
timestamp 1587416550
transform 0 -1 207593 1 0 454900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2728
timestamp 1587416550
transform 0 -1 207593 1 0 455100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2729
timestamp 1587416550
transform 0 -1 207593 1 0 455300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2730
timestamp 1587416550
transform 0 -1 207593 1 0 455500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2731
timestamp 1587416550
transform 0 -1 207593 1 0 455700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2732
timestamp 1587416550
transform 0 -1 207593 1 0 455900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2733
timestamp 1587416550
transform 0 -1 207593 1 0 456100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2734
timestamp 1587416550
transform 0 -1 207593 1 0 456300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2736
timestamp 1587416550
transform 0 -1 207593 1 0 456700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2735
timestamp 1587416550
transform 0 -1 207593 1 0 456500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2737
timestamp 1587416550
transform 0 -1 207593 1 0 456900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2738
timestamp 1587416550
transform 0 -1 207593 1 0 457100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2739
timestamp 1587416550
transform 0 -1 207593 1 0 457300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2740
timestamp 1587416550
transform 0 -1 207593 1 0 457500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2742
timestamp 1587416550
transform 0 -1 207593 1 0 457900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2741
timestamp 1587416550
transform 0 -1 207593 1 0 457700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2743
timestamp 1587416550
transform 0 -1 207593 1 0 458100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2744
timestamp 1587416550
transform 0 -1 207593 1 0 458300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2746
timestamp 1587416550
transform 0 -1 207593 1 0 474500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2747
timestamp 1587416550
transform 0 -1 207593 1 0 474700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2748
timestamp 1587416550
transform 0 -1 207593 1 0 474900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2749
timestamp 1587416550
transform 0 -1 207593 1 0 475100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2750
timestamp 1587416550
transform 0 -1 207593 1 0 475300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2751
timestamp 1587416550
transform 0 -1 207593 1 0 475500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2752
timestamp 1587416550
transform 0 -1 207593 1 0 475700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2753
timestamp 1587416550
transform 0 -1 207593 1 0 475900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2754
timestamp 1587416550
transform 0 -1 207593 1 0 476100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2755
timestamp 1587416550
transform 0 -1 207593 1 0 476300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2756
timestamp 1587416550
transform 0 -1 207593 1 0 476500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2757
timestamp 1587416550
transform 0 -1 207593 1 0 476700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2758
timestamp 1587416550
transform 0 -1 207593 1 0 476900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2759
timestamp 1587416550
transform 0 -1 207593 1 0 477100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2760
timestamp 1587416550
transform 0 -1 207593 1 0 477300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2761
timestamp 1587416550
transform 0 -1 207593 1 0 477500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2762
timestamp 1587416550
transform 0 -1 207593 1 0 477700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2763
timestamp 1587416550
transform 0 -1 207593 1 0 477900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2764
timestamp 1587416550
transform 0 -1 207593 1 0 478100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2766
timestamp 1587416550
transform 0 -1 207593 1 0 478500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2765
timestamp 1587416550
transform 0 -1 207593 1 0 478300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2767
timestamp 1587416550
transform 0 -1 207593 1 0 478700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2768
timestamp 1587416550
transform 0 -1 207593 1 0 478900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2770
timestamp 1587416550
transform 0 -1 207593 1 0 479300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2769
timestamp 1587416550
transform 0 -1 207593 1 0 479100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2771
timestamp 1587416550
transform 0 -1 207593 1 0 479500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2772
timestamp 1587416550
transform 0 -1 207593 1 0 479700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2773
timestamp 1587416550
transform 0 -1 207593 1 0 479900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2774
timestamp 1587416550
transform 0 -1 207593 1 0 480100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2775
timestamp 1587416550
transform 0 -1 207593 1 0 480300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2776
timestamp 1587416550
transform 0 -1 207593 1 0 480500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2777
timestamp 1587416550
transform 0 -1 207593 1 0 480700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2778
timestamp 1587416550
transform 0 -1 207593 1 0 480900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2779
timestamp 1587416550
transform 0 -1 207593 1 0 481100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2780
timestamp 1587416550
transform 0 -1 207593 1 0 481300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2781
timestamp 1587416550
transform 0 -1 207593 1 0 481500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2782
timestamp 1587416550
transform 0 -1 207593 1 0 481700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2783
timestamp 1587416550
transform 0 -1 207593 1 0 481900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2784
timestamp 1587416550
transform 0 -1 207593 1 0 482100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2785
timestamp 1587416550
transform 0 -1 207593 1 0 482300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2786
timestamp 1587416550
transform 0 -1 207593 1 0 482500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2787
timestamp 1587416550
transform 0 -1 207593 1 0 482700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2788
timestamp 1587416550
transform 0 -1 207593 1 0 482900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2789
timestamp 1587416550
transform 0 -1 207593 1 0 483100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2790
timestamp 1587416550
transform 0 -1 207593 1 0 483300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2791
timestamp 1587416550
transform 0 -1 207593 1 0 483500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2792
timestamp 1587416550
transform 0 -1 207593 1 0 483700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2793
timestamp 1587416550
transform 0 -1 207593 1 0 483900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2794
timestamp 1587416550
transform 0 -1 207593 1 0 484100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2795
timestamp 1587416550
transform 0 -1 207593 1 0 484300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2796
timestamp 1587416550
transform 0 -1 207593 1 0 484500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2797
timestamp 1587416550
transform 0 -1 207593 1 0 484700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2798
timestamp 1587416550
transform 0 -1 207593 1 0 484900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2799
timestamp 1587416550
transform 0 -1 207593 1 0 485100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2800
timestamp 1587416550
transform 0 -1 207593 1 0 485300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2801
timestamp 1587416550
transform 0 -1 207593 1 0 485500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2802
timestamp 1587416550
transform 0 -1 207593 1 0 485700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2803
timestamp 1587416550
transform 0 -1 207593 1 0 485900
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad  comp_inp_pad /usr/share/pdk/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1587416550
transform 0 -1 207593 1 0 377300
box -143 -414 16134 39593
use sky130_ef_io__gpiov2_pad  CSB_pad
timestamp 1587416550
transform 0 -1 207593 1 0 431100
box -143 -414 16134 39593
use sky130_ef_io__gpiov2_pad  SCK_pad
timestamp 1587416550
transform 0 -1 207593 1 0 458500
box -143 -414 16134 39593
use sky130_ef_io__gpiov2_pad  xclk_pad
timestamp 1587416550
transform 0 -1 207593 1 0 486100
box -143 -414 16134 39593
use striVe_soc  core
timestamp 1587660775
transform 1 0 252543 0 1 280300
box 0 0 366785 366785
use sky130_ef_io__com_bus_slice_1um  FILLER_1449
timestamp 1587416550
transform -1 0 367000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1450
timestamp 1587416550
transform -1 0 367200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1451
timestamp 1587416550
transform -1 0 367400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1452
timestamp 1587416550
transform -1 0 367600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1453
timestamp 1587416550
transform -1 0 367800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1454
timestamp 1587416550
transform -1 0 368000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1455
timestamp 1587416550
transform -1 0 368200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1456
timestamp 1587416550
transform -1 0 368400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1457
timestamp 1587416550
transform -1 0 368600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1458
timestamp 1587416550
transform -1 0 368800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1459
timestamp 1587416550
transform -1 0 369000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1460
timestamp 1587416550
transform -1 0 369200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1461
timestamp 1587416550
transform -1 0 369400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1462
timestamp 1587416550
transform -1 0 369600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1463
timestamp 1587416550
transform -1 0 369800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1464
timestamp 1587416550
transform -1 0 370000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1465
timestamp 1587416550
transform -1 0 370200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1466
timestamp 1587416550
transform -1 0 370400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1467
timestamp 1587416550
transform -1 0 370600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1468
timestamp 1587416550
transform -1 0 370800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1469
timestamp 1587416550
transform -1 0 371000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1470
timestamp 1587416550
transform -1 0 371200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1471
timestamp 1587416550
transform -1 0 371400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1472
timestamp 1587416550
transform -1 0 371600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1473
timestamp 1587416550
transform -1 0 371800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1474
timestamp 1587416550
transform -1 0 372000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1475
timestamp 1587416550
transform -1 0 372200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1476
timestamp 1587416550
transform -1 0 372400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1477
timestamp 1587416550
transform -1 0 372600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1478
timestamp 1587416550
transform -1 0 372800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1479
timestamp 1587416550
transform -1 0 373000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1480
timestamp 1587416550
transform -1 0 373200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1481
timestamp 1587416550
transform -1 0 373400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1482
timestamp 1587416550
transform -1 0 373600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1483
timestamp 1587416550
transform -1 0 373800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1484
timestamp 1587416550
transform -1 0 374000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1485
timestamp 1587416550
transform -1 0 374200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1486
timestamp 1587416550
transform -1 0 374400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1487
timestamp 1587416550
transform -1 0 374600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1488
timestamp 1587416550
transform -1 0 374800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1489
timestamp 1587416550
transform -1 0 375000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1490
timestamp 1587416550
transform -1 0 375200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1491
timestamp 1587416550
transform -1 0 375400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1492
timestamp 1587416550
transform -1 0 375600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1493
timestamp 1587416550
transform -1 0 375800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1494
timestamp 1587416550
transform -1 0 376000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1495
timestamp 1587416550
transform -1 0 376200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1496
timestamp 1587416550
transform -1 0 376400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1497
timestamp 1587416550
transform -1 0 376600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1498
timestamp 1587416550
transform -1 0 376800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1499
timestamp 1587416550
transform -1 0 377000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1500
timestamp 1587416550
transform -1 0 377200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1501
timestamp 1587416550
transform -1 0 377400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1502
timestamp 1587416550
transform -1 0 377600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1503
timestamp 1587416550
transform -1 0 377800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1504
timestamp 1587416550
transform -1 0 378000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1505
timestamp 1587416550
transform -1 0 378200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1506
timestamp 1587416550
transform -1 0 378400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1507
timestamp 1587416550
transform -1 0 378600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1508
timestamp 1587416550
transform -1 0 378800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1509
timestamp 1587416550
transform -1 0 379000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1510
timestamp 1587416550
transform -1 0 379200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1511
timestamp 1587416550
transform -1 0 379400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1512
timestamp 1587416550
transform -1 0 379600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1513
timestamp 1587416550
transform -1 0 379800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1514
timestamp 1587416550
transform -1 0 380000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1515
timestamp 1587416550
transform -1 0 380200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1516
timestamp 1587416550
transform -1 0 380400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1517
timestamp 1587416550
transform -1 0 380600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1518
timestamp 1587416550
transform -1 0 380800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1519
timestamp 1587416550
transform -1 0 381000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1520
timestamp 1587416550
transform -1 0 381200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1521
timestamp 1587416550
transform -1 0 381400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1522
timestamp 1587416550
transform -1 0 381600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1523
timestamp 1587416550
transform -1 0 381800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1524
timestamp 1587416550
transform -1 0 382000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1525
timestamp 1587416550
transform -1 0 382200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1526
timestamp 1587416550
transform -1 0 382400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1528
timestamp 1587416550
transform -1 0 398600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1530
timestamp 1587416550
transform -1 0 399000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1529
timestamp 1587416550
transform -1 0 398800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1531
timestamp 1587416550
transform -1 0 399200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1532
timestamp 1587416550
transform -1 0 399400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1534
timestamp 1587416550
transform -1 0 399800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1533
timestamp 1587416550
transform -1 0 399600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1535
timestamp 1587416550
transform -1 0 400000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1536
timestamp 1587416550
transform -1 0 400200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1537
timestamp 1587416550
transform -1 0 400400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1538
timestamp 1587416550
transform -1 0 400600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1539
timestamp 1587416550
transform -1 0 400800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1541
timestamp 1587416550
transform -1 0 401200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1540
timestamp 1587416550
transform -1 0 401000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1542
timestamp 1587416550
transform -1 0 401400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1543
timestamp 1587416550
transform -1 0 401600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1544
timestamp 1587416550
transform -1 0 401800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1545
timestamp 1587416550
transform -1 0 402000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1546
timestamp 1587416550
transform -1 0 402200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1547
timestamp 1587416550
transform -1 0 402400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1548
timestamp 1587416550
transform -1 0 402600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1549
timestamp 1587416550
transform -1 0 402800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1551
timestamp 1587416550
transform -1 0 403200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1550
timestamp 1587416550
transform -1 0 403000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1552
timestamp 1587416550
transform -1 0 403400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1553
timestamp 1587416550
transform -1 0 403600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1554
timestamp 1587416550
transform -1 0 403800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1555
timestamp 1587416550
transform -1 0 404000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1556
timestamp 1587416550
transform -1 0 404200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1557
timestamp 1587416550
transform -1 0 404400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1558
timestamp 1587416550
transform -1 0 404600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1560
timestamp 1587416550
transform -1 0 405000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1559
timestamp 1587416550
transform -1 0 404800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1562
timestamp 1587416550
transform -1 0 405400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1561
timestamp 1587416550
transform -1 0 405200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1564
timestamp 1587416550
transform -1 0 405800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1563
timestamp 1587416550
transform -1 0 405600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1566
timestamp 1587416550
transform -1 0 406200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1565
timestamp 1587416550
transform -1 0 406000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1567
timestamp 1587416550
transform -1 0 406400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1568
timestamp 1587416550
transform -1 0 406600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1569
timestamp 1587416550
transform -1 0 406800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1571
timestamp 1587416550
transform -1 0 407200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1570
timestamp 1587416550
transform -1 0 407000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1573
timestamp 1587416550
transform -1 0 407600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1572
timestamp 1587416550
transform -1 0 407400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1575
timestamp 1587416550
transform -1 0 408000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1574
timestamp 1587416550
transform -1 0 407800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1576
timestamp 1587416550
transform -1 0 408200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1577
timestamp 1587416550
transform -1 0 408400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1578
timestamp 1587416550
transform -1 0 408600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1579
timestamp 1587416550
transform -1 0 408800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1580
timestamp 1587416550
transform -1 0 409000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1581
timestamp 1587416550
transform -1 0 409200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1582
timestamp 1587416550
transform -1 0 409400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1583
timestamp 1587416550
transform -1 0 409600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1584
timestamp 1587416550
transform -1 0 409800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1585
timestamp 1587416550
transform -1 0 410000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1586
timestamp 1587416550
transform -1 0 410200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1588
timestamp 1587416550
transform -1 0 410600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1587
timestamp 1587416550
transform -1 0 410400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1589
timestamp 1587416550
transform -1 0 410800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1590
timestamp 1587416550
transform -1 0 411000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1591
timestamp 1587416550
transform -1 0 411200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1592
timestamp 1587416550
transform -1 0 411400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1593
timestamp 1587416550
transform -1 0 411600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1594
timestamp 1587416550
transform -1 0 411800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1595
timestamp 1587416550
transform -1 0 412000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1596
timestamp 1587416550
transform -1 0 412200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1597
timestamp 1587416550
transform -1 0 412400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1598
timestamp 1587416550
transform -1 0 412600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1599
timestamp 1587416550
transform -1 0 412800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1600
timestamp 1587416550
transform -1 0 413000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1601
timestamp 1587416550
transform -1 0 413200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1602
timestamp 1587416550
transform -1 0 413400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1603
timestamp 1587416550
transform -1 0 413600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1604
timestamp 1587416550
transform -1 0 413800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1605
timestamp 1587416550
transform -1 0 414000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1606
timestamp 1587416550
transform -1 0 414200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1607
timestamp 1587416550
transform -1 0 414400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1608
timestamp 1587416550
transform -1 0 414600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1609
timestamp 1587416550
transform -1 0 414800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1610
timestamp 1587416550
transform -1 0 415000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1612
timestamp 1587416550
transform -1 0 431200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1613
timestamp 1587416550
transform -1 0 431400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1614
timestamp 1587416550
transform -1 0 431600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1615
timestamp 1587416550
transform -1 0 431800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1616
timestamp 1587416550
transform -1 0 432000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1617
timestamp 1587416550
transform -1 0 432200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1618
timestamp 1587416550
transform -1 0 432400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1619
timestamp 1587416550
transform -1 0 432600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1620
timestamp 1587416550
transform -1 0 432800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1621
timestamp 1587416550
transform -1 0 433000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1622
timestamp 1587416550
transform -1 0 433200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1623
timestamp 1587416550
transform -1 0 433400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1624
timestamp 1587416550
transform -1 0 433600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1625
timestamp 1587416550
transform -1 0 433800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1626
timestamp 1587416550
transform -1 0 434000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1627
timestamp 1587416550
transform -1 0 434200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1628
timestamp 1587416550
transform -1 0 434400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1629
timestamp 1587416550
transform -1 0 434600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1630
timestamp 1587416550
transform -1 0 434800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1631
timestamp 1587416550
transform -1 0 435000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1632
timestamp 1587416550
transform -1 0 435200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1633
timestamp 1587416550
transform -1 0 435400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1634
timestamp 1587416550
transform -1 0 435600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1635
timestamp 1587416550
transform -1 0 435800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1637
timestamp 1587416550
transform -1 0 436200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1636
timestamp 1587416550
transform -1 0 436000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1638
timestamp 1587416550
transform -1 0 436400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1639
timestamp 1587416550
transform -1 0 436600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1640
timestamp 1587416550
transform -1 0 436800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1642
timestamp 1587416550
transform -1 0 437200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1641
timestamp 1587416550
transform -1 0 437000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1643
timestamp 1587416550
transform -1 0 437400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1644
timestamp 1587416550
transform -1 0 437600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1645
timestamp 1587416550
transform -1 0 437800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1646
timestamp 1587416550
transform -1 0 438000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1647
timestamp 1587416550
transform -1 0 438200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1648
timestamp 1587416550
transform -1 0 438400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1649
timestamp 1587416550
transform -1 0 438600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1650
timestamp 1587416550
transform -1 0 438800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1651
timestamp 1587416550
transform -1 0 439000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1652
timestamp 1587416550
transform -1 0 439200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1653
timestamp 1587416550
transform -1 0 439400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1654
timestamp 1587416550
transform -1 0 439600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1655
timestamp 1587416550
transform -1 0 439800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1656
timestamp 1587416550
transform -1 0 440000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1657
timestamp 1587416550
transform -1 0 440200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1658
timestamp 1587416550
transform -1 0 440400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1659
timestamp 1587416550
transform -1 0 440600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1660
timestamp 1587416550
transform -1 0 440800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1661
timestamp 1587416550
transform -1 0 441000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1662
timestamp 1587416550
transform -1 0 441200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1663
timestamp 1587416550
transform -1 0 441400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1664
timestamp 1587416550
transform -1 0 441600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1665
timestamp 1587416550
transform -1 0 441800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1666
timestamp 1587416550
transform -1 0 442000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1667
timestamp 1587416550
transform -1 0 442200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1668
timestamp 1587416550
transform -1 0 442400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1669
timestamp 1587416550
transform -1 0 442600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1670
timestamp 1587416550
transform -1 0 442800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1671
timestamp 1587416550
transform -1 0 443000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1672
timestamp 1587416550
transform -1 0 443200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1673
timestamp 1587416550
transform -1 0 443400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1674
timestamp 1587416550
transform -1 0 443600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1675
timestamp 1587416550
transform -1 0 443800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1676
timestamp 1587416550
transform -1 0 444000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1677
timestamp 1587416550
transform -1 0 444200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1678
timestamp 1587416550
transform -1 0 444400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1679
timestamp 1587416550
transform -1 0 444600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1680
timestamp 1587416550
transform -1 0 444800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1681
timestamp 1587416550
transform -1 0 445000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1682
timestamp 1587416550
transform -1 0 445200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1683
timestamp 1587416550
transform -1 0 445400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1684
timestamp 1587416550
transform -1 0 445600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1685
timestamp 1587416550
transform -1 0 445800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1686
timestamp 1587416550
transform -1 0 446000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1687
timestamp 1587416550
transform -1 0 446200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1688
timestamp 1587416550
transform -1 0 446400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1689
timestamp 1587416550
transform -1 0 446600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1690
timestamp 1587416550
transform -1 0 446800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1691
timestamp 1587416550
transform -1 0 447000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1692
timestamp 1587416550
transform -1 0 447200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1693
timestamp 1587416550
transform -1 0 447400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1696
timestamp 1587416550
transform -1 0 463800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1697
timestamp 1587416550
transform -1 0 464000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1695
timestamp 1587416550
transform -1 0 463600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1699
timestamp 1587416550
transform -1 0 464400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1700
timestamp 1587416550
transform -1 0 464600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1698
timestamp 1587416550
transform -1 0 464200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1701
timestamp 1587416550
transform -1 0 464800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1702
timestamp 1587416550
transform -1 0 465000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1703
timestamp 1587416550
transform -1 0 465200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1704
timestamp 1587416550
transform -1 0 465400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1705
timestamp 1587416550
transform -1 0 465600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1706
timestamp 1587416550
transform -1 0 465800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1707
timestamp 1587416550
transform -1 0 466000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1708
timestamp 1587416550
transform -1 0 466200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1709
timestamp 1587416550
transform -1 0 466400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1710
timestamp 1587416550
transform -1 0 466600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1711
timestamp 1587416550
transform -1 0 466800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1712
timestamp 1587416550
transform -1 0 467000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1713
timestamp 1587416550
transform -1 0 467200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1714
timestamp 1587416550
transform -1 0 467400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1715
timestamp 1587416550
transform -1 0 467600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1716
timestamp 1587416550
transform -1 0 467800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1717
timestamp 1587416550
transform -1 0 468000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1718
timestamp 1587416550
transform -1 0 468200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1719
timestamp 1587416550
transform -1 0 468400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1720
timestamp 1587416550
transform -1 0 468600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1721
timestamp 1587416550
transform -1 0 468800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1722
timestamp 1587416550
transform -1 0 469000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1723
timestamp 1587416550
transform -1 0 469200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1724
timestamp 1587416550
transform -1 0 469400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1725
timestamp 1587416550
transform -1 0 469600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1726
timestamp 1587416550
transform -1 0 469800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1727
timestamp 1587416550
transform -1 0 470000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1728
timestamp 1587416550
transform -1 0 470200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1729
timestamp 1587416550
transform -1 0 470400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1730
timestamp 1587416550
transform -1 0 470600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1731
timestamp 1587416550
transform -1 0 470800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1732
timestamp 1587416550
transform -1 0 471000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1733
timestamp 1587416550
transform -1 0 471200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1734
timestamp 1587416550
transform -1 0 471400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1735
timestamp 1587416550
transform -1 0 471600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1736
timestamp 1587416550
transform -1 0 471800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1737
timestamp 1587416550
transform -1 0 472000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1738
timestamp 1587416550
transform -1 0 472200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1739
timestamp 1587416550
transform -1 0 472400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1740
timestamp 1587416550
transform -1 0 472600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1741
timestamp 1587416550
transform -1 0 472800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1742
timestamp 1587416550
transform -1 0 473000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1743
timestamp 1587416550
transform -1 0 473200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1744
timestamp 1587416550
transform -1 0 473400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1745
timestamp 1587416550
transform -1 0 473600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1746
timestamp 1587416550
transform -1 0 473800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1747
timestamp 1587416550
transform -1 0 474000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1748
timestamp 1587416550
transform -1 0 474200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1749
timestamp 1587416550
transform -1 0 474400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1750
timestamp 1587416550
transform -1 0 474600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1751
timestamp 1587416550
transform -1 0 474800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1752
timestamp 1587416550
transform -1 0 475000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1753
timestamp 1587416550
transform -1 0 475200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1754
timestamp 1587416550
transform -1 0 475400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1755
timestamp 1587416550
transform -1 0 475600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1756
timestamp 1587416550
transform -1 0 475800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1757
timestamp 1587416550
transform -1 0 476000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1758
timestamp 1587416550
transform -1 0 476200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1759
timestamp 1587416550
transform -1 0 476400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1760
timestamp 1587416550
transform -1 0 476600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1761
timestamp 1587416550
transform -1 0 476800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1762
timestamp 1587416550
transform -1 0 477000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1763
timestamp 1587416550
transform -1 0 477200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1764
timestamp 1587416550
transform -1 0 477400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1765
timestamp 1587416550
transform -1 0 477600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1766
timestamp 1587416550
transform -1 0 477800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1767
timestamp 1587416550
transform -1 0 478000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1768
timestamp 1587416550
transform -1 0 478200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1769
timestamp 1587416550
transform -1 0 478400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1770
timestamp 1587416550
transform -1 0 478600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1771
timestamp 1587416550
transform -1 0 478800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1772
timestamp 1587416550
transform -1 0 479000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1774
timestamp 1587416550
transform -1 0 479400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1773
timestamp 1587416550
transform -1 0 479200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1775
timestamp 1587416550
transform -1 0 479600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1776
timestamp 1587416550
transform -1 0 479800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1777
timestamp 1587416550
transform -1 0 480000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1779
timestamp 1587416550
transform -1 0 496200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1780
timestamp 1587416550
transform -1 0 496400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1781
timestamp 1587416550
transform -1 0 496600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1782
timestamp 1587416550
transform -1 0 496800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1783
timestamp 1587416550
transform -1 0 497000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1784
timestamp 1587416550
transform -1 0 497200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1785
timestamp 1587416550
transform -1 0 497400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1786
timestamp 1587416550
transform -1 0 497600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1787
timestamp 1587416550
transform -1 0 497800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1788
timestamp 1587416550
transform -1 0 498000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1789
timestamp 1587416550
transform -1 0 498200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1790
timestamp 1587416550
transform -1 0 498400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1791
timestamp 1587416550
transform -1 0 498600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1792
timestamp 1587416550
transform -1 0 498800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1793
timestamp 1587416550
transform -1 0 499000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1794
timestamp 1587416550
transform -1 0 499200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1795
timestamp 1587416550
transform -1 0 499400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1796
timestamp 1587416550
transform -1 0 499600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1797
timestamp 1587416550
transform -1 0 499800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1799
timestamp 1587416550
transform -1 0 500200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1798
timestamp 1587416550
transform -1 0 500000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1800
timestamp 1587416550
transform -1 0 500400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1801
timestamp 1587416550
transform -1 0 500600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1802
timestamp 1587416550
transform -1 0 500800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1803
timestamp 1587416550
transform -1 0 501000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1804
timestamp 1587416550
transform -1 0 501200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1806
timestamp 1587416550
transform -1 0 501600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1805
timestamp 1587416550
transform -1 0 501400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1807
timestamp 1587416550
transform -1 0 501800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1808
timestamp 1587416550
transform -1 0 502000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1809
timestamp 1587416550
transform -1 0 502200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1810
timestamp 1587416550
transform -1 0 502400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1811
timestamp 1587416550
transform -1 0 502600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1812
timestamp 1587416550
transform -1 0 502800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1813
timestamp 1587416550
transform -1 0 503000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1814
timestamp 1587416550
transform -1 0 503200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1815
timestamp 1587416550
transform -1 0 503400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1816
timestamp 1587416550
transform -1 0 503600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1817
timestamp 1587416550
transform -1 0 503800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1818
timestamp 1587416550
transform -1 0 504000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1819
timestamp 1587416550
transform -1 0 504200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1820
timestamp 1587416550
transform -1 0 504400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1821
timestamp 1587416550
transform -1 0 504600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1822
timestamp 1587416550
transform -1 0 504800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1823
timestamp 1587416550
transform -1 0 505000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1825
timestamp 1587416550
transform -1 0 505400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1824
timestamp 1587416550
transform -1 0 505200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1826
timestamp 1587416550
transform -1 0 505600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1827
timestamp 1587416550
transform -1 0 505800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1828
timestamp 1587416550
transform -1 0 506000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1829
timestamp 1587416550
transform -1 0 506200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1830
timestamp 1587416550
transform -1 0 506400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1831
timestamp 1587416550
transform -1 0 506600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1832
timestamp 1587416550
transform -1 0 506800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1833
timestamp 1587416550
transform -1 0 507000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1834
timestamp 1587416550
transform -1 0 507200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1835
timestamp 1587416550
transform -1 0 507400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1836
timestamp 1587416550
transform -1 0 507600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1837
timestamp 1587416550
transform -1 0 507800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1838
timestamp 1587416550
transform -1 0 508000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1839
timestamp 1587416550
transform -1 0 508200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1840
timestamp 1587416550
transform -1 0 508400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1841
timestamp 1587416550
transform -1 0 508600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1842
timestamp 1587416550
transform -1 0 508800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1843
timestamp 1587416550
transform -1 0 509000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1844
timestamp 1587416550
transform -1 0 509200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1845
timestamp 1587416550
transform -1 0 509400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1846
timestamp 1587416550
transform -1 0 509600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1847
timestamp 1587416550
transform -1 0 509800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1848
timestamp 1587416550
transform -1 0 510000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1849
timestamp 1587416550
transform -1 0 510200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1850
timestamp 1587416550
transform -1 0 510400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1851
timestamp 1587416550
transform -1 0 510600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1852
timestamp 1587416550
transform -1 0 510800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1853
timestamp 1587416550
transform -1 0 511000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1854
timestamp 1587416550
transform -1 0 511200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1855
timestamp 1587416550
transform -1 0 511400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1856
timestamp 1587416550
transform -1 0 511600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1857
timestamp 1587416550
transform -1 0 511800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1858
timestamp 1587416550
transform -1 0 512000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1859
timestamp 1587416550
transform -1 0 512200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1860
timestamp 1587416550
transform -1 0 512400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1861
timestamp 1587416550
transform -1 0 512600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1864
timestamp 1587416550
transform -1 0 529000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1863
timestamp 1587416550
transform -1 0 528800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1867
timestamp 1587416550
transform -1 0 529600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1865
timestamp 1587416550
transform -1 0 529200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1866
timestamp 1587416550
transform -1 0 529400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1868
timestamp 1587416550
transform -1 0 529800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1869
timestamp 1587416550
transform -1 0 530000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1870
timestamp 1587416550
transform -1 0 530200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1871
timestamp 1587416550
transform -1 0 530400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1872
timestamp 1587416550
transform -1 0 530600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1873
timestamp 1587416550
transform -1 0 530800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1874
timestamp 1587416550
transform -1 0 531000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1875
timestamp 1587416550
transform -1 0 531200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1876
timestamp 1587416550
transform -1 0 531400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1877
timestamp 1587416550
transform -1 0 531600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1878
timestamp 1587416550
transform -1 0 531800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1879
timestamp 1587416550
transform -1 0 532000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1880
timestamp 1587416550
transform -1 0 532200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1881
timestamp 1587416550
transform -1 0 532400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1882
timestamp 1587416550
transform -1 0 532600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1883
timestamp 1587416550
transform -1 0 532800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1884
timestamp 1587416550
transform -1 0 533000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1885
timestamp 1587416550
transform -1 0 533200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1886
timestamp 1587416550
transform -1 0 533400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1887
timestamp 1587416550
transform -1 0 533600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1888
timestamp 1587416550
transform -1 0 533800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1889
timestamp 1587416550
transform -1 0 534000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1890
timestamp 1587416550
transform -1 0 534200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1891
timestamp 1587416550
transform -1 0 534400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1892
timestamp 1587416550
transform -1 0 534600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1893
timestamp 1587416550
transform -1 0 534800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1894
timestamp 1587416550
transform -1 0 535000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1895
timestamp 1587416550
transform -1 0 535200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1896
timestamp 1587416550
transform -1 0 535400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1897
timestamp 1587416550
transform -1 0 535600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1898
timestamp 1587416550
transform -1 0 535800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1899
timestamp 1587416550
transform -1 0 536000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1900
timestamp 1587416550
transform -1 0 536200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1901
timestamp 1587416550
transform -1 0 536400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1902
timestamp 1587416550
transform -1 0 536600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1903
timestamp 1587416550
transform -1 0 536800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1904
timestamp 1587416550
transform -1 0 537000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1905
timestamp 1587416550
transform -1 0 537200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1906
timestamp 1587416550
transform -1 0 537400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1907
timestamp 1587416550
transform -1 0 537600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1908
timestamp 1587416550
transform -1 0 537800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1909
timestamp 1587416550
transform -1 0 538000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1910
timestamp 1587416550
transform -1 0 538200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1911
timestamp 1587416550
transform -1 0 538400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1912
timestamp 1587416550
transform -1 0 538600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1913
timestamp 1587416550
transform -1 0 538800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1914
timestamp 1587416550
transform -1 0 539000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1915
timestamp 1587416550
transform -1 0 539200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1916
timestamp 1587416550
transform -1 0 539400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1917
timestamp 1587416550
transform -1 0 539600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1918
timestamp 1587416550
transform -1 0 539800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1919
timestamp 1587416550
transform -1 0 540000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1920
timestamp 1587416550
transform -1 0 540200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1921
timestamp 1587416550
transform -1 0 540400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1922
timestamp 1587416550
transform -1 0 540600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1923
timestamp 1587416550
transform -1 0 540800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1924
timestamp 1587416550
transform -1 0 541000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1925
timestamp 1587416550
transform -1 0 541200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1926
timestamp 1587416550
transform -1 0 541400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1927
timestamp 1587416550
transform -1 0 541600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1928
timestamp 1587416550
transform -1 0 541800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1929
timestamp 1587416550
transform -1 0 542000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1930
timestamp 1587416550
transform -1 0 542200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1931
timestamp 1587416550
transform -1 0 542400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1932
timestamp 1587416550
transform -1 0 542600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1933
timestamp 1587416550
transform -1 0 542800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1934
timestamp 1587416550
transform -1 0 543000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1935
timestamp 1587416550
transform -1 0 543200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1936
timestamp 1587416550
transform -1 0 543400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1937
timestamp 1587416550
transform -1 0 543600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1938
timestamp 1587416550
transform -1 0 543800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1939
timestamp 1587416550
transform -1 0 544000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1940
timestamp 1587416550
transform -1 0 544200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1941
timestamp 1587416550
transform -1 0 544400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1942
timestamp 1587416550
transform -1 0 544600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1943
timestamp 1587416550
transform -1 0 544800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1944
timestamp 1587416550
transform -1 0 545000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1945
timestamp 1587416550
transform -1 0 545200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1947
timestamp 1587416550
transform -1 0 561400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1950
timestamp 1587416550
transform -1 0 562000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1948
timestamp 1587416550
transform -1 0 561600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1949
timestamp 1587416550
transform -1 0 561800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1951
timestamp 1587416550
transform -1 0 562200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1953
timestamp 1587416550
transform -1 0 562600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1952
timestamp 1587416550
transform -1 0 562400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1954
timestamp 1587416550
transform -1 0 562800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1955
timestamp 1587416550
transform -1 0 563000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1956
timestamp 1587416550
transform -1 0 563200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1957
timestamp 1587416550
transform -1 0 563400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1959
timestamp 1587416550
transform -1 0 563800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1958
timestamp 1587416550
transform -1 0 563600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1960
timestamp 1587416550
transform -1 0 564000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1962
timestamp 1587416550
transform -1 0 564400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1961
timestamp 1587416550
transform -1 0 564200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1963
timestamp 1587416550
transform -1 0 564600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1964
timestamp 1587416550
transform -1 0 564800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1966
timestamp 1587416550
transform -1 0 565200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1965
timestamp 1587416550
transform -1 0 565000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1967
timestamp 1587416550
transform -1 0 565400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1968
timestamp 1587416550
transform -1 0 565600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1969
timestamp 1587416550
transform -1 0 565800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1970
timestamp 1587416550
transform -1 0 566000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1972
timestamp 1587416550
transform -1 0 566400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1971
timestamp 1587416550
transform -1 0 566200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1973
timestamp 1587416550
transform -1 0 566600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1974
timestamp 1587416550
transform -1 0 566800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1975
timestamp 1587416550
transform -1 0 567000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1976
timestamp 1587416550
transform -1 0 567200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1977
timestamp 1587416550
transform -1 0 567400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1978
timestamp 1587416550
transform -1 0 567600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1979
timestamp 1587416550
transform -1 0 567800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1981
timestamp 1587416550
transform -1 0 568200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1980
timestamp 1587416550
transform -1 0 568000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1983
timestamp 1587416550
transform -1 0 568600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1982
timestamp 1587416550
transform -1 0 568400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1985
timestamp 1587416550
transform -1 0 569000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1984
timestamp 1587416550
transform -1 0 568800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1987
timestamp 1587416550
transform -1 0 569400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1986
timestamp 1587416550
transform -1 0 569200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1988
timestamp 1587416550
transform -1 0 569600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1989
timestamp 1587416550
transform -1 0 569800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1990
timestamp 1587416550
transform -1 0 570000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1992
timestamp 1587416550
transform -1 0 570400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1991
timestamp 1587416550
transform -1 0 570200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1994
timestamp 1587416550
transform -1 0 570800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1993
timestamp 1587416550
transform -1 0 570600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1996
timestamp 1587416550
transform -1 0 571200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1995
timestamp 1587416550
transform -1 0 571000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1997
timestamp 1587416550
transform -1 0 571400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1998
timestamp 1587416550
transform -1 0 571600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1999
timestamp 1587416550
transform -1 0 571800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2000
timestamp 1587416550
transform -1 0 572000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2001
timestamp 1587416550
transform -1 0 572200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2002
timestamp 1587416550
transform -1 0 572400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2003
timestamp 1587416550
transform -1 0 572600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2004
timestamp 1587416550
transform -1 0 572800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2005
timestamp 1587416550
transform -1 0 573000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2006
timestamp 1587416550
transform -1 0 573200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2007
timestamp 1587416550
transform -1 0 573400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2008
timestamp 1587416550
transform -1 0 573600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2009
timestamp 1587416550
transform -1 0 573800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2010
timestamp 1587416550
transform -1 0 574000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2011
timestamp 1587416550
transform -1 0 574200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2012
timestamp 1587416550
transform -1 0 574400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2013
timestamp 1587416550
transform -1 0 574600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2014
timestamp 1587416550
transform -1 0 574800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2015
timestamp 1587416550
transform -1 0 575000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2016
timestamp 1587416550
transform -1 0 575200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2017
timestamp 1587416550
transform -1 0 575400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2018
timestamp 1587416550
transform -1 0 575600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2019
timestamp 1587416550
transform -1 0 575800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2020
timestamp 1587416550
transform -1 0 576000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2021
timestamp 1587416550
transform -1 0 576200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2022
timestamp 1587416550
transform -1 0 576400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2023
timestamp 1587416550
transform -1 0 576600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2024
timestamp 1587416550
transform -1 0 576800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2025
timestamp 1587416550
transform -1 0 577000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2026
timestamp 1587416550
transform -1 0 577200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2027
timestamp 1587416550
transform -1 0 577400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2028
timestamp 1587416550
transform -1 0 577600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2029
timestamp 1587416550
transform -1 0 577800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2031
timestamp 1587416550
transform -1 0 594000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2032
timestamp 1587416550
transform -1 0 594200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2034
timestamp 1587416550
transform -1 0 594600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2033
timestamp 1587416550
transform -1 0 594400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2035
timestamp 1587416550
transform -1 0 594800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2036
timestamp 1587416550
transform -1 0 595000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2037
timestamp 1587416550
transform -1 0 595200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2038
timestamp 1587416550
transform -1 0 595400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2039
timestamp 1587416550
transform -1 0 595600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2040
timestamp 1587416550
transform -1 0 595800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2041
timestamp 1587416550
transform -1 0 596000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2042
timestamp 1587416550
transform -1 0 596200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2043
timestamp 1587416550
transform -1 0 596400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2044
timestamp 1587416550
transform -1 0 596600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2045
timestamp 1587416550
transform -1 0 596800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2046
timestamp 1587416550
transform -1 0 597000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2047
timestamp 1587416550
transform -1 0 597200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2048
timestamp 1587416550
transform -1 0 597400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2049
timestamp 1587416550
transform -1 0 597600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2050
timestamp 1587416550
transform -1 0 597800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2052
timestamp 1587416550
transform -1 0 598200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2051
timestamp 1587416550
transform -1 0 598000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2053
timestamp 1587416550
transform -1 0 598400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2054
timestamp 1587416550
transform -1 0 598600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2055
timestamp 1587416550
transform -1 0 598800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2056
timestamp 1587416550
transform -1 0 599000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2057
timestamp 1587416550
transform -1 0 599200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2058
timestamp 1587416550
transform -1 0 599400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2059
timestamp 1587416550
transform -1 0 599600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2060
timestamp 1587416550
transform -1 0 599800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2061
timestamp 1587416550
transform -1 0 600000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2062
timestamp 1587416550
transform -1 0 600200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2063
timestamp 1587416550
transform -1 0 600400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2064
timestamp 1587416550
transform -1 0 600600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2065
timestamp 1587416550
transform -1 0 600800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2066
timestamp 1587416550
transform -1 0 601000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2067
timestamp 1587416550
transform -1 0 601200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2068
timestamp 1587416550
transform -1 0 601400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2069
timestamp 1587416550
transform -1 0 601600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2070
timestamp 1587416550
transform -1 0 601800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2071
timestamp 1587416550
transform -1 0 602000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2072
timestamp 1587416550
transform -1 0 602200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2073
timestamp 1587416550
transform -1 0 602400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2074
timestamp 1587416550
transform -1 0 602600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2075
timestamp 1587416550
transform -1 0 602800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2076
timestamp 1587416550
transform -1 0 603000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2077
timestamp 1587416550
transform -1 0 603200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2078
timestamp 1587416550
transform -1 0 603400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2079
timestamp 1587416550
transform -1 0 603600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2080
timestamp 1587416550
transform -1 0 603800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2081
timestamp 1587416550
transform -1 0 604000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2082
timestamp 1587416550
transform -1 0 604200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2083
timestamp 1587416550
transform -1 0 604400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2084
timestamp 1587416550
transform -1 0 604600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2085
timestamp 1587416550
transform -1 0 604800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2086
timestamp 1587416550
transform -1 0 605000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2087
timestamp 1587416550
transform -1 0 605200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2088
timestamp 1587416550
transform -1 0 605400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2089
timestamp 1587416550
transform -1 0 605600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2090
timestamp 1587416550
transform -1 0 605800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2091
timestamp 1587416550
transform -1 0 606000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2092
timestamp 1587416550
transform -1 0 606200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2093
timestamp 1587416550
transform -1 0 606400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2095
timestamp 1587416550
transform -1 0 606800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2094
timestamp 1587416550
transform -1 0 606600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2096
timestamp 1587416550
transform -1 0 607000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2097
timestamp 1587416550
transform -1 0 607200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2098
timestamp 1587416550
transform -1 0 607400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2099
timestamp 1587416550
transform -1 0 607600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2100
timestamp 1587416550
transform -1 0 607800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2101
timestamp 1587416550
transform -1 0 608000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2102
timestamp 1587416550
transform -1 0 608200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2103
timestamp 1587416550
transform -1 0 608400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2104
timestamp 1587416550
transform -1 0 608600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2105
timestamp 1587416550
transform -1 0 608800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2106
timestamp 1587416550
transform -1 0 609000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2107
timestamp 1587416550
transform -1 0 609200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2108
timestamp 1587416550
transform -1 0 609400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2109
timestamp 1587416550
transform -1 0 609600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2110
timestamp 1587416550
transform -1 0 609800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2111
timestamp 1587416550
transform -1 0 610000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2112
timestamp 1587416550
transform -1 0 610200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2113
timestamp 1587416550
transform -1 0 610400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2115
timestamp 1587416550
transform -1 0 626600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2116
timestamp 1587416550
transform -1 0 626800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2118
timestamp 1587416550
transform -1 0 627200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2119
timestamp 1587416550
transform -1 0 627400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2117
timestamp 1587416550
transform -1 0 627000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2121
timestamp 1587416550
transform -1 0 627800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2120
timestamp 1587416550
transform -1 0 627600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2122
timestamp 1587416550
transform -1 0 628000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2123
timestamp 1587416550
transform -1 0 628200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2124
timestamp 1587416550
transform -1 0 628400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2125
timestamp 1587416550
transform -1 0 628600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2126
timestamp 1587416550
transform -1 0 628800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2127
timestamp 1587416550
transform -1 0 629000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2128
timestamp 1587416550
transform -1 0 629200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2129
timestamp 1587416550
transform -1 0 629400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2130
timestamp 1587416550
transform -1 0 629600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2131
timestamp 1587416550
transform -1 0 629800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2132
timestamp 1587416550
transform -1 0 630000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2133
timestamp 1587416550
transform -1 0 630200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2134
timestamp 1587416550
transform -1 0 630400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2135
timestamp 1587416550
transform -1 0 630600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2136
timestamp 1587416550
transform -1 0 630800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2137
timestamp 1587416550
transform -1 0 631000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2138
timestamp 1587416550
transform -1 0 631200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2139
timestamp 1587416550
transform -1 0 631400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2140
timestamp 1587416550
transform -1 0 631600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2141
timestamp 1587416550
transform -1 0 631800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2142
timestamp 1587416550
transform -1 0 632000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2143
timestamp 1587416550
transform -1 0 632200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2144
timestamp 1587416550
transform -1 0 632400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2145
timestamp 1587416550
transform -1 0 632600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2146
timestamp 1587416550
transform -1 0 632800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2147
timestamp 1587416550
transform -1 0 633000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2148
timestamp 1587416550
transform -1 0 633200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2149
timestamp 1587416550
transform -1 0 633400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2150
timestamp 1587416550
transform -1 0 633600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2151
timestamp 1587416550
transform -1 0 633800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2152
timestamp 1587416550
transform -1 0 634000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2153
timestamp 1587416550
transform -1 0 634200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2154
timestamp 1587416550
transform -1 0 634400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2155
timestamp 1587416550
transform -1 0 634600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2156
timestamp 1587416550
transform -1 0 634800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2157
timestamp 1587416550
transform -1 0 635000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2158
timestamp 1587416550
transform -1 0 635200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2159
timestamp 1587416550
transform -1 0 635400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2160
timestamp 1587416550
transform -1 0 635600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2161
timestamp 1587416550
transform -1 0 635800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2162
timestamp 1587416550
transform -1 0 636000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2163
timestamp 1587416550
transform -1 0 636200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2164
timestamp 1587416550
transform -1 0 636400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2165
timestamp 1587416550
transform -1 0 636600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2166
timestamp 1587416550
transform -1 0 636800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2167
timestamp 1587416550
transform -1 0 637000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2168
timestamp 1587416550
transform -1 0 637200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2169
timestamp 1587416550
transform -1 0 637400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2170
timestamp 1587416550
transform -1 0 637600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2171
timestamp 1587416550
transform -1 0 637800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2172
timestamp 1587416550
transform -1 0 638000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2173
timestamp 1587416550
transform -1 0 638200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2174
timestamp 1587416550
transform -1 0 638400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2175
timestamp 1587416550
transform -1 0 638600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2176
timestamp 1587416550
transform -1 0 638800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2177
timestamp 1587416550
transform -1 0 639000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2178
timestamp 1587416550
transform -1 0 639200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2179
timestamp 1587416550
transform -1 0 639400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2180
timestamp 1587416550
transform -1 0 639600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2181
timestamp 1587416550
transform -1 0 639800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2182
timestamp 1587416550
transform -1 0 640000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2183
timestamp 1587416550
transform -1 0 640200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2184
timestamp 1587416550
transform -1 0 640400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2185
timestamp 1587416550
transform -1 0 640600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2186
timestamp 1587416550
transform -1 0 640800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2187
timestamp 1587416550
transform -1 0 641000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2188
timestamp 1587416550
transform -1 0 641200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2189
timestamp 1587416550
transform -1 0 641400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2190
timestamp 1587416550
transform -1 0 641600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2191
timestamp 1587416550
transform -1 0 641800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2192
timestamp 1587416550
transform -1 0 642000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2193
timestamp 1587416550
transform -1 0 642200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2194
timestamp 1587416550
transform -1 0 642400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2195
timestamp 1587416550
transform -1 0 642600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2196
timestamp 1587416550
transform -1 0 642800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2197
timestamp 1587416550
transform -1 0 643000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2199
timestamp 1587416550
transform -1 0 659200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2200
timestamp 1587416550
transform -1 0 659400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2201
timestamp 1587416550
transform -1 0 659600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2202
timestamp 1587416550
transform -1 0 659800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2204
timestamp 1587416550
transform -1 0 660200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2203
timestamp 1587416550
transform -1 0 660000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2205
timestamp 1587416550
transform -1 0 660400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2206
timestamp 1587416550
transform -1 0 660600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2207
timestamp 1587416550
transform -1 0 660800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2208
timestamp 1587416550
transform -1 0 661000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2209
timestamp 1587416550
transform -1 0 661200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2210
timestamp 1587416550
transform -1 0 661400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2211
timestamp 1587416550
transform -1 0 661600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2212
timestamp 1587416550
transform -1 0 661800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2213
timestamp 1587416550
transform -1 0 662000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2214
timestamp 1587416550
transform -1 0 662200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2215
timestamp 1587416550
transform -1 0 662400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2216
timestamp 1587416550
transform -1 0 662600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2217
timestamp 1587416550
transform -1 0 662800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2218
timestamp 1587416550
transform -1 0 663000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2219
timestamp 1587416550
transform -1 0 663200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2220
timestamp 1587416550
transform -1 0 663400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2221
timestamp 1587416550
transform -1 0 663600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2222
timestamp 1587416550
transform -1 0 663800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2223
timestamp 1587416550
transform -1 0 664000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2224
timestamp 1587416550
transform -1 0 664200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2225
timestamp 1587416550
transform -1 0 664400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2226
timestamp 1587416550
transform -1 0 664600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2227
timestamp 1587416550
transform -1 0 664800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2228
timestamp 1587416550
transform -1 0 665000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2229
timestamp 1587416550
transform -1 0 665200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2230
timestamp 1587416550
transform -1 0 665400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2231
timestamp 1587416550
transform -1 0 665600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2232
timestamp 1587416550
transform -1 0 665800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2233
timestamp 1587416550
transform -1 0 666000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2234
timestamp 1587416550
transform -1 0 666200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2235
timestamp 1587416550
transform -1 0 666400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2236
timestamp 1587416550
transform -1 0 666600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2237
timestamp 1587416550
transform -1 0 666800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2238
timestamp 1587416550
transform -1 0 667000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2239
timestamp 1587416550
transform -1 0 667200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2240
timestamp 1587416550
transform -1 0 667400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2241
timestamp 1587416550
transform -1 0 667600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2242
timestamp 1587416550
transform -1 0 667800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2243
timestamp 1587416550
transform -1 0 668000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2244
timestamp 1587416550
transform -1 0 668200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2245
timestamp 1587416550
transform -1 0 668400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2247
timestamp 1587416550
transform -1 0 668800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2246
timestamp 1587416550
transform -1 0 668600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2248
timestamp 1587416550
transform -1 0 669000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2249
timestamp 1587416550
transform -1 0 669200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2250
timestamp 1587416550
transform -1 0 669400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2251
timestamp 1587416550
transform -1 0 669600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2252
timestamp 1587416550
transform -1 0 669800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2253
timestamp 1587416550
transform -1 0 670000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2254
timestamp 1587416550
transform -1 0 670200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2255
timestamp 1587416550
transform -1 0 670400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2256
timestamp 1587416550
transform -1 0 670600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2257
timestamp 1587416550
transform -1 0 670800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2258
timestamp 1587416550
transform -1 0 671000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2259
timestamp 1587416550
transform -1 0 671200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2260
timestamp 1587416550
transform -1 0 671400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2261
timestamp 1587416550
transform -1 0 671600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2263
timestamp 1587416550
transform -1 0 672000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2262
timestamp 1587416550
transform -1 0 671800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2264
timestamp 1587416550
transform -1 0 672200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2265
timestamp 1587416550
transform -1 0 672400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2266
timestamp 1587416550
transform -1 0 672600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2267
timestamp 1587416550
transform -1 0 672800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2269
timestamp 1587416550
transform -1 0 673200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2268
timestamp 1587416550
transform -1 0 673000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2270
timestamp 1587416550
transform -1 0 673400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2271
timestamp 1587416550
transform -1 0 673600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2272
timestamp 1587416550
transform -1 0 673800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2274
timestamp 1587416550
transform -1 0 674200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2273
timestamp 1587416550
transform -1 0 674000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2275
timestamp 1587416550
transform -1 0 674400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2276
timestamp 1587416550
transform -1 0 674600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2277
timestamp 1587416550
transform -1 0 674800 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2278
timestamp 1587416550
transform -1 0 675000 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2280
timestamp 1587416550
transform -1 0 675400 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2279
timestamp 1587416550
transform -1 0 675200 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2281
timestamp 1587416550
transform -1 0 675600 0 -1 259093
box 0 0 200 39593
use sky130_ef_io__corner_pad  corner[0]
timestamp 1587416550
transform 0 1 675600 -1 0 259500
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_1um  FILLER_3269
timestamp 1587416550
transform 0 1 676807 -1 0 259700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3270
timestamp 1587416550
transform 0 1 676807 -1 0 259900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3271
timestamp 1587416550
transform 0 1 676807 -1 0 260100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3272
timestamp 1587416550
transform 0 1 676807 -1 0 260300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3273
timestamp 1587416550
transform 0 1 676807 -1 0 260500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3274
timestamp 1587416550
transform 0 1 676807 -1 0 260700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3275
timestamp 1587416550
transform 0 1 676807 -1 0 260900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3276
timestamp 1587416550
transform 0 1 676807 -1 0 261100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3277
timestamp 1587416550
transform 0 1 676807 -1 0 261300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3278
timestamp 1587416550
transform 0 1 676807 -1 0 261500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3279
timestamp 1587416550
transform 0 1 676807 -1 0 261700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3280
timestamp 1587416550
transform 0 1 676807 -1 0 261900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3281
timestamp 1587416550
transform 0 1 676807 -1 0 262100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3282
timestamp 1587416550
transform 0 1 676807 -1 0 262300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3283
timestamp 1587416550
transform 0 1 676807 -1 0 262500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3284
timestamp 1587416550
transform 0 1 676807 -1 0 262700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3285
timestamp 1587416550
transform 0 1 676807 -1 0 262900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3286
timestamp 1587416550
transform 0 1 676807 -1 0 263100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3287
timestamp 1587416550
transform 0 1 676807 -1 0 263300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3288
timestamp 1587416550
transform 0 1 676807 -1 0 263500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3289
timestamp 1587416550
transform 0 1 676807 -1 0 263700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3290
timestamp 1587416550
transform 0 1 676807 -1 0 263900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3291
timestamp 1587416550
transform 0 1 676807 -1 0 264100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3292
timestamp 1587416550
transform 0 1 676807 -1 0 264300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3293
timestamp 1587416550
transform 0 1 676807 -1 0 264500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3294
timestamp 1587416550
transform 0 1 676807 -1 0 264700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3295
timestamp 1587416550
transform 0 1 676807 -1 0 264900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3296
timestamp 1587416550
transform 0 1 676807 -1 0 265100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3297
timestamp 1587416550
transform 0 1 676807 -1 0 265300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3298
timestamp 1587416550
transform 0 1 676807 -1 0 265500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3299
timestamp 1587416550
transform 0 1 676807 -1 0 265700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3300
timestamp 1587416550
transform 0 1 676807 -1 0 265900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3301
timestamp 1587416550
transform 0 1 676807 -1 0 266100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3302
timestamp 1587416550
transform 0 1 676807 -1 0 266300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3303
timestamp 1587416550
transform 0 1 676807 -1 0 266500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3304
timestamp 1587416550
transform 0 1 676807 -1 0 266700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3305
timestamp 1587416550
transform 0 1 676807 -1 0 266900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3306
timestamp 1587416550
transform 0 1 676807 -1 0 267100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3307
timestamp 1587416550
transform 0 1 676807 -1 0 267300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3308
timestamp 1587416550
transform 0 1 676807 -1 0 267500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3309
timestamp 1587416550
transform 0 1 676807 -1 0 267700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3310
timestamp 1587416550
transform 0 1 676807 -1 0 267900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3311
timestamp 1587416550
transform 0 1 676807 -1 0 268100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3312
timestamp 1587416550
transform 0 1 676807 -1 0 268300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3313
timestamp 1587416550
transform 0 1 676807 -1 0 268500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3314
timestamp 1587416550
transform 0 1 676807 -1 0 268700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3315
timestamp 1587416550
transform 0 1 676807 -1 0 268900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3316
timestamp 1587416550
transform 0 1 676807 -1 0 269100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3317
timestamp 1587416550
transform 0 1 676807 -1 0 269300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3318
timestamp 1587416550
transform 0 1 676807 -1 0 269500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3319
timestamp 1587416550
transform 0 1 676807 -1 0 269700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3320
timestamp 1587416550
transform 0 1 676807 -1 0 269900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3321
timestamp 1587416550
transform 0 1 676807 -1 0 270100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3322
timestamp 1587416550
transform 0 1 676807 -1 0 270300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3323
timestamp 1587416550
transform 0 1 676807 -1 0 270500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3324
timestamp 1587416550
transform 0 1 676807 -1 0 270700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3325
timestamp 1587416550
transform 0 1 676807 -1 0 270900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3326
timestamp 1587416550
transform 0 1 676807 -1 0 271100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3327
timestamp 1587416550
transform 0 1 676807 -1 0 271300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3328
timestamp 1587416550
transform 0 1 676807 -1 0 271500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3329
timestamp 1587416550
transform 0 1 676807 -1 0 271700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3330
timestamp 1587416550
transform 0 1 676807 -1 0 271900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3331
timestamp 1587416550
transform 0 1 676807 -1 0 272100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3332
timestamp 1587416550
transform 0 1 676807 -1 0 272300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3333
timestamp 1587416550
transform 0 1 676807 -1 0 272500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3334
timestamp 1587416550
transform 0 1 676807 -1 0 272700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3335
timestamp 1587416550
transform 0 1 676807 -1 0 272900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3336
timestamp 1587416550
transform 0 1 676807 -1 0 273100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3337
timestamp 1587416550
transform 0 1 676807 -1 0 273300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3338
timestamp 1587416550
transform 0 1 676807 -1 0 273500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3339
timestamp 1587416550
transform 0 1 676807 -1 0 273700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3340
timestamp 1587416550
transform 0 1 676807 -1 0 273900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3341
timestamp 1587416550
transform 0 1 676807 -1 0 274100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3342
timestamp 1587416550
transform 0 1 676807 -1 0 274300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3343
timestamp 1587416550
transform 0 1 676807 -1 0 274500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3344
timestamp 1587416550
transform 0 1 676807 -1 0 274700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3345
timestamp 1587416550
transform 0 1 676807 -1 0 274900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3346
timestamp 1587416550
transform 0 1 676807 -1 0 275100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3347
timestamp 1587416550
transform 0 1 676807 -1 0 275300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3348
timestamp 1587416550
transform 0 1 676807 -1 0 275500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3349
timestamp 1587416550
transform 0 1 676807 -1 0 275700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3350
timestamp 1587416550
transform 0 1 676807 -1 0 275900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3351
timestamp 1587416550
transform 0 1 676807 -1 0 276100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3352
timestamp 1587416550
transform 0 1 676807 -1 0 276300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3353
timestamp 1587416550
transform 0 1 676807 -1 0 276500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3354
timestamp 1587416550
transform 0 1 676807 -1 0 276700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3355
timestamp 1587416550
transform 0 1 676807 -1 0 276900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3356
timestamp 1587416550
transform 0 1 676807 -1 0 277100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3357
timestamp 1587416550
transform 0 1 676807 -1 0 277300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3358
timestamp 1587416550
transform 0 1 676807 -1 0 277500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3359
timestamp 1587416550
transform 0 1 676807 -1 0 277700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3360
timestamp 1587416550
transform 0 1 676807 -1 0 277900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3361
timestamp 1587416550
transform 0 1 676807 -1 0 278100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3362
timestamp 1587416550
transform 0 1 676807 -1 0 278300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3363
timestamp 1587416550
transform 0 1 676807 -1 0 278500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3364
timestamp 1587416550
transform 0 1 676807 -1 0 278700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3365
timestamp 1587416550
transform 0 1 676807 -1 0 278900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3366
timestamp 1587416550
transform 0 1 676807 -1 0 279100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3367
timestamp 1587416550
transform 0 1 676807 -1 0 279300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3368
timestamp 1587416550
transform 0 1 676807 -1 0 279500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3369
timestamp 1587416550
transform 0 1 676807 -1 0 279700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3370
timestamp 1587416550
transform 0 1 676807 -1 0 279900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3371
timestamp 1587416550
transform 0 1 676807 -1 0 280100
box 0 0 200 39593
use sky130_fd_sc_hd__conb_1  mask_rev_value[0] /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1587416520
transform 1 0 639328 0 1 280300
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1587416520
transform 1 0 639604 0 1 280300
box -38 -48 130 592
use sky130_ef_io__com_bus_slice_1um  FILLER_3372
timestamp 1587416550
transform 0 1 676807 -1 0 280300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3373
timestamp 1587416550
transform 0 1 676807 -1 0 280500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3374
timestamp 1587416550
transform 0 1 676807 -1 0 280700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3375
timestamp 1587416550
transform 0 1 676807 -1 0 280900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3376
timestamp 1587416550
transform 0 1 676807 -1 0 281100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3377
timestamp 1587416550
transform 0 1 676807 -1 0 281300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3378
timestamp 1587416550
transform 0 1 676807 -1 0 281500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3379
timestamp 1587416550
transform 0 1 676807 -1 0 281700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3380
timestamp 1587416550
transform 0 1 676807 -1 0 281900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3382
timestamp 1587416550
transform 0 1 676807 -1 0 282300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3381
timestamp 1587416550
transform 0 1 676807 -1 0 282100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3383
timestamp 1587416550
transform 0 1 676807 -1 0 282500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3384
timestamp 1587416550
transform 0 1 676807 -1 0 282700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3385
timestamp 1587416550
transform 0 1 676807 -1 0 282900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3386
timestamp 1587416550
transform 0 1 676807 -1 0 283100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3387
timestamp 1587416550
transform 0 1 676807 -1 0 283300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3388
timestamp 1587416550
transform 0 1 676807 -1 0 283500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3389
timestamp 1587416550
transform 0 1 676807 -1 0 283700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3390
timestamp 1587416550
transform 0 1 676807 -1 0 283900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3391
timestamp 1587416550
transform 0 1 676807 -1 0 284100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3392
timestamp 1587416550
transform 0 1 676807 -1 0 284300
box 0 0 200 39593
use sky130_ef_io__vdda_hvc_pad  vdd3v3hclamp[1]
timestamp 1587416550
transform 0 1 676807 -1 0 299300
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3394
timestamp 1587416550
transform 0 1 676807 -1 0 299500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3395
timestamp 1587416550
transform 0 1 676807 -1 0 299700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3396
timestamp 1587416550
transform 0 1 676807 -1 0 299900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3397
timestamp 1587416550
transform 0 1 676807 -1 0 300100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3398
timestamp 1587416550
transform 0 1 676807 -1 0 300300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3399
timestamp 1587416550
transform 0 1 676807 -1 0 300500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3400
timestamp 1587416550
transform 0 1 676807 -1 0 300700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3401
timestamp 1587416550
transform 0 1 676807 -1 0 300900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3402
timestamp 1587416550
transform 0 1 676807 -1 0 301100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3403
timestamp 1587416550
transform 0 1 676807 -1 0 301300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3404
timestamp 1587416550
transform 0 1 676807 -1 0 301500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3405
timestamp 1587416550
transform 0 1 676807 -1 0 301700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3406
timestamp 1587416550
transform 0 1 676807 -1 0 301900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3407
timestamp 1587416550
transform 0 1 676807 -1 0 302100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3408
timestamp 1587416550
transform 0 1 676807 -1 0 302300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3409
timestamp 1587416550
transform 0 1 676807 -1 0 302500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3410
timestamp 1587416550
transform 0 1 676807 -1 0 302700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3411
timestamp 1587416550
transform 0 1 676807 -1 0 302900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3412
timestamp 1587416550
transform 0 1 676807 -1 0 303100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3413
timestamp 1587416550
transform 0 1 676807 -1 0 303300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3414
timestamp 1587416550
transform 0 1 676807 -1 0 303500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3415
timestamp 1587416550
transform 0 1 676807 -1 0 303700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3416
timestamp 1587416550
transform 0 1 676807 -1 0 303900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3417
timestamp 1587416550
transform 0 1 676807 -1 0 304100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3418
timestamp 1587416550
transform 0 1 676807 -1 0 304300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3419
timestamp 1587416550
transform 0 1 676807 -1 0 304500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3420
timestamp 1587416550
transform 0 1 676807 -1 0 304700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3421
timestamp 1587416550
transform 0 1 676807 -1 0 304900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3422
timestamp 1587416550
transform 0 1 676807 -1 0 305100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3423
timestamp 1587416550
transform 0 1 676807 -1 0 305300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3424
timestamp 1587416550
transform 0 1 676807 -1 0 305500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3425
timestamp 1587416550
transform 0 1 676807 -1 0 305700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3426
timestamp 1587416550
transform 0 1 676807 -1 0 305900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3427
timestamp 1587416550
transform 0 1 676807 -1 0 306100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3428
timestamp 1587416550
transform 0 1 676807 -1 0 306300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3429
timestamp 1587416550
transform 0 1 676807 -1 0 306500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3430
timestamp 1587416550
transform 0 1 676807 -1 0 306700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3431
timestamp 1587416550
transform 0 1 676807 -1 0 306900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3432
timestamp 1587416550
transform 0 1 676807 -1 0 307100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3433
timestamp 1587416550
transform 0 1 676807 -1 0 307300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3434
timestamp 1587416550
transform 0 1 676807 -1 0 307500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3435
timestamp 1587416550
transform 0 1 676807 -1 0 307700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3436
timestamp 1587416550
transform 0 1 676807 -1 0 307900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3437
timestamp 1587416550
transform 0 1 676807 -1 0 308100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3438
timestamp 1587416550
transform 0 1 676807 -1 0 308300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3439
timestamp 1587416550
transform 0 1 676807 -1 0 308500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3440
timestamp 1587416550
transform 0 1 676807 -1 0 308700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3441
timestamp 1587416550
transform 0 1 676807 -1 0 308900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3442
timestamp 1587416550
transform 0 1 676807 -1 0 309100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3443
timestamp 1587416550
transform 0 1 676807 -1 0 309300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3444
timestamp 1587416550
transform 0 1 676807 -1 0 309500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3445
timestamp 1587416550
transform 0 1 676807 -1 0 309700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3446
timestamp 1587416550
transform 0 1 676807 -1 0 309900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3447
timestamp 1587416550
transform 0 1 676807 -1 0 310100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3448
timestamp 1587416550
transform 0 1 676807 -1 0 310300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3449
timestamp 1587416550
transform 0 1 676807 -1 0 310500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3450
timestamp 1587416550
transform 0 1 676807 -1 0 310700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3451
timestamp 1587416550
transform 0 1 676807 -1 0 310900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3452
timestamp 1587416550
transform 0 1 676807 -1 0 311100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3453
timestamp 1587416550
transform 0 1 676807 -1 0 311300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3454
timestamp 1587416550
transform 0 1 676807 -1 0 311500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3455
timestamp 1587416550
transform 0 1 676807 -1 0 311700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3456
timestamp 1587416550
transform 0 1 676807 -1 0 311900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3457
timestamp 1587416550
transform 0 1 676807 -1 0 312100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3458
timestamp 1587416550
transform 0 1 676807 -1 0 312300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3459
timestamp 1587416550
transform 0 1 676807 -1 0 312500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3460
timestamp 1587416550
transform 0 1 676807 -1 0 312700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3461
timestamp 1587416550
transform 0 1 676807 -1 0 312900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3462
timestamp 1587416550
transform 0 1 676807 -1 0 313100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3463
timestamp 1587416550
transform 0 1 676807 -1 0 313300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3464
timestamp 1587416550
transform 0 1 676807 -1 0 313500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3465
timestamp 1587416550
transform 0 1 676807 -1 0 313700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3466
timestamp 1587416550
transform 0 1 676807 -1 0 313900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3467
timestamp 1587416550
transform 0 1 676807 -1 0 314100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3468
timestamp 1587416550
transform 0 1 676807 -1 0 314300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3469
timestamp 1587416550
transform 0 1 676807 -1 0 314500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3470
timestamp 1587416550
transform 0 1 676807 -1 0 314700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3471
timestamp 1587416550
transform 0 1 676807 -1 0 314900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3472
timestamp 1587416550
transform 0 1 676807 -1 0 315100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3473
timestamp 1587416550
transform 0 1 676807 -1 0 315300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3474
timestamp 1587416550
transform 0 1 676807 -1 0 315500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3475
timestamp 1587416550
transform 0 1 676807 -1 0 315700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3476
timestamp 1587416550
transform 0 1 676807 -1 0 315900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3477
timestamp 1587416550
transform 0 1 676807 -1 0 316100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3478
timestamp 1587416550
transform 0 1 676807 -1 0 316300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3479
timestamp 1587416550
transform 0 1 676807 -1 0 316500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3480
timestamp 1587416550
transform 0 1 676807 -1 0 316700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3481
timestamp 1587416550
transform 0 1 676807 -1 0 316900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3482
timestamp 1587416550
transform 0 1 676807 -1 0 317100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3483
timestamp 1587416550
transform 0 1 676807 -1 0 317300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3484
timestamp 1587416550
transform 0 1 676807 -1 0 317500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3485
timestamp 1587416550
transform 0 1 676807 -1 0 317700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3486
timestamp 1587416550
transform 0 1 676807 -1 0 317900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3487
timestamp 1587416550
transform 0 1 676807 -1 0 318100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3488
timestamp 1587416550
transform 0 1 676807 -1 0 318300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3489
timestamp 1587416550
transform 0 1 676807 -1 0 318500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3490
timestamp 1587416550
transform 0 1 676807 -1 0 318700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3491
timestamp 1587416550
transform 0 1 676807 -1 0 318900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3492
timestamp 1587416550
transform 0 1 676807 -1 0 319100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3493
timestamp 1587416550
transform 0 1 676807 -1 0 319300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3494
timestamp 1587416550
transform 0 1 676807 -1 0 319500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3495
timestamp 1587416550
transform 0 1 676807 -1 0 319700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3496
timestamp 1587416550
transform 0 1 676807 -1 0 319900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3497
timestamp 1587416550
transform 0 1 676807 -1 0 320100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3498
timestamp 1587416550
transform 0 1 676807 -1 0 320300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3499
timestamp 1587416550
transform 0 1 676807 -1 0 320500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3500
timestamp 1587416550
transform 0 1 676807 -1 0 320700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3501
timestamp 1587416550
transform 0 1 676807 -1 0 320900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3502
timestamp 1587416550
transform 0 1 676807 -1 0 321100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3503
timestamp 1587416550
transform 0 1 676807 -1 0 321300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3504
timestamp 1587416550
transform 0 1 676807 -1 0 321500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3505
timestamp 1587416550
transform 0 1 676807 -1 0 321700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3506
timestamp 1587416550
transform 0 1 676807 -1 0 321900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3507
timestamp 1587416550
transform 0 1 676807 -1 0 322100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3508
timestamp 1587416550
transform 0 1 676807 -1 0 322300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3509
timestamp 1587416550
transform 0 1 676807 -1 0 322500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3510
timestamp 1587416550
transform 0 1 676807 -1 0 322700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3511
timestamp 1587416550
transform 0 1 676807 -1 0 322900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3512
timestamp 1587416550
transform 0 1 676807 -1 0 323100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3513
timestamp 1587416550
transform 0 1 676807 -1 0 323300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3514
timestamp 1587416550
transform 0 1 676807 -1 0 323500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3515
timestamp 1587416550
transform 0 1 676807 -1 0 323700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3516
timestamp 1587416550
transform 0 1 676807 -1 0 323900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3517
timestamp 1587416550
transform 0 1 676807 -1 0 324100
box 0 0 200 39593
use sky130_ef_io__vdda_lvc_pad  vdd3v3lclamp[1]
timestamp 1587416550
transform 0 1 676807 -1 0 339100
box 0 -7 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3519
timestamp 1587416550
transform 0 1 676807 -1 0 339300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3520
timestamp 1587416550
transform 0 1 676807 -1 0 339500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3521
timestamp 1587416550
transform 0 1 676807 -1 0 339700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3523
timestamp 1587416550
transform 0 1 676807 -1 0 340100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3522
timestamp 1587416550
transform 0 1 676807 -1 0 339900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3524
timestamp 1587416550
transform 0 1 676807 -1 0 340300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3525
timestamp 1587416550
transform 0 1 676807 -1 0 340500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3526
timestamp 1587416550
transform 0 1 676807 -1 0 340700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3527
timestamp 1587416550
transform 0 1 676807 -1 0 340900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3528
timestamp 1587416550
transform 0 1 676807 -1 0 341100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3529
timestamp 1587416550
transform 0 1 676807 -1 0 341300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3530
timestamp 1587416550
transform 0 1 676807 -1 0 341500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3531
timestamp 1587416550
transform 0 1 676807 -1 0 341700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3532
timestamp 1587416550
transform 0 1 676807 -1 0 341900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3533
timestamp 1587416550
transform 0 1 676807 -1 0 342100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3534
timestamp 1587416550
transform 0 1 676807 -1 0 342300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3535
timestamp 1587416550
transform 0 1 676807 -1 0 342500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3536
timestamp 1587416550
transform 0 1 676807 -1 0 342700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3537
timestamp 1587416550
transform 0 1 676807 -1 0 342900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3538
timestamp 1587416550
transform 0 1 676807 -1 0 343100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3539
timestamp 1587416550
transform 0 1 676807 -1 0 343300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3540
timestamp 1587416550
transform 0 1 676807 -1 0 343500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3541
timestamp 1587416550
transform 0 1 676807 -1 0 343700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3542
timestamp 1587416550
transform 0 1 676807 -1 0 343900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3543
timestamp 1587416550
transform 0 1 676807 -1 0 344100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3544
timestamp 1587416550
transform 0 1 676807 -1 0 344300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3545
timestamp 1587416550
transform 0 1 676807 -1 0 344500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3546
timestamp 1587416550
transform 0 1 676807 -1 0 344700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3547
timestamp 1587416550
transform 0 1 676807 -1 0 344900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3548
timestamp 1587416550
transform 0 1 676807 -1 0 345100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3549
timestamp 1587416550
transform 0 1 676807 -1 0 345300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3550
timestamp 1587416550
transform 0 1 676807 -1 0 345500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3551
timestamp 1587416550
transform 0 1 676807 -1 0 345700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3552
timestamp 1587416550
transform 0 1 676807 -1 0 345900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3553
timestamp 1587416550
transform 0 1 676807 -1 0 346100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3554
timestamp 1587416550
transform 0 1 676807 -1 0 346300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3555
timestamp 1587416550
transform 0 1 676807 -1 0 346500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3556
timestamp 1587416550
transform 0 1 676807 -1 0 346700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3557
timestamp 1587416550
transform 0 1 676807 -1 0 346900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3558
timestamp 1587416550
transform 0 1 676807 -1 0 347100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3559
timestamp 1587416550
transform 0 1 676807 -1 0 347300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3560
timestamp 1587416550
transform 0 1 676807 -1 0 347500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3561
timestamp 1587416550
transform 0 1 676807 -1 0 347700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3562
timestamp 1587416550
transform 0 1 676807 -1 0 347900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3563
timestamp 1587416550
transform 0 1 676807 -1 0 348100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3564
timestamp 1587416550
transform 0 1 676807 -1 0 348300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3565
timestamp 1587416550
transform 0 1 676807 -1 0 348500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3566
timestamp 1587416550
transform 0 1 676807 -1 0 348700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3567
timestamp 1587416550
transform 0 1 676807 -1 0 348900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3568
timestamp 1587416550
transform 0 1 676807 -1 0 349100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3569
timestamp 1587416550
transform 0 1 676807 -1 0 349300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3570
timestamp 1587416550
transform 0 1 676807 -1 0 349500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3571
timestamp 1587416550
transform 0 1 676807 -1 0 349700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3572
timestamp 1587416550
transform 0 1 676807 -1 0 349900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3573
timestamp 1587416550
transform 0 1 676807 -1 0 350100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3574
timestamp 1587416550
transform 0 1 676807 -1 0 350300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3575
timestamp 1587416550
transform 0 1 676807 -1 0 350500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3576
timestamp 1587416550
transform 0 1 676807 -1 0 350700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3577
timestamp 1587416550
transform 0 1 676807 -1 0 350900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3578
timestamp 1587416550
transform 0 1 676807 -1 0 351100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3579
timestamp 1587416550
transform 0 1 676807 -1 0 351300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3580
timestamp 1587416550
transform 0 1 676807 -1 0 351500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3581
timestamp 1587416550
transform 0 1 676807 -1 0 351700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3582
timestamp 1587416550
transform 0 1 676807 -1 0 351900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3583
timestamp 1587416550
transform 0 1 676807 -1 0 352100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3584
timestamp 1587416550
transform 0 1 676807 -1 0 352300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3585
timestamp 1587416550
transform 0 1 676807 -1 0 352500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3586
timestamp 1587416550
transform 0 1 676807 -1 0 352700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3587
timestamp 1587416550
transform 0 1 676807 -1 0 352900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3588
timestamp 1587416550
transform 0 1 676807 -1 0 353100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3589
timestamp 1587416550
transform 0 1 676807 -1 0 353300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3590
timestamp 1587416550
transform 0 1 676807 -1 0 353500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3591
timestamp 1587416550
transform 0 1 676807 -1 0 353700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3592
timestamp 1587416550
transform 0 1 676807 -1 0 353900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3593
timestamp 1587416550
transform 0 1 676807 -1 0 354100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3594
timestamp 1587416550
transform 0 1 676807 -1 0 354300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3595
timestamp 1587416550
transform 0 1 676807 -1 0 354500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3596
timestamp 1587416550
transform 0 1 676807 -1 0 354700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3597
timestamp 1587416550
transform 0 1 676807 -1 0 354900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3598
timestamp 1587416550
transform 0 1 676807 -1 0 355100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3599
timestamp 1587416550
transform 0 1 676807 -1 0 355300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3600
timestamp 1587416550
transform 0 1 676807 -1 0 355500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3601
timestamp 1587416550
transform 0 1 676807 -1 0 355700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3602
timestamp 1587416550
transform 0 1 676807 -1 0 355900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3603
timestamp 1587416550
transform 0 1 676807 -1 0 356100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3604
timestamp 1587416550
transform 0 1 676807 -1 0 356300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3605
timestamp 1587416550
transform 0 1 676807 -1 0 356500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3606
timestamp 1587416550
transform 0 1 676807 -1 0 356700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3607
timestamp 1587416550
transform 0 1 676807 -1 0 356900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3608
timestamp 1587416550
transform 0 1 676807 -1 0 357100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3609
timestamp 1587416550
transform 0 1 676807 -1 0 357300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3610
timestamp 1587416550
transform 0 1 676807 -1 0 357500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3611
timestamp 1587416550
transform 0 1 676807 -1 0 357700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3612
timestamp 1587416550
transform 0 1 676807 -1 0 357900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3613
timestamp 1587416550
transform 0 1 676807 -1 0 358100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3614
timestamp 1587416550
transform 0 1 676807 -1 0 358300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3615
timestamp 1587416550
transform 0 1 676807 -1 0 358500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3616
timestamp 1587416550
transform 0 1 676807 -1 0 358700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3617
timestamp 1587416550
transform 0 1 676807 -1 0 358900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3618
timestamp 1587416550
transform 0 1 676807 -1 0 359100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3619
timestamp 1587416550
transform 0 1 676807 -1 0 359300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3620
timestamp 1587416550
transform 0 1 676807 -1 0 359500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3621
timestamp 1587416550
transform 0 1 676807 -1 0 359700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3622
timestamp 1587416550
transform 0 1 676807 -1 0 359900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3623
timestamp 1587416550
transform 0 1 676807 -1 0 360100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3624
timestamp 1587416550
transform 0 1 676807 -1 0 360300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3625
timestamp 1587416550
transform 0 1 676807 -1 0 360500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3626
timestamp 1587416550
transform 0 1 676807 -1 0 360700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3627
timestamp 1587416550
transform 0 1 676807 -1 0 360900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3628
timestamp 1587416550
transform 0 1 676807 -1 0 361100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3629
timestamp 1587416550
transform 0 1 676807 -1 0 361300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3630
timestamp 1587416550
transform 0 1 676807 -1 0 361500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3631
timestamp 1587416550
transform 0 1 676807 -1 0 361700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3632
timestamp 1587416550
transform 0 1 676807 -1 0 361900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3633
timestamp 1587416550
transform 0 1 676807 -1 0 362100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3634
timestamp 1587416550
transform 0 1 676807 -1 0 362300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3635
timestamp 1587416550
transform 0 1 676807 -1 0 362500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3636
timestamp 1587416550
transform 0 1 676807 -1 0 362700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3637
timestamp 1587416550
transform 0 1 676807 -1 0 362900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3638
timestamp 1587416550
transform 0 1 676807 -1 0 363100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3639
timestamp 1587416550
transform 0 1 676807 -1 0 363300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3640
timestamp 1587416550
transform 0 1 676807 -1 0 363500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3641
timestamp 1587416550
transform 0 1 676807 -1 0 363700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3642
timestamp 1587416550
transform 0 1 676807 -1 0 363900
box 0 0 200 39593
use sky130_ef_io__vccd_hvc_pad  vdd1v8hclamp[1] /usr/share/pdk/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1587416550
transform 0 1 676807 -1 0 378900
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3644
timestamp 1587416550
transform 0 1 676807 -1 0 379100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3645
timestamp 1587416550
transform 0 1 676807 -1 0 379300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3646
timestamp 1587416550
transform 0 1 676807 -1 0 379500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3647
timestamp 1587416550
transform 0 1 676807 -1 0 379700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3648
timestamp 1587416550
transform 0 1 676807 -1 0 379900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3649
timestamp 1587416550
transform 0 1 676807 -1 0 380100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3650
timestamp 1587416550
transform 0 1 676807 -1 0 380300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3651
timestamp 1587416550
transform 0 1 676807 -1 0 380500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3652
timestamp 1587416550
transform 0 1 676807 -1 0 380700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3653
timestamp 1587416550
transform 0 1 676807 -1 0 380900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3654
timestamp 1587416550
transform 0 1 676807 -1 0 381100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3655
timestamp 1587416550
transform 0 1 676807 -1 0 381300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3656
timestamp 1587416550
transform 0 1 676807 -1 0 381500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3657
timestamp 1587416550
transform 0 1 676807 -1 0 381700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3658
timestamp 1587416550
transform 0 1 676807 -1 0 381900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3659
timestamp 1587416550
transform 0 1 676807 -1 0 382100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3660
timestamp 1587416550
transform 0 1 676807 -1 0 382300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3661
timestamp 1587416550
transform 0 1 676807 -1 0 382500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3662
timestamp 1587416550
transform 0 1 676807 -1 0 382700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3663
timestamp 1587416550
transform 0 1 676807 -1 0 382900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3664
timestamp 1587416550
transform 0 1 676807 -1 0 383100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3665
timestamp 1587416550
transform 0 1 676807 -1 0 383300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3666
timestamp 1587416550
transform 0 1 676807 -1 0 383500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3667
timestamp 1587416550
transform 0 1 676807 -1 0 383700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3668
timestamp 1587416550
transform 0 1 676807 -1 0 383900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3669
timestamp 1587416550
transform 0 1 676807 -1 0 384100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3670
timestamp 1587416550
transform 0 1 676807 -1 0 384300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3671
timestamp 1587416550
transform 0 1 676807 -1 0 384500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3672
timestamp 1587416550
transform 0 1 676807 -1 0 384700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3673
timestamp 1587416550
transform 0 1 676807 -1 0 384900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3674
timestamp 1587416550
transform 0 1 676807 -1 0 385100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3675
timestamp 1587416550
transform 0 1 676807 -1 0 385300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3676
timestamp 1587416550
transform 0 1 676807 -1 0 385500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3677
timestamp 1587416550
transform 0 1 676807 -1 0 385700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3678
timestamp 1587416550
transform 0 1 676807 -1 0 385900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3679
timestamp 1587416550
transform 0 1 676807 -1 0 386100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3680
timestamp 1587416550
transform 0 1 676807 -1 0 386300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3681
timestamp 1587416550
transform 0 1 676807 -1 0 386500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3682
timestamp 1587416550
transform 0 1 676807 -1 0 386700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3683
timestamp 1587416550
transform 0 1 676807 -1 0 386900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3684
timestamp 1587416550
transform 0 1 676807 -1 0 387100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3685
timestamp 1587416550
transform 0 1 676807 -1 0 387300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3686
timestamp 1587416550
transform 0 1 676807 -1 0 387500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3687
timestamp 1587416550
transform 0 1 676807 -1 0 387700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3688
timestamp 1587416550
transform 0 1 676807 -1 0 387900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3689
timestamp 1587416550
transform 0 1 676807 -1 0 388100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3690
timestamp 1587416550
transform 0 1 676807 -1 0 388300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3691
timestamp 1587416550
transform 0 1 676807 -1 0 388500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3692
timestamp 1587416550
transform 0 1 676807 -1 0 388700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3693
timestamp 1587416550
transform 0 1 676807 -1 0 388900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3694
timestamp 1587416550
transform 0 1 676807 -1 0 389100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3695
timestamp 1587416550
transform 0 1 676807 -1 0 389300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3696
timestamp 1587416550
transform 0 1 676807 -1 0 389500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3697
timestamp 1587416550
transform 0 1 676807 -1 0 389700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3698
timestamp 1587416550
transform 0 1 676807 -1 0 389900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3699
timestamp 1587416550
transform 0 1 676807 -1 0 390100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3700
timestamp 1587416550
transform 0 1 676807 -1 0 390300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3701
timestamp 1587416550
transform 0 1 676807 -1 0 390500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3702
timestamp 1587416550
transform 0 1 676807 -1 0 390700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3703
timestamp 1587416550
transform 0 1 676807 -1 0 390900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3704
timestamp 1587416550
transform 0 1 676807 -1 0 391100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3705
timestamp 1587416550
transform 0 1 676807 -1 0 391300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3706
timestamp 1587416550
transform 0 1 676807 -1 0 391500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3707
timestamp 1587416550
transform 0 1 676807 -1 0 391700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3708
timestamp 1587416550
transform 0 1 676807 -1 0 391900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3709
timestamp 1587416550
transform 0 1 676807 -1 0 392100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3710
timestamp 1587416550
transform 0 1 676807 -1 0 392300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3711
timestamp 1587416550
transform 0 1 676807 -1 0 392500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3712
timestamp 1587416550
transform 0 1 676807 -1 0 392700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3713
timestamp 1587416550
transform 0 1 676807 -1 0 392900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3714
timestamp 1587416550
transform 0 1 676807 -1 0 393100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3715
timestamp 1587416550
transform 0 1 676807 -1 0 393300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3716
timestamp 1587416550
transform 0 1 676807 -1 0 393500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3717
timestamp 1587416550
transform 0 1 676807 -1 0 393700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3718
timestamp 1587416550
transform 0 1 676807 -1 0 393900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3719
timestamp 1587416550
transform 0 1 676807 -1 0 394100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3720
timestamp 1587416550
transform 0 1 676807 -1 0 394300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3721
timestamp 1587416550
transform 0 1 676807 -1 0 394500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3722
timestamp 1587416550
transform 0 1 676807 -1 0 394700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3723
timestamp 1587416550
transform 0 1 676807 -1 0 394900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3724
timestamp 1587416550
transform 0 1 676807 -1 0 395100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3725
timestamp 1587416550
transform 0 1 676807 -1 0 395300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3726
timestamp 1587416550
transform 0 1 676807 -1 0 395500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3727
timestamp 1587416550
transform 0 1 676807 -1 0 395700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3728
timestamp 1587416550
transform 0 1 676807 -1 0 395900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3729
timestamp 1587416550
transform 0 1 676807 -1 0 396100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3730
timestamp 1587416550
transform 0 1 676807 -1 0 396300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3731
timestamp 1587416550
transform 0 1 676807 -1 0 396500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3732
timestamp 1587416550
transform 0 1 676807 -1 0 396700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3733
timestamp 1587416550
transform 0 1 676807 -1 0 396900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3734
timestamp 1587416550
transform 0 1 676807 -1 0 397100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3735
timestamp 1587416550
transform 0 1 676807 -1 0 397300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3736
timestamp 1587416550
transform 0 1 676807 -1 0 397500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3737
timestamp 1587416550
transform 0 1 676807 -1 0 397700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3738
timestamp 1587416550
transform 0 1 676807 -1 0 397900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3739
timestamp 1587416550
transform 0 1 676807 -1 0 398100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3740
timestamp 1587416550
transform 0 1 676807 -1 0 398300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3741
timestamp 1587416550
transform 0 1 676807 -1 0 398500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3742
timestamp 1587416550
transform 0 1 676807 -1 0 398700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3743
timestamp 1587416550
transform 0 1 676807 -1 0 398900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3744
timestamp 1587416550
transform 0 1 676807 -1 0 399100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3745
timestamp 1587416550
transform 0 1 676807 -1 0 399300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3746
timestamp 1587416550
transform 0 1 676807 -1 0 399500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3747
timestamp 1587416550
transform 0 1 676807 -1 0 399700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3748
timestamp 1587416550
transform 0 1 676807 -1 0 399900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3749
timestamp 1587416550
transform 0 1 676807 -1 0 400100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3750
timestamp 1587416550
transform 0 1 676807 -1 0 400300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3751
timestamp 1587416550
transform 0 1 676807 -1 0 400500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3752
timestamp 1587416550
transform 0 1 676807 -1 0 400700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3753
timestamp 1587416550
transform 0 1 676807 -1 0 400900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3754
timestamp 1587416550
transform 0 1 676807 -1 0 401100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3755
timestamp 1587416550
transform 0 1 676807 -1 0 401300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3756
timestamp 1587416550
transform 0 1 676807 -1 0 401500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3757
timestamp 1587416550
transform 0 1 676807 -1 0 401700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3758
timestamp 1587416550
transform 0 1 676807 -1 0 401900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3759
timestamp 1587416550
transform 0 1 676807 -1 0 402100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3760
timestamp 1587416550
transform 0 1 676807 -1 0 402300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3761
timestamp 1587416550
transform 0 1 676807 -1 0 402500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3762
timestamp 1587416550
transform 0 1 676807 -1 0 402700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3763
timestamp 1587416550
transform 0 1 676807 -1 0 402900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3764
timestamp 1587416550
transform 0 1 676807 -1 0 403100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3765
timestamp 1587416550
transform 0 1 676807 -1 0 403300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3766
timestamp 1587416550
transform 0 1 676807 -1 0 403500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3767
timestamp 1587416550
transform 0 1 676807 -1 0 403700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3768
timestamp 1587416550
transform 0 1 676807 -1 0 403900
box 0 0 200 39593
use sky130_ef_io__vssa_hvc_pad  vsshclamp[3]
timestamp 1587416550
transform 0 1 676807 -1 0 418900
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3770
timestamp 1587416550
transform 0 1 676807 -1 0 419100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3771
timestamp 1587416550
transform 0 1 676807 -1 0 419300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3773
timestamp 1587416550
transform 0 1 676807 -1 0 419700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3772
timestamp 1587416550
transform 0 1 676807 -1 0 419500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3774
timestamp 1587416550
transform 0 1 676807 -1 0 419900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3775
timestamp 1587416550
transform 0 1 676807 -1 0 420100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3776
timestamp 1587416550
transform 0 1 676807 -1 0 420300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3777
timestamp 1587416550
transform 0 1 676807 -1 0 420500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3778
timestamp 1587416550
transform 0 1 676807 -1 0 420700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3779
timestamp 1587416550
transform 0 1 676807 -1 0 420900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3781
timestamp 1587416550
transform 0 1 676807 -1 0 421300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3780
timestamp 1587416550
transform 0 1 676807 -1 0 421100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3782
timestamp 1587416550
transform 0 1 676807 -1 0 421500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3783
timestamp 1587416550
transform 0 1 676807 -1 0 421700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3785
timestamp 1587416550
transform 0 1 676807 -1 0 422100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3784
timestamp 1587416550
transform 0 1 676807 -1 0 421900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3786
timestamp 1587416550
transform 0 1 676807 -1 0 422300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3787
timestamp 1587416550
transform 0 1 676807 -1 0 422500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3788
timestamp 1587416550
transform 0 1 676807 -1 0 422700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3789
timestamp 1587416550
transform 0 1 676807 -1 0 422900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3790
timestamp 1587416550
transform 0 1 676807 -1 0 423100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3791
timestamp 1587416550
transform 0 1 676807 -1 0 423300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3792
timestamp 1587416550
transform 0 1 676807 -1 0 423500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3793
timestamp 1587416550
transform 0 1 676807 -1 0 423700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3794
timestamp 1587416550
transform 0 1 676807 -1 0 423900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3795
timestamp 1587416550
transform 0 1 676807 -1 0 424100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3796
timestamp 1587416550
transform 0 1 676807 -1 0 424300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3797
timestamp 1587416550
transform 0 1 676807 -1 0 424500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3798
timestamp 1587416550
transform 0 1 676807 -1 0 424700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3799
timestamp 1587416550
transform 0 1 676807 -1 0 424900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3800
timestamp 1587416550
transform 0 1 676807 -1 0 425100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3801
timestamp 1587416550
transform 0 1 676807 -1 0 425300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3802
timestamp 1587416550
transform 0 1 676807 -1 0 425500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3803
timestamp 1587416550
transform 0 1 676807 -1 0 425700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3804
timestamp 1587416550
transform 0 1 676807 -1 0 425900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3805
timestamp 1587416550
transform 0 1 676807 -1 0 426100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3806
timestamp 1587416550
transform 0 1 676807 -1 0 426300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3807
timestamp 1587416550
transform 0 1 676807 -1 0 426500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3808
timestamp 1587416550
transform 0 1 676807 -1 0 426700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3809
timestamp 1587416550
transform 0 1 676807 -1 0 426900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3810
timestamp 1587416550
transform 0 1 676807 -1 0 427100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3811
timestamp 1587416550
transform 0 1 676807 -1 0 427300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3812
timestamp 1587416550
transform 0 1 676807 -1 0 427500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3813
timestamp 1587416550
transform 0 1 676807 -1 0 427700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3814
timestamp 1587416550
transform 0 1 676807 -1 0 427900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3815
timestamp 1587416550
transform 0 1 676807 -1 0 428100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3816
timestamp 1587416550
transform 0 1 676807 -1 0 428300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3817
timestamp 1587416550
transform 0 1 676807 -1 0 428500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3818
timestamp 1587416550
transform 0 1 676807 -1 0 428700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3819
timestamp 1587416550
transform 0 1 676807 -1 0 428900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3820
timestamp 1587416550
transform 0 1 676807 -1 0 429100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3821
timestamp 1587416550
transform 0 1 676807 -1 0 429300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3822
timestamp 1587416550
transform 0 1 676807 -1 0 429500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3823
timestamp 1587416550
transform 0 1 676807 -1 0 429700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3824
timestamp 1587416550
transform 0 1 676807 -1 0 429900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3825
timestamp 1587416550
transform 0 1 676807 -1 0 430100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3826
timestamp 1587416550
transform 0 1 676807 -1 0 430300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3827
timestamp 1587416550
transform 0 1 676807 -1 0 430500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3828
timestamp 1587416550
transform 0 1 676807 -1 0 430700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3829
timestamp 1587416550
transform 0 1 676807 -1 0 430900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3830
timestamp 1587416550
transform 0 1 676807 -1 0 431100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3831
timestamp 1587416550
transform 0 1 676807 -1 0 431300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3832
timestamp 1587416550
transform 0 1 676807 -1 0 431500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3833
timestamp 1587416550
transform 0 1 676807 -1 0 431700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3834
timestamp 1587416550
transform 0 1 676807 -1 0 431900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3835
timestamp 1587416550
transform 0 1 676807 -1 0 432100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3836
timestamp 1587416550
transform 0 1 676807 -1 0 432300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3837
timestamp 1587416550
transform 0 1 676807 -1 0 432500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3838
timestamp 1587416550
transform 0 1 676807 -1 0 432700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3839
timestamp 1587416550
transform 0 1 676807 -1 0 432900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3840
timestamp 1587416550
transform 0 1 676807 -1 0 433100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3841
timestamp 1587416550
transform 0 1 676807 -1 0 433300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3842
timestamp 1587416550
transform 0 1 676807 -1 0 433500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3843
timestamp 1587416550
transform 0 1 676807 -1 0 433700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3844
timestamp 1587416550
transform 0 1 676807 -1 0 433900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3845
timestamp 1587416550
transform 0 1 676807 -1 0 434100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3846
timestamp 1587416550
transform 0 1 676807 -1 0 434300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3847
timestamp 1587416550
transform 0 1 676807 -1 0 434500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3848
timestamp 1587416550
transform 0 1 676807 -1 0 434700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3849
timestamp 1587416550
transform 0 1 676807 -1 0 434900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3850
timestamp 1587416550
transform 0 1 676807 -1 0 435100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3851
timestamp 1587416550
transform 0 1 676807 -1 0 435300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3852
timestamp 1587416550
transform 0 1 676807 -1 0 435500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3853
timestamp 1587416550
transform 0 1 676807 -1 0 435700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3854
timestamp 1587416550
transform 0 1 676807 -1 0 435900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3855
timestamp 1587416550
transform 0 1 676807 -1 0 436100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3856
timestamp 1587416550
transform 0 1 676807 -1 0 436300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3857
timestamp 1587416550
transform 0 1 676807 -1 0 436500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3858
timestamp 1587416550
transform 0 1 676807 -1 0 436700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3859
timestamp 1587416550
transform 0 1 676807 -1 0 436900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3860
timestamp 1587416550
transform 0 1 676807 -1 0 437100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3861
timestamp 1587416550
transform 0 1 676807 -1 0 437300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3862
timestamp 1587416550
transform 0 1 676807 -1 0 437500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3863
timestamp 1587416550
transform 0 1 676807 -1 0 437700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3864
timestamp 1587416550
transform 0 1 676807 -1 0 437900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3865
timestamp 1587416550
transform 0 1 676807 -1 0 438100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3866
timestamp 1587416550
transform 0 1 676807 -1 0 438300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3867
timestamp 1587416550
transform 0 1 676807 -1 0 438500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3868
timestamp 1587416550
transform 0 1 676807 -1 0 438700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3869
timestamp 1587416550
transform 0 1 676807 -1 0 438900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3870
timestamp 1587416550
transform 0 1 676807 -1 0 439100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3871
timestamp 1587416550
transform 0 1 676807 -1 0 439300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3872
timestamp 1587416550
transform 0 1 676807 -1 0 439500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3873
timestamp 1587416550
transform 0 1 676807 -1 0 439700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3874
timestamp 1587416550
transform 0 1 676807 -1 0 439900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3875
timestamp 1587416550
transform 0 1 676807 -1 0 440100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3876
timestamp 1587416550
transform 0 1 676807 -1 0 440300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3877
timestamp 1587416550
transform 0 1 676807 -1 0 440500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3878
timestamp 1587416550
transform 0 1 676807 -1 0 440700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3879
timestamp 1587416550
transform 0 1 676807 -1 0 440900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3880
timestamp 1587416550
transform 0 1 676807 -1 0 441100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3881
timestamp 1587416550
transform 0 1 676807 -1 0 441300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3882
timestamp 1587416550
transform 0 1 676807 -1 0 441500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3883
timestamp 1587416550
transform 0 1 676807 -1 0 441700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3884
timestamp 1587416550
transform 0 1 676807 -1 0 441900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3885
timestamp 1587416550
transform 0 1 676807 -1 0 442100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3886
timestamp 1587416550
transform 0 1 676807 -1 0 442300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3887
timestamp 1587416550
transform 0 1 676807 -1 0 442500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3888
timestamp 1587416550
transform 0 1 676807 -1 0 442700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3889
timestamp 1587416550
transform 0 1 676807 -1 0 442900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3890
timestamp 1587416550
transform 0 1 676807 -1 0 443100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3891
timestamp 1587416550
transform 0 1 676807 -1 0 443300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3892
timestamp 1587416550
transform 0 1 676807 -1 0 443500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3893
timestamp 1587416550
transform 0 1 676807 -1 0 443700
box 0 0 200 39593
use sky130_ef_io__vssa_lvc_pad  sky130_ef_io__vssa_lvc_pad_0 /usr/share/pdk/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1587416550
transform 0 1 676807 -1 0 458700
box 0 -7 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3895
timestamp 1587416550
transform 0 1 676807 -1 0 458900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3896
timestamp 1587416550
transform 0 1 676807 -1 0 459100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3897
timestamp 1587416550
transform 0 1 676807 -1 0 459300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3898
timestamp 1587416550
transform 0 1 676807 -1 0 459500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3900
timestamp 1587416550
transform 0 1 676807 -1 0 459900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3899
timestamp 1587416550
transform 0 1 676807 -1 0 459700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3901
timestamp 1587416550
transform 0 1 676807 -1 0 460100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3902
timestamp 1587416550
transform 0 1 676807 -1 0 460300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3904
timestamp 1587416550
transform 0 1 676807 -1 0 460700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3903
timestamp 1587416550
transform 0 1 676807 -1 0 460500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3905
timestamp 1587416550
transform 0 1 676807 -1 0 460900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3906
timestamp 1587416550
transform 0 1 676807 -1 0 461100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3907
timestamp 1587416550
transform 0 1 676807 -1 0 461300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3908
timestamp 1587416550
transform 0 1 676807 -1 0 461500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3909
timestamp 1587416550
transform 0 1 676807 -1 0 461700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3910
timestamp 1587416550
transform 0 1 676807 -1 0 461900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3912
timestamp 1587416550
transform 0 1 676807 -1 0 462300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3911
timestamp 1587416550
transform 0 1 676807 -1 0 462100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3913
timestamp 1587416550
transform 0 1 676807 -1 0 462500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3914
timestamp 1587416550
transform 0 1 676807 -1 0 462700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3916
timestamp 1587416550
transform 0 1 676807 -1 0 463100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3915
timestamp 1587416550
transform 0 1 676807 -1 0 462900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3917
timestamp 1587416550
transform 0 1 676807 -1 0 463300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3918
timestamp 1587416550
transform 0 1 676807 -1 0 463500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3919
timestamp 1587416550
transform 0 1 676807 -1 0 463700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3920
timestamp 1587416550
transform 0 1 676807 -1 0 463900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3921
timestamp 1587416550
transform 0 1 676807 -1 0 464100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3922
timestamp 1587416550
transform 0 1 676807 -1 0 464300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3923
timestamp 1587416550
transform 0 1 676807 -1 0 464500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3924
timestamp 1587416550
transform 0 1 676807 -1 0 464700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3925
timestamp 1587416550
transform 0 1 676807 -1 0 464900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3926
timestamp 1587416550
transform 0 1 676807 -1 0 465100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3927
timestamp 1587416550
transform 0 1 676807 -1 0 465300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3928
timestamp 1587416550
transform 0 1 676807 -1 0 465500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3929
timestamp 1587416550
transform 0 1 676807 -1 0 465700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3930
timestamp 1587416550
transform 0 1 676807 -1 0 465900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3931
timestamp 1587416550
transform 0 1 676807 -1 0 466100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3932
timestamp 1587416550
transform 0 1 676807 -1 0 466300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3933
timestamp 1587416550
transform 0 1 676807 -1 0 466500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3934
timestamp 1587416550
transform 0 1 676807 -1 0 466700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3935
timestamp 1587416550
transform 0 1 676807 -1 0 466900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3936
timestamp 1587416550
transform 0 1 676807 -1 0 467100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3937
timestamp 1587416550
transform 0 1 676807 -1 0 467300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3938
timestamp 1587416550
transform 0 1 676807 -1 0 467500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3939
timestamp 1587416550
transform 0 1 676807 -1 0 467700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3940
timestamp 1587416550
transform 0 1 676807 -1 0 467900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3941
timestamp 1587416550
transform 0 1 676807 -1 0 468100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3942
timestamp 1587416550
transform 0 1 676807 -1 0 468300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3943
timestamp 1587416550
transform 0 1 676807 -1 0 468500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3944
timestamp 1587416550
transform 0 1 676807 -1 0 468700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3945
timestamp 1587416550
transform 0 1 676807 -1 0 468900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3946
timestamp 1587416550
transform 0 1 676807 -1 0 469100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3947
timestamp 1587416550
transform 0 1 676807 -1 0 469300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3948
timestamp 1587416550
transform 0 1 676807 -1 0 469500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3949
timestamp 1587416550
transform 0 1 676807 -1 0 469700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3950
timestamp 1587416550
transform 0 1 676807 -1 0 469900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3951
timestamp 1587416550
transform 0 1 676807 -1 0 470100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3952
timestamp 1587416550
transform 0 1 676807 -1 0 470300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3953
timestamp 1587416550
transform 0 1 676807 -1 0 470500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3954
timestamp 1587416550
transform 0 1 676807 -1 0 470700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3955
timestamp 1587416550
transform 0 1 676807 -1 0 470900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3956
timestamp 1587416550
transform 0 1 676807 -1 0 471100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3957
timestamp 1587416550
transform 0 1 676807 -1 0 471300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3958
timestamp 1587416550
transform 0 1 676807 -1 0 471500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3959
timestamp 1587416550
transform 0 1 676807 -1 0 471700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3960
timestamp 1587416550
transform 0 1 676807 -1 0 471900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3961
timestamp 1587416550
transform 0 1 676807 -1 0 472100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3962
timestamp 1587416550
transform 0 1 676807 -1 0 472300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3963
timestamp 1587416550
transform 0 1 676807 -1 0 472500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3964
timestamp 1587416550
transform 0 1 676807 -1 0 472700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3965
timestamp 1587416550
transform 0 1 676807 -1 0 472900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3966
timestamp 1587416550
transform 0 1 676807 -1 0 473100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3967
timestamp 1587416550
transform 0 1 676807 -1 0 473300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3968
timestamp 1587416550
transform 0 1 676807 -1 0 473500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3969
timestamp 1587416550
transform 0 1 676807 -1 0 473700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3970
timestamp 1587416550
transform 0 1 676807 -1 0 473900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3971
timestamp 1587416550
transform 0 1 676807 -1 0 474100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3972
timestamp 1587416550
transform 0 1 676807 -1 0 474300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3973
timestamp 1587416550
transform 0 1 676807 -1 0 474500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3974
timestamp 1587416550
transform 0 1 676807 -1 0 474700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3975
timestamp 1587416550
transform 0 1 676807 -1 0 474900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3976
timestamp 1587416550
transform 0 1 676807 -1 0 475100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3977
timestamp 1587416550
transform 0 1 676807 -1 0 475300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3978
timestamp 1587416550
transform 0 1 676807 -1 0 475500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3979
timestamp 1587416550
transform 0 1 676807 -1 0 475700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3980
timestamp 1587416550
transform 0 1 676807 -1 0 475900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3981
timestamp 1587416550
transform 0 1 676807 -1 0 476100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3982
timestamp 1587416550
transform 0 1 676807 -1 0 476300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3983
timestamp 1587416550
transform 0 1 676807 -1 0 476500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3984
timestamp 1587416550
transform 0 1 676807 -1 0 476700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3985
timestamp 1587416550
transform 0 1 676807 -1 0 476900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3986
timestamp 1587416550
transform 0 1 676807 -1 0 477100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3987
timestamp 1587416550
transform 0 1 676807 -1 0 477300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3988
timestamp 1587416550
transform 0 1 676807 -1 0 477500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3989
timestamp 1587416550
transform 0 1 676807 -1 0 477700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3990
timestamp 1587416550
transform 0 1 676807 -1 0 477900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3991
timestamp 1587416550
transform 0 1 676807 -1 0 478100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3992
timestamp 1587416550
transform 0 1 676807 -1 0 478300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3993
timestamp 1587416550
transform 0 1 676807 -1 0 478500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3994
timestamp 1587416550
transform 0 1 676807 -1 0 478700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3995
timestamp 1587416550
transform 0 1 676807 -1 0 478900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3996
timestamp 1587416550
transform 0 1 676807 -1 0 479100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3997
timestamp 1587416550
transform 0 1 676807 -1 0 479300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3998
timestamp 1587416550
transform 0 1 676807 -1 0 479500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3999
timestamp 1587416550
transform 0 1 676807 -1 0 479700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4000
timestamp 1587416550
transform 0 1 676807 -1 0 479900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4001
timestamp 1587416550
transform 0 1 676807 -1 0 480100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4002
timestamp 1587416550
transform 0 1 676807 -1 0 480300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4003
timestamp 1587416550
transform 0 1 676807 -1 0 480500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4004
timestamp 1587416550
transform 0 1 676807 -1 0 480700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4006
timestamp 1587416550
transform 0 1 676807 -1 0 481100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4005
timestamp 1587416550
transform 0 1 676807 -1 0 480900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4007
timestamp 1587416550
transform 0 1 676807 -1 0 481300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4008
timestamp 1587416550
transform 0 1 676807 -1 0 481500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4009
timestamp 1587416550
transform 0 1 676807 -1 0 481700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4010
timestamp 1587416550
transform 0 1 676807 -1 0 481900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4012
timestamp 1587416550
transform 0 1 676807 -1 0 482300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4011
timestamp 1587416550
transform 0 1 676807 -1 0 482100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4013
timestamp 1587416550
transform 0 1 676807 -1 0 482500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4014
timestamp 1587416550
transform 0 1 676807 -1 0 482700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4015
timestamp 1587416550
transform 0 1 676807 -1 0 482900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4016
timestamp 1587416550
transform 0 1 676807 -1 0 483100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4017
timestamp 1587416550
transform 0 1 676807 -1 0 483300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4018
timestamp 1587416550
transform 0 1 676807 -1 0 483500
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad  gpio_pad[4]
timestamp 1587416550
transform 0 1 676807 -1 0 499500
box -143 -414 16134 39593
use sky130_ef_io__gpiov2_pad  comp_inn_pad
timestamp 1587416550
transform -1 0 398400 0 -1 259093
box -143 -414 16134 39593
use sky130_ef_io__gpiov2_pad  adc_low_pad
timestamp 1587416550
transform -1 0 431000 0 -1 259093
box -143 -414 16134 39593
use sky130_ef_io__gpiov2_pad  adc_high_pad
timestamp 1587416550
transform -1 0 463400 0 -1 259093
box -143 -414 16134 39593
use sky130_ef_io__gpiov2_pad  adc1_in_pad
timestamp 1587416550
transform -1 0 496000 0 -1 259093
box -143 -414 16134 39593
use sky130_ef_io__gpiov2_pad  adc0_in_pad
timestamp 1587416550
transform -1 0 528600 0 -1 259093
box -143 -414 16134 39593
use sky130_ef_io__gpiov2_pad  xo_pad
timestamp 1587416550
transform -1 0 561200 0 -1 259093
box -143 -414 16134 39593
use sky130_ef_io__gpiov2_pad  xi_pad
timestamp 1587416550
transform -1 0 593800 0 -1 259093
box -143 -414 16134 39593
use sky130_ef_io__gpiov2_pad  gpio_pad[10]
timestamp 1587416550
transform -1 0 626400 0 -1 259093
box -143 -414 16134 39593
use sky130_ef_io__gpiov2_pad  gpio_pad[9]
timestamp 1587416550
transform -1 0 659000 0 -1 259093
box -143 -414 16134 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2806
timestamp 1587416550
transform 0 -1 207593 1 0 502300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2805
timestamp 1587416550
transform 0 -1 207593 1 0 502100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2807
timestamp 1587416550
transform 0 -1 207593 1 0 502500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2808
timestamp 1587416550
transform 0 -1 207593 1 0 502700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2809
timestamp 1587416550
transform 0 -1 207593 1 0 502900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2811
timestamp 1587416550
transform 0 -1 207593 1 0 503300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2810
timestamp 1587416550
transform 0 -1 207593 1 0 503100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2813
timestamp 1587416550
transform 0 -1 207593 1 0 503700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2812
timestamp 1587416550
transform 0 -1 207593 1 0 503500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2815
timestamp 1587416550
transform 0 -1 207593 1 0 504100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2814
timestamp 1587416550
transform 0 -1 207593 1 0 503900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2817
timestamp 1587416550
transform 0 -1 207593 1 0 504500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2816
timestamp 1587416550
transform 0 -1 207593 1 0 504300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2819
timestamp 1587416550
transform 0 -1 207593 1 0 504900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2818
timestamp 1587416550
transform 0 -1 207593 1 0 504700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2820
timestamp 1587416550
transform 0 -1 207593 1 0 505100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2821
timestamp 1587416550
transform 0 -1 207593 1 0 505300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2822
timestamp 1587416550
transform 0 -1 207593 1 0 505500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2824
timestamp 1587416550
transform 0 -1 207593 1 0 505900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2823
timestamp 1587416550
transform 0 -1 207593 1 0 505700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2826
timestamp 1587416550
transform 0 -1 207593 1 0 506300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2825
timestamp 1587416550
transform 0 -1 207593 1 0 506100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2828
timestamp 1587416550
transform 0 -1 207593 1 0 506700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2827
timestamp 1587416550
transform 0 -1 207593 1 0 506500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2830
timestamp 1587416550
transform 0 -1 207593 1 0 507100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2829
timestamp 1587416550
transform 0 -1 207593 1 0 506900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2832
timestamp 1587416550
transform 0 -1 207593 1 0 507500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2831
timestamp 1587416550
transform 0 -1 207593 1 0 507300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2833
timestamp 1587416550
transform 0 -1 207593 1 0 507700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2834
timestamp 1587416550
transform 0 -1 207593 1 0 507900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2835
timestamp 1587416550
transform 0 -1 207593 1 0 508100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2836
timestamp 1587416550
transform 0 -1 207593 1 0 508300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2837
timestamp 1587416550
transform 0 -1 207593 1 0 508500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2839
timestamp 1587416550
transform 0 -1 207593 1 0 508900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2838
timestamp 1587416550
transform 0 -1 207593 1 0 508700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2841
timestamp 1587416550
transform 0 -1 207593 1 0 509300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2840
timestamp 1587416550
transform 0 -1 207593 1 0 509100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2843
timestamp 1587416550
transform 0 -1 207593 1 0 509700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2842
timestamp 1587416550
transform 0 -1 207593 1 0 509500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2845
timestamp 1587416550
transform 0 -1 207593 1 0 510100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2844
timestamp 1587416550
transform 0 -1 207593 1 0 509900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2846
timestamp 1587416550
transform 0 -1 207593 1 0 510300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2847
timestamp 1587416550
transform 0 -1 207593 1 0 510500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2850
timestamp 1587416550
transform 0 -1 207593 1 0 511100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2848
timestamp 1587416550
transform 0 -1 207593 1 0 510700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2849
timestamp 1587416550
transform 0 -1 207593 1 0 510900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2853
timestamp 1587416550
transform 0 -1 207593 1 0 511700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2851
timestamp 1587416550
transform 0 -1 207593 1 0 511300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2852
timestamp 1587416550
transform 0 -1 207593 1 0 511500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2854
timestamp 1587416550
transform 0 -1 207593 1 0 511900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2855
timestamp 1587416550
transform 0 -1 207593 1 0 512100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2856
timestamp 1587416550
transform 0 -1 207593 1 0 512300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2857
timestamp 1587416550
transform 0 -1 207593 1 0 512500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2858
timestamp 1587416550
transform 0 -1 207593 1 0 512700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2859
timestamp 1587416550
transform 0 -1 207593 1 0 512900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2860
timestamp 1587416550
transform 0 -1 207593 1 0 513100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2861
timestamp 1587416550
transform 0 -1 207593 1 0 513300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2863
timestamp 1587416550
transform 0 -1 207593 1 0 529500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2864
timestamp 1587416550
transform 0 -1 207593 1 0 529700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2866
timestamp 1587416550
transform 0 -1 207593 1 0 530100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2865
timestamp 1587416550
transform 0 -1 207593 1 0 529900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2867
timestamp 1587416550
transform 0 -1 207593 1 0 530300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2869
timestamp 1587416550
transform 0 -1 207593 1 0 530700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2868
timestamp 1587416550
transform 0 -1 207593 1 0 530500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2870
timestamp 1587416550
transform 0 -1 207593 1 0 530900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2871
timestamp 1587416550
transform 0 -1 207593 1 0 531100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2872
timestamp 1587416550
transform 0 -1 207593 1 0 531300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2874
timestamp 1587416550
transform 0 -1 207593 1 0 531700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2873
timestamp 1587416550
transform 0 -1 207593 1 0 531500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2875
timestamp 1587416550
transform 0 -1 207593 1 0 531900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2877
timestamp 1587416550
transform 0 -1 207593 1 0 532300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2876
timestamp 1587416550
transform 0 -1 207593 1 0 532100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2878
timestamp 1587416550
transform 0 -1 207593 1 0 532500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2879
timestamp 1587416550
transform 0 -1 207593 1 0 532700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2880
timestamp 1587416550
transform 0 -1 207593 1 0 532900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2882
timestamp 1587416550
transform 0 -1 207593 1 0 533300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2881
timestamp 1587416550
transform 0 -1 207593 1 0 533100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2883
timestamp 1587416550
transform 0 -1 207593 1 0 533500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2885
timestamp 1587416550
transform 0 -1 207593 1 0 533900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2884
timestamp 1587416550
transform 0 -1 207593 1 0 533700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2886
timestamp 1587416550
transform 0 -1 207593 1 0 534100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2887
timestamp 1587416550
transform 0 -1 207593 1 0 534300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2888
timestamp 1587416550
transform 0 -1 207593 1 0 534500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2890
timestamp 1587416550
transform 0 -1 207593 1 0 534900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2889
timestamp 1587416550
transform 0 -1 207593 1 0 534700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2891
timestamp 1587416550
transform 0 -1 207593 1 0 535100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2892
timestamp 1587416550
transform 0 -1 207593 1 0 535300
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad  flash_clk_pad
timestamp 1587416550
transform 0 -1 207593 1 0 513500
box -143 -414 16134 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4020
timestamp 1587416550
transform 0 1 676807 -1 0 499700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4022
timestamp 1587416550
transform 0 1 676807 -1 0 500100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4021
timestamp 1587416550
transform 0 1 676807 -1 0 499900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4023
timestamp 1587416550
transform 0 1 676807 -1 0 500300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4024
timestamp 1587416550
transform 0 1 676807 -1 0 500500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4025
timestamp 1587416550
transform 0 1 676807 -1 0 500700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4026
timestamp 1587416550
transform 0 1 676807 -1 0 500900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4027
timestamp 1587416550
transform 0 1 676807 -1 0 501100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4029
timestamp 1587416550
transform 0 1 676807 -1 0 501500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4028
timestamp 1587416550
transform 0 1 676807 -1 0 501300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4030
timestamp 1587416550
transform 0 1 676807 -1 0 501700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4032
timestamp 1587416550
transform 0 1 676807 -1 0 502100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4031
timestamp 1587416550
transform 0 1 676807 -1 0 501900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4033
timestamp 1587416550
transform 0 1 676807 -1 0 502300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4034
timestamp 1587416550
transform 0 1 676807 -1 0 502500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4035
timestamp 1587416550
transform 0 1 676807 -1 0 502700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4036
timestamp 1587416550
transform 0 1 676807 -1 0 502900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4037
timestamp 1587416550
transform 0 1 676807 -1 0 503100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4039
timestamp 1587416550
transform 0 1 676807 -1 0 503500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4038
timestamp 1587416550
transform 0 1 676807 -1 0 503300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4040
timestamp 1587416550
transform 0 1 676807 -1 0 503700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4042
timestamp 1587416550
transform 0 1 676807 -1 0 504100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4041
timestamp 1587416550
transform 0 1 676807 -1 0 503900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4043
timestamp 1587416550
transform 0 1 676807 -1 0 504300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4044
timestamp 1587416550
transform 0 1 676807 -1 0 504500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4045
timestamp 1587416550
transform 0 1 676807 -1 0 504700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4046
timestamp 1587416550
transform 0 1 676807 -1 0 504900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4047
timestamp 1587416550
transform 0 1 676807 -1 0 505100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4049
timestamp 1587416550
transform 0 1 676807 -1 0 505500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4048
timestamp 1587416550
transform 0 1 676807 -1 0 505300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4050
timestamp 1587416550
transform 0 1 676807 -1 0 505700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4051
timestamp 1587416550
transform 0 1 676807 -1 0 505900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4052
timestamp 1587416550
transform 0 1 676807 -1 0 506100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4053
timestamp 1587416550
transform 0 1 676807 -1 0 506300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4054
timestamp 1587416550
transform 0 1 676807 -1 0 506500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4055
timestamp 1587416550
transform 0 1 676807 -1 0 506700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4056
timestamp 1587416550
transform 0 1 676807 -1 0 506900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4057
timestamp 1587416550
transform 0 1 676807 -1 0 507100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4059
timestamp 1587416550
transform 0 1 676807 -1 0 507500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4058
timestamp 1587416550
transform 0 1 676807 -1 0 507300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4060
timestamp 1587416550
transform 0 1 676807 -1 0 507700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4061
timestamp 1587416550
transform 0 1 676807 -1 0 507900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4062
timestamp 1587416550
transform 0 1 676807 -1 0 508100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4063
timestamp 1587416550
transform 0 1 676807 -1 0 508300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4064
timestamp 1587416550
transform 0 1 676807 -1 0 508500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4065
timestamp 1587416550
transform 0 1 676807 -1 0 508700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4066
timestamp 1587416550
transform 0 1 676807 -1 0 508900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4067
timestamp 1587416550
transform 0 1 676807 -1 0 509100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4069
timestamp 1587416550
transform 0 1 676807 -1 0 509500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4068
timestamp 1587416550
transform 0 1 676807 -1 0 509300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4070
timestamp 1587416550
transform 0 1 676807 -1 0 509700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4071
timestamp 1587416550
transform 0 1 676807 -1 0 509900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4072
timestamp 1587416550
transform 0 1 676807 -1 0 510100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4073
timestamp 1587416550
transform 0 1 676807 -1 0 510300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4074
timestamp 1587416550
transform 0 1 676807 -1 0 510500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4075
timestamp 1587416550
transform 0 1 676807 -1 0 510700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4076
timestamp 1587416550
transform 0 1 676807 -1 0 510900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4077
timestamp 1587416550
transform 0 1 676807 -1 0 511100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4078
timestamp 1587416550
transform 0 1 676807 -1 0 511300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4079
timestamp 1587416550
transform 0 1 676807 -1 0 511500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4080
timestamp 1587416550
transform 0 1 676807 -1 0 511700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4081
timestamp 1587416550
transform 0 1 676807 -1 0 511900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4082
timestamp 1587416550
transform 0 1 676807 -1 0 512100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4083
timestamp 1587416550
transform 0 1 676807 -1 0 512300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4084
timestamp 1587416550
transform 0 1 676807 -1 0 512500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4085
timestamp 1587416550
transform 0 1 676807 -1 0 512700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4086
timestamp 1587416550
transform 0 1 676807 -1 0 512900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4087
timestamp 1587416550
transform 0 1 676807 -1 0 513100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4088
timestamp 1587416550
transform 0 1 676807 -1 0 513300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4089
timestamp 1587416550
transform 0 1 676807 -1 0 513500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4090
timestamp 1587416550
transform 0 1 676807 -1 0 513700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4091
timestamp 1587416550
transform 0 1 676807 -1 0 513900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4092
timestamp 1587416550
transform 0 1 676807 -1 0 514100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4093
timestamp 1587416550
transform 0 1 676807 -1 0 514300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4094
timestamp 1587416550
transform 0 1 676807 -1 0 514500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4095
timestamp 1587416550
transform 0 1 676807 -1 0 514700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4096
timestamp 1587416550
transform 0 1 676807 -1 0 514900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4097
timestamp 1587416550
transform 0 1 676807 -1 0 515100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4098
timestamp 1587416550
transform 0 1 676807 -1 0 515300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4099
timestamp 1587416550
transform 0 1 676807 -1 0 515500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4100
timestamp 1587416550
transform 0 1 676807 -1 0 515700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4101
timestamp 1587416550
transform 0 1 676807 -1 0 515900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4102
timestamp 1587416550
transform 0 1 676807 -1 0 516100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4103
timestamp 1587416550
transform 0 1 676807 -1 0 516300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4104
timestamp 1587416550
transform 0 1 676807 -1 0 516500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4105
timestamp 1587416550
transform 0 1 676807 -1 0 516700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4106
timestamp 1587416550
transform 0 1 676807 -1 0 516900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4107
timestamp 1587416550
transform 0 1 676807 -1 0 517100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4108
timestamp 1587416550
transform 0 1 676807 -1 0 517300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4109
timestamp 1587416550
transform 0 1 676807 -1 0 517500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4110
timestamp 1587416550
transform 0 1 676807 -1 0 517700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4111
timestamp 1587416550
transform 0 1 676807 -1 0 517900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4112
timestamp 1587416550
transform 0 1 676807 -1 0 518100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4113
timestamp 1587416550
transform 0 1 676807 -1 0 518300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4114
timestamp 1587416550
transform 0 1 676807 -1 0 518500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4115
timestamp 1587416550
transform 0 1 676807 -1 0 518700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4116
timestamp 1587416550
transform 0 1 676807 -1 0 518900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4118
timestamp 1587416550
transform 0 1 676807 -1 0 519300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4117
timestamp 1587416550
transform 0 1 676807 -1 0 519100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4119
timestamp 1587416550
transform 0 1 676807 -1 0 519500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4121
timestamp 1587416550
transform 0 1 676807 -1 0 519900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4120
timestamp 1587416550
transform 0 1 676807 -1 0 519700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4122
timestamp 1587416550
transform 0 1 676807 -1 0 520100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4124
timestamp 1587416550
transform 0 1 676807 -1 0 520500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4123
timestamp 1587416550
transform 0 1 676807 -1 0 520300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4125
timestamp 1587416550
transform 0 1 676807 -1 0 520700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4126
timestamp 1587416550
transform 0 1 676807 -1 0 520900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4128
timestamp 1587416550
transform 0 1 676807 -1 0 521300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4127
timestamp 1587416550
transform 0 1 676807 -1 0 521100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4129
timestamp 1587416550
transform 0 1 676807 -1 0 521500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4131
timestamp 1587416550
transform 0 1 676807 -1 0 521900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4130
timestamp 1587416550
transform 0 1 676807 -1 0 521700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4132
timestamp 1587416550
transform 0 1 676807 -1 0 522100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4134
timestamp 1587416550
transform 0 1 676807 -1 0 522500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4133
timestamp 1587416550
transform 0 1 676807 -1 0 522300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4135
timestamp 1587416550
transform 0 1 676807 -1 0 522700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4136
timestamp 1587416550
transform 0 1 676807 -1 0 522900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4138
timestamp 1587416550
transform 0 1 676807 -1 0 523300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4137
timestamp 1587416550
transform 0 1 676807 -1 0 523100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4139
timestamp 1587416550
transform 0 1 676807 -1 0 523500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4141
timestamp 1587416550
transform 0 1 676807 -1 0 523900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4140
timestamp 1587416550
transform 0 1 676807 -1 0 523700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4142
timestamp 1587416550
transform 0 1 676807 -1 0 524100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4143
timestamp 1587416550
transform 0 1 676807 -1 0 524300
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad  gpio_pad[3]
timestamp 1587416550
transform 0 1 676807 -1 0 540300
box -143 -414 16134 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2893
timestamp 1587416550
transform 0 -1 207593 1 0 535500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2894
timestamp 1587416550
transform 0 -1 207593 1 0 535700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2895
timestamp 1587416550
transform 0 -1 207593 1 0 535900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2896
timestamp 1587416550
transform 0 -1 207593 1 0 536100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2897
timestamp 1587416550
transform 0 -1 207593 1 0 536300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2898
timestamp 1587416550
transform 0 -1 207593 1 0 536500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2899
timestamp 1587416550
transform 0 -1 207593 1 0 536700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2900
timestamp 1587416550
transform 0 -1 207593 1 0 536900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2901
timestamp 1587416550
transform 0 -1 207593 1 0 537100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2902
timestamp 1587416550
transform 0 -1 207593 1 0 537300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2903
timestamp 1587416550
transform 0 -1 207593 1 0 537500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2904
timestamp 1587416550
transform 0 -1 207593 1 0 537700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2905
timestamp 1587416550
transform 0 -1 207593 1 0 537900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2906
timestamp 1587416550
transform 0 -1 207593 1 0 538100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2907
timestamp 1587416550
transform 0 -1 207593 1 0 538300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2908
timestamp 1587416550
transform 0 -1 207593 1 0 538500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2909
timestamp 1587416550
transform 0 -1 207593 1 0 538700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2910
timestamp 1587416550
transform 0 -1 207593 1 0 538900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2911
timestamp 1587416550
transform 0 -1 207593 1 0 539100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2912
timestamp 1587416550
transform 0 -1 207593 1 0 539300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2913
timestamp 1587416550
transform 0 -1 207593 1 0 539500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2914
timestamp 1587416550
transform 0 -1 207593 1 0 539700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2915
timestamp 1587416550
transform 0 -1 207593 1 0 539900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2916
timestamp 1587416550
transform 0 -1 207593 1 0 540100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2917
timestamp 1587416550
transform 0 -1 207593 1 0 540300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2918
timestamp 1587416550
transform 0 -1 207593 1 0 540500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2919
timestamp 1587416550
transform 0 -1 207593 1 0 540700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2921
timestamp 1587416550
transform 0 -1 207593 1 0 556900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2922
timestamp 1587416550
transform 0 -1 207593 1 0 557100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2923
timestamp 1587416550
transform 0 -1 207593 1 0 557300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2924
timestamp 1587416550
transform 0 -1 207593 1 0 557500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2925
timestamp 1587416550
transform 0 -1 207593 1 0 557700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2926
timestamp 1587416550
transform 0 -1 207593 1 0 557900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2927
timestamp 1587416550
transform 0 -1 207593 1 0 558100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2928
timestamp 1587416550
transform 0 -1 207593 1 0 558300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2929
timestamp 1587416550
transform 0 -1 207593 1 0 558500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2930
timestamp 1587416550
transform 0 -1 207593 1 0 558700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2931
timestamp 1587416550
transform 0 -1 207593 1 0 558900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2932
timestamp 1587416550
transform 0 -1 207593 1 0 559100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2933
timestamp 1587416550
transform 0 -1 207593 1 0 559300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2934
timestamp 1587416550
transform 0 -1 207593 1 0 559500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2935
timestamp 1587416550
transform 0 -1 207593 1 0 559700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2936
timestamp 1587416550
transform 0 -1 207593 1 0 559900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2937
timestamp 1587416550
transform 0 -1 207593 1 0 560100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2938
timestamp 1587416550
transform 0 -1 207593 1 0 560300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2939
timestamp 1587416550
transform 0 -1 207593 1 0 560500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2940
timestamp 1587416550
transform 0 -1 207593 1 0 560700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2941
timestamp 1587416550
transform 0 -1 207593 1 0 560900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2942
timestamp 1587416550
transform 0 -1 207593 1 0 561100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2943
timestamp 1587416550
transform 0 -1 207593 1 0 561300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2944
timestamp 1587416550
transform 0 -1 207593 1 0 561500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2945
timestamp 1587416550
transform 0 -1 207593 1 0 561700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2946
timestamp 1587416550
transform 0 -1 207593 1 0 561900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2947
timestamp 1587416550
transform 0 -1 207593 1 0 562100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2948
timestamp 1587416550
transform 0 -1 207593 1 0 562300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2949
timestamp 1587416550
transform 0 -1 207593 1 0 562500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2950
timestamp 1587416550
transform 0 -1 207593 1 0 562700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2951
timestamp 1587416550
transform 0 -1 207593 1 0 562900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2952
timestamp 1587416550
transform 0 -1 207593 1 0 563100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2953
timestamp 1587416550
transform 0 -1 207593 1 0 563300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2954
timestamp 1587416550
transform 0 -1 207593 1 0 563500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2955
timestamp 1587416550
transform 0 -1 207593 1 0 563700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2956
timestamp 1587416550
transform 0 -1 207593 1 0 563900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2957
timestamp 1587416550
transform 0 -1 207593 1 0 564100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2958
timestamp 1587416550
transform 0 -1 207593 1 0 564300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2959
timestamp 1587416550
transform 0 -1 207593 1 0 564500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2960
timestamp 1587416550
transform 0 -1 207593 1 0 564700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2961
timestamp 1587416550
transform 0 -1 207593 1 0 564900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2962
timestamp 1587416550
transform 0 -1 207593 1 0 565100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2963
timestamp 1587416550
transform 0 -1 207593 1 0 565300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2964
timestamp 1587416550
transform 0 -1 207593 1 0 565500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2965
timestamp 1587416550
transform 0 -1 207593 1 0 565700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2966
timestamp 1587416550
transform 0 -1 207593 1 0 565900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2967
timestamp 1587416550
transform 0 -1 207593 1 0 566100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2968
timestamp 1587416550
transform 0 -1 207593 1 0 566300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2969
timestamp 1587416550
transform 0 -1 207593 1 0 566500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2970
timestamp 1587416550
transform 0 -1 207593 1 0 566700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2971
timestamp 1587416550
transform 0 -1 207593 1 0 566900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2972
timestamp 1587416550
transform 0 -1 207593 1 0 567100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2973
timestamp 1587416550
transform 0 -1 207593 1 0 567300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2974
timestamp 1587416550
transform 0 -1 207593 1 0 567500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2975
timestamp 1587416550
transform 0 -1 207593 1 0 567700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2976
timestamp 1587416550
transform 0 -1 207593 1 0 567900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2977
timestamp 1587416550
transform 0 -1 207593 1 0 568100
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad  flash_io0_pad
timestamp 1587416550
transform 0 -1 207593 1 0 540900
box -143 -414 16134 39593
use sky130_ef_io__gpiov2_pad  flash_io1_pad
timestamp 1587416550
transform 0 -1 207593 1 0 568300
box -143 -414 16134 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4145
timestamp 1587416550
transform 0 1 676807 -1 0 540500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4147
timestamp 1587416550
transform 0 1 676807 -1 0 540900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4146
timestamp 1587416550
transform 0 1 676807 -1 0 540700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4148
timestamp 1587416550
transform 0 1 676807 -1 0 541100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4149
timestamp 1587416550
transform 0 1 676807 -1 0 541300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4150
timestamp 1587416550
transform 0 1 676807 -1 0 541500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4151
timestamp 1587416550
transform 0 1 676807 -1 0 541700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4152
timestamp 1587416550
transform 0 1 676807 -1 0 541900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4154
timestamp 1587416550
transform 0 1 676807 -1 0 542300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4153
timestamp 1587416550
transform 0 1 676807 -1 0 542100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4155
timestamp 1587416550
transform 0 1 676807 -1 0 542500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4157
timestamp 1587416550
transform 0 1 676807 -1 0 542900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4156
timestamp 1587416550
transform 0 1 676807 -1 0 542700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4158
timestamp 1587416550
transform 0 1 676807 -1 0 543100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4159
timestamp 1587416550
transform 0 1 676807 -1 0 543300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4160
timestamp 1587416550
transform 0 1 676807 -1 0 543500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4161
timestamp 1587416550
transform 0 1 676807 -1 0 543700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4162
timestamp 1587416550
transform 0 1 676807 -1 0 543900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4164
timestamp 1587416550
transform 0 1 676807 -1 0 544300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4163
timestamp 1587416550
transform 0 1 676807 -1 0 544100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4165
timestamp 1587416550
transform 0 1 676807 -1 0 544500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4167
timestamp 1587416550
transform 0 1 676807 -1 0 544900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4166
timestamp 1587416550
transform 0 1 676807 -1 0 544700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4168
timestamp 1587416550
transform 0 1 676807 -1 0 545100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4169
timestamp 1587416550
transform 0 1 676807 -1 0 545300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4170
timestamp 1587416550
transform 0 1 676807 -1 0 545500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4171
timestamp 1587416550
transform 0 1 676807 -1 0 545700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4172
timestamp 1587416550
transform 0 1 676807 -1 0 545900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4174
timestamp 1587416550
transform 0 1 676807 -1 0 546300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4173
timestamp 1587416550
transform 0 1 676807 -1 0 546100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4175
timestamp 1587416550
transform 0 1 676807 -1 0 546500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4177
timestamp 1587416550
transform 0 1 676807 -1 0 546900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4176
timestamp 1587416550
transform 0 1 676807 -1 0 546700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4178
timestamp 1587416550
transform 0 1 676807 -1 0 547100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4179
timestamp 1587416550
transform 0 1 676807 -1 0 547300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4180
timestamp 1587416550
transform 0 1 676807 -1 0 547500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4181
timestamp 1587416550
transform 0 1 676807 -1 0 547700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4182
timestamp 1587416550
transform 0 1 676807 -1 0 547900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4184
timestamp 1587416550
transform 0 1 676807 -1 0 548300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4183
timestamp 1587416550
transform 0 1 676807 -1 0 548100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4185
timestamp 1587416550
transform 0 1 676807 -1 0 548500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4186
timestamp 1587416550
transform 0 1 676807 -1 0 548700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4187
timestamp 1587416550
transform 0 1 676807 -1 0 548900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4188
timestamp 1587416550
transform 0 1 676807 -1 0 549100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4189
timestamp 1587416550
transform 0 1 676807 -1 0 549300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4190
timestamp 1587416550
transform 0 1 676807 -1 0 549500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4191
timestamp 1587416550
transform 0 1 676807 -1 0 549700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4192
timestamp 1587416550
transform 0 1 676807 -1 0 549900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4194
timestamp 1587416550
transform 0 1 676807 -1 0 550300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4193
timestamp 1587416550
transform 0 1 676807 -1 0 550100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4195
timestamp 1587416550
transform 0 1 676807 -1 0 550500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4196
timestamp 1587416550
transform 0 1 676807 -1 0 550700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4197
timestamp 1587416550
transform 0 1 676807 -1 0 550900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4198
timestamp 1587416550
transform 0 1 676807 -1 0 551100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4199
timestamp 1587416550
transform 0 1 676807 -1 0 551300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4200
timestamp 1587416550
transform 0 1 676807 -1 0 551500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4201
timestamp 1587416550
transform 0 1 676807 -1 0 551700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4202
timestamp 1587416550
transform 0 1 676807 -1 0 551900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4203
timestamp 1587416550
transform 0 1 676807 -1 0 552100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4204
timestamp 1587416550
transform 0 1 676807 -1 0 552300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4205
timestamp 1587416550
transform 0 1 676807 -1 0 552500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4206
timestamp 1587416550
transform 0 1 676807 -1 0 552700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4207
timestamp 1587416550
transform 0 1 676807 -1 0 552900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4208
timestamp 1587416550
transform 0 1 676807 -1 0 553100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4209
timestamp 1587416550
transform 0 1 676807 -1 0 553300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4210
timestamp 1587416550
transform 0 1 676807 -1 0 553500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4211
timestamp 1587416550
transform 0 1 676807 -1 0 553700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4212
timestamp 1587416550
transform 0 1 676807 -1 0 553900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4213
timestamp 1587416550
transform 0 1 676807 -1 0 554100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4214
timestamp 1587416550
transform 0 1 676807 -1 0 554300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4215
timestamp 1587416550
transform 0 1 676807 -1 0 554500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4216
timestamp 1587416550
transform 0 1 676807 -1 0 554700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4217
timestamp 1587416550
transform 0 1 676807 -1 0 554900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4218
timestamp 1587416550
transform 0 1 676807 -1 0 555100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4219
timestamp 1587416550
transform 0 1 676807 -1 0 555300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4220
timestamp 1587416550
transform 0 1 676807 -1 0 555500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4221
timestamp 1587416550
transform 0 1 676807 -1 0 555700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4222
timestamp 1587416550
transform 0 1 676807 -1 0 555900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4223
timestamp 1587416550
transform 0 1 676807 -1 0 556100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4224
timestamp 1587416550
transform 0 1 676807 -1 0 556300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4225
timestamp 1587416550
transform 0 1 676807 -1 0 556500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4226
timestamp 1587416550
transform 0 1 676807 -1 0 556700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4227
timestamp 1587416550
transform 0 1 676807 -1 0 556900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4228
timestamp 1587416550
transform 0 1 676807 -1 0 557100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4229
timestamp 1587416550
transform 0 1 676807 -1 0 557300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4230
timestamp 1587416550
transform 0 1 676807 -1 0 557500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4231
timestamp 1587416550
transform 0 1 676807 -1 0 557700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4232
timestamp 1587416550
transform 0 1 676807 -1 0 557900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4233
timestamp 1587416550
transform 0 1 676807 -1 0 558100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4234
timestamp 1587416550
transform 0 1 676807 -1 0 558300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4235
timestamp 1587416550
transform 0 1 676807 -1 0 558500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4236
timestamp 1587416550
transform 0 1 676807 -1 0 558700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4237
timestamp 1587416550
transform 0 1 676807 -1 0 558900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4238
timestamp 1587416550
transform 0 1 676807 -1 0 559100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4239
timestamp 1587416550
transform 0 1 676807 -1 0 559300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4240
timestamp 1587416550
transform 0 1 676807 -1 0 559500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4241
timestamp 1587416550
transform 0 1 676807 -1 0 559700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4243
timestamp 1587416550
transform 0 1 676807 -1 0 560100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4242
timestamp 1587416550
transform 0 1 676807 -1 0 559900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4244
timestamp 1587416550
transform 0 1 676807 -1 0 560300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4246
timestamp 1587416550
transform 0 1 676807 -1 0 560700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4245
timestamp 1587416550
transform 0 1 676807 -1 0 560500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4247
timestamp 1587416550
transform 0 1 676807 -1 0 560900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4248
timestamp 1587416550
transform 0 1 676807 -1 0 561100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4250
timestamp 1587416550
transform 0 1 676807 -1 0 561500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4249
timestamp 1587416550
transform 0 1 676807 -1 0 561300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4251
timestamp 1587416550
transform 0 1 676807 -1 0 561700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4252
timestamp 1587416550
transform 0 1 676807 -1 0 561900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4254
timestamp 1587416550
transform 0 1 676807 -1 0 562300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4253
timestamp 1587416550
transform 0 1 676807 -1 0 562100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4255
timestamp 1587416550
transform 0 1 676807 -1 0 562500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4257
timestamp 1587416550
transform 0 1 676807 -1 0 562900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4256
timestamp 1587416550
transform 0 1 676807 -1 0 562700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4258
timestamp 1587416550
transform 0 1 676807 -1 0 563100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4259
timestamp 1587416550
transform 0 1 676807 -1 0 563300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4261
timestamp 1587416550
transform 0 1 676807 -1 0 563700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4260
timestamp 1587416550
transform 0 1 676807 -1 0 563500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4262
timestamp 1587416550
transform 0 1 676807 -1 0 563900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4264
timestamp 1587416550
transform 0 1 676807 -1 0 564300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4263
timestamp 1587416550
transform 0 1 676807 -1 0 564100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4265
timestamp 1587416550
transform 0 1 676807 -1 0 564500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4266
timestamp 1587416550
transform 0 1 676807 -1 0 564700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4268
timestamp 1587416550
transform 0 1 676807 -1 0 565100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4267
timestamp 1587416550
transform 0 1 676807 -1 0 564900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4269
timestamp 1587416550
transform 0 1 676807 -1 0 565300
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad  gpio_pad[2]
timestamp 1587416550
transform 0 1 676807 -1 0 581300
box -143 -414 16134 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2980
timestamp 1587416550
transform 0 -1 207593 1 0 584500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2979
timestamp 1587416550
transform 0 -1 207593 1 0 584300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2982
timestamp 1587416550
transform 0 -1 207593 1 0 584900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2981
timestamp 1587416550
transform 0 -1 207593 1 0 584700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2984
timestamp 1587416550
transform 0 -1 207593 1 0 585300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2983
timestamp 1587416550
transform 0 -1 207593 1 0 585100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2986
timestamp 1587416550
transform 0 -1 207593 1 0 585700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2985
timestamp 1587416550
transform 0 -1 207593 1 0 585500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2988
timestamp 1587416550
transform 0 -1 207593 1 0 586100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2987
timestamp 1587416550
transform 0 -1 207593 1 0 585900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2990
timestamp 1587416550
transform 0 -1 207593 1 0 586500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2989
timestamp 1587416550
transform 0 -1 207593 1 0 586300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2992
timestamp 1587416550
transform 0 -1 207593 1 0 586900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2991
timestamp 1587416550
transform 0 -1 207593 1 0 586700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2994
timestamp 1587416550
transform 0 -1 207593 1 0 587300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2993
timestamp 1587416550
transform 0 -1 207593 1 0 587100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2996
timestamp 1587416550
transform 0 -1 207593 1 0 587700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2995
timestamp 1587416550
transform 0 -1 207593 1 0 587500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2998
timestamp 1587416550
transform 0 -1 207593 1 0 588100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2997
timestamp 1587416550
transform 0 -1 207593 1 0 587900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3000
timestamp 1587416550
transform 0 -1 207593 1 0 588500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_2999
timestamp 1587416550
transform 0 -1 207593 1 0 588300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3002
timestamp 1587416550
transform 0 -1 207593 1 0 588900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3001
timestamp 1587416550
transform 0 -1 207593 1 0 588700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3004
timestamp 1587416550
transform 0 -1 207593 1 0 589300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3003
timestamp 1587416550
transform 0 -1 207593 1 0 589100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3006
timestamp 1587416550
transform 0 -1 207593 1 0 589700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3005
timestamp 1587416550
transform 0 -1 207593 1 0 589500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3008
timestamp 1587416550
transform 0 -1 207593 1 0 590100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3007
timestamp 1587416550
transform 0 -1 207593 1 0 589900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3010
timestamp 1587416550
transform 0 -1 207593 1 0 590500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3009
timestamp 1587416550
transform 0 -1 207593 1 0 590300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3012
timestamp 1587416550
transform 0 -1 207593 1 0 590900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3011
timestamp 1587416550
transform 0 -1 207593 1 0 590700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3014
timestamp 1587416550
transform 0 -1 207593 1 0 591300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3013
timestamp 1587416550
transform 0 -1 207593 1 0 591100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3016
timestamp 1587416550
transform 0 -1 207593 1 0 591700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3015
timestamp 1587416550
transform 0 -1 207593 1 0 591500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3018
timestamp 1587416550
transform 0 -1 207593 1 0 592100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3017
timestamp 1587416550
transform 0 -1 207593 1 0 591900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3019
timestamp 1587416550
transform 0 -1 207593 1 0 592300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3020
timestamp 1587416550
transform 0 -1 207593 1 0 592500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3023
timestamp 1587416550
transform 0 -1 207593 1 0 593100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3021
timestamp 1587416550
transform 0 -1 207593 1 0 592700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3022
timestamp 1587416550
transform 0 -1 207593 1 0 592900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3024
timestamp 1587416550
transform 0 -1 207593 1 0 593300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3025
timestamp 1587416550
transform 0 -1 207593 1 0 593500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3026
timestamp 1587416550
transform 0 -1 207593 1 0 593700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3027
timestamp 1587416550
transform 0 -1 207593 1 0 593900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3030
timestamp 1587416550
transform 0 -1 207593 1 0 594500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3028
timestamp 1587416550
transform 0 -1 207593 1 0 594100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3029
timestamp 1587416550
transform 0 -1 207593 1 0 594300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3031
timestamp 1587416550
transform 0 -1 207593 1 0 594700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3032
timestamp 1587416550
transform 0 -1 207593 1 0 594900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3033
timestamp 1587416550
transform 0 -1 207593 1 0 595100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3034
timestamp 1587416550
transform 0 -1 207593 1 0 595300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3035
timestamp 1587416550
transform 0 -1 207593 1 0 595500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3037
timestamp 1587416550
transform 0 -1 207593 1 0 611700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3039
timestamp 1587416550
transform 0 -1 207593 1 0 612100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3038
timestamp 1587416550
transform 0 -1 207593 1 0 611900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3040
timestamp 1587416550
transform 0 -1 207593 1 0 612300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3042
timestamp 1587416550
transform 0 -1 207593 1 0 612700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3041
timestamp 1587416550
transform 0 -1 207593 1 0 612500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3043
timestamp 1587416550
transform 0 -1 207593 1 0 612900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3045
timestamp 1587416550
transform 0 -1 207593 1 0 613300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3044
timestamp 1587416550
transform 0 -1 207593 1 0 613100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3046
timestamp 1587416550
transform 0 -1 207593 1 0 613500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3048
timestamp 1587416550
transform 0 -1 207593 1 0 613900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3047
timestamp 1587416550
transform 0 -1 207593 1 0 613700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3049
timestamp 1587416550
transform 0 -1 207593 1 0 614100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3051
timestamp 1587416550
transform 0 -1 207593 1 0 614500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3050
timestamp 1587416550
transform 0 -1 207593 1 0 614300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3052
timestamp 1587416550
transform 0 -1 207593 1 0 614700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3054
timestamp 1587416550
transform 0 -1 207593 1 0 615100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3053
timestamp 1587416550
transform 0 -1 207593 1 0 614900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3055
timestamp 1587416550
transform 0 -1 207593 1 0 615300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3057
timestamp 1587416550
transform 0 -1 207593 1 0 615700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3056
timestamp 1587416550
transform 0 -1 207593 1 0 615500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3058
timestamp 1587416550
transform 0 -1 207593 1 0 615900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3060
timestamp 1587416550
transform 0 -1 207593 1 0 616300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3059
timestamp 1587416550
transform 0 -1 207593 1 0 616100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3061
timestamp 1587416550
transform 0 -1 207593 1 0 616500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3063
timestamp 1587416550
transform 0 -1 207593 1 0 616900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3062
timestamp 1587416550
transform 0 -1 207593 1 0 616700
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad  flash_io2_pad
timestamp 1587416550
transform 0 -1 207593 1 0 595700
box -143 -414 16134 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4271
timestamp 1587416550
transform 0 1 676807 -1 0 581500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4272
timestamp 1587416550
transform 0 1 676807 -1 0 581700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4274
timestamp 1587416550
transform 0 1 676807 -1 0 582100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4273
timestamp 1587416550
transform 0 1 676807 -1 0 581900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4275
timestamp 1587416550
transform 0 1 676807 -1 0 582300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4276
timestamp 1587416550
transform 0 1 676807 -1 0 582500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4277
timestamp 1587416550
transform 0 1 676807 -1 0 582700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4278
timestamp 1587416550
transform 0 1 676807 -1 0 582900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4279
timestamp 1587416550
transform 0 1 676807 -1 0 583100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4280
timestamp 1587416550
transform 0 1 676807 -1 0 583300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4281
timestamp 1587416550
transform 0 1 676807 -1 0 583500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4282
timestamp 1587416550
transform 0 1 676807 -1 0 583700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4284
timestamp 1587416550
transform 0 1 676807 -1 0 584100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4283
timestamp 1587416550
transform 0 1 676807 -1 0 583900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4285
timestamp 1587416550
transform 0 1 676807 -1 0 584300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4287
timestamp 1587416550
transform 0 1 676807 -1 0 584700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4286
timestamp 1587416550
transform 0 1 676807 -1 0 584500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4288
timestamp 1587416550
transform 0 1 676807 -1 0 584900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4289
timestamp 1587416550
transform 0 1 676807 -1 0 585100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4290
timestamp 1587416550
transform 0 1 676807 -1 0 585300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4291
timestamp 1587416550
transform 0 1 676807 -1 0 585500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4292
timestamp 1587416550
transform 0 1 676807 -1 0 585700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4293
timestamp 1587416550
transform 0 1 676807 -1 0 585900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4294
timestamp 1587416550
transform 0 1 676807 -1 0 586100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4295
timestamp 1587416550
transform 0 1 676807 -1 0 586300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4296
timestamp 1587416550
transform 0 1 676807 -1 0 586500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4297
timestamp 1587416550
transform 0 1 676807 -1 0 586700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4298
timestamp 1587416550
transform 0 1 676807 -1 0 586900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4299
timestamp 1587416550
transform 0 1 676807 -1 0 587100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4300
timestamp 1587416550
transform 0 1 676807 -1 0 587300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4301
timestamp 1587416550
transform 0 1 676807 -1 0 587500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4303
timestamp 1587416550
transform 0 1 676807 -1 0 587900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4302
timestamp 1587416550
transform 0 1 676807 -1 0 587700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4304
timestamp 1587416550
transform 0 1 676807 -1 0 588100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4305
timestamp 1587416550
transform 0 1 676807 -1 0 588300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4306
timestamp 1587416550
transform 0 1 676807 -1 0 588500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4307
timestamp 1587416550
transform 0 1 676807 -1 0 588700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4308
timestamp 1587416550
transform 0 1 676807 -1 0 588900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4309
timestamp 1587416550
transform 0 1 676807 -1 0 589100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4310
timestamp 1587416550
transform 0 1 676807 -1 0 589300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4311
timestamp 1587416550
transform 0 1 676807 -1 0 589500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4312
timestamp 1587416550
transform 0 1 676807 -1 0 589700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4313
timestamp 1587416550
transform 0 1 676807 -1 0 589900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4314
timestamp 1587416550
transform 0 1 676807 -1 0 590100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4315
timestamp 1587416550
transform 0 1 676807 -1 0 590300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4316
timestamp 1587416550
transform 0 1 676807 -1 0 590500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4317
timestamp 1587416550
transform 0 1 676807 -1 0 590700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4318
timestamp 1587416550
transform 0 1 676807 -1 0 590900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4319
timestamp 1587416550
transform 0 1 676807 -1 0 591100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4320
timestamp 1587416550
transform 0 1 676807 -1 0 591300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4321
timestamp 1587416550
transform 0 1 676807 -1 0 591500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4322
timestamp 1587416550
transform 0 1 676807 -1 0 591700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4323
timestamp 1587416550
transform 0 1 676807 -1 0 591900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4324
timestamp 1587416550
transform 0 1 676807 -1 0 592100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4325
timestamp 1587416550
transform 0 1 676807 -1 0 592300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4326
timestamp 1587416550
transform 0 1 676807 -1 0 592500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4327
timestamp 1587416550
transform 0 1 676807 -1 0 592700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4328
timestamp 1587416550
transform 0 1 676807 -1 0 592900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4329
timestamp 1587416550
transform 0 1 676807 -1 0 593100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4330
timestamp 1587416550
transform 0 1 676807 -1 0 593300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4331
timestamp 1587416550
transform 0 1 676807 -1 0 593500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4332
timestamp 1587416550
transform 0 1 676807 -1 0 593700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4333
timestamp 1587416550
transform 0 1 676807 -1 0 593900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4334
timestamp 1587416550
transform 0 1 676807 -1 0 594100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4335
timestamp 1587416550
transform 0 1 676807 -1 0 594300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4336
timestamp 1587416550
transform 0 1 676807 -1 0 594500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4337
timestamp 1587416550
transform 0 1 676807 -1 0 594700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4338
timestamp 1587416550
transform 0 1 676807 -1 0 594900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4339
timestamp 1587416550
transform 0 1 676807 -1 0 595100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4340
timestamp 1587416550
transform 0 1 676807 -1 0 595300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4341
timestamp 1587416550
transform 0 1 676807 -1 0 595500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4342
timestamp 1587416550
transform 0 1 676807 -1 0 595700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4343
timestamp 1587416550
transform 0 1 676807 -1 0 595900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4344
timestamp 1587416550
transform 0 1 676807 -1 0 596100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4345
timestamp 1587416550
transform 0 1 676807 -1 0 596300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4346
timestamp 1587416550
transform 0 1 676807 -1 0 596500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4347
timestamp 1587416550
transform 0 1 676807 -1 0 596700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4348
timestamp 1587416550
transform 0 1 676807 -1 0 596900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4349
timestamp 1587416550
transform 0 1 676807 -1 0 597100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4350
timestamp 1587416550
transform 0 1 676807 -1 0 597300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4351
timestamp 1587416550
transform 0 1 676807 -1 0 597500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4352
timestamp 1587416550
transform 0 1 676807 -1 0 597700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4353
timestamp 1587416550
transform 0 1 676807 -1 0 597900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4354
timestamp 1587416550
transform 0 1 676807 -1 0 598100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4355
timestamp 1587416550
transform 0 1 676807 -1 0 598300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4356
timestamp 1587416550
transform 0 1 676807 -1 0 598500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4357
timestamp 1587416550
transform 0 1 676807 -1 0 598700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4358
timestamp 1587416550
transform 0 1 676807 -1 0 598900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4359
timestamp 1587416550
transform 0 1 676807 -1 0 599100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4360
timestamp 1587416550
transform 0 1 676807 -1 0 599300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4361
timestamp 1587416550
transform 0 1 676807 -1 0 599500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4362
timestamp 1587416550
transform 0 1 676807 -1 0 599700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4363
timestamp 1587416550
transform 0 1 676807 -1 0 599900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4364
timestamp 1587416550
transform 0 1 676807 -1 0 600100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4365
timestamp 1587416550
transform 0 1 676807 -1 0 600300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4366
timestamp 1587416550
transform 0 1 676807 -1 0 600500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4368
timestamp 1587416550
transform 0 1 676807 -1 0 600900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4367
timestamp 1587416550
transform 0 1 676807 -1 0 600700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4369
timestamp 1587416550
transform 0 1 676807 -1 0 601100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4371
timestamp 1587416550
transform 0 1 676807 -1 0 601500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4370
timestamp 1587416550
transform 0 1 676807 -1 0 601300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4372
timestamp 1587416550
transform 0 1 676807 -1 0 601700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4373
timestamp 1587416550
transform 0 1 676807 -1 0 601900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4375
timestamp 1587416550
transform 0 1 676807 -1 0 602300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4374
timestamp 1587416550
transform 0 1 676807 -1 0 602100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4376
timestamp 1587416550
transform 0 1 676807 -1 0 602500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4377
timestamp 1587416550
transform 0 1 676807 -1 0 602700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4379
timestamp 1587416550
transform 0 1 676807 -1 0 603100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4378
timestamp 1587416550
transform 0 1 676807 -1 0 602900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4380
timestamp 1587416550
transform 0 1 676807 -1 0 603300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4382
timestamp 1587416550
transform 0 1 676807 -1 0 603700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4381
timestamp 1587416550
transform 0 1 676807 -1 0 603500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4383
timestamp 1587416550
transform 0 1 676807 -1 0 603900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4384
timestamp 1587416550
transform 0 1 676807 -1 0 604100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4386
timestamp 1587416550
transform 0 1 676807 -1 0 604500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4385
timestamp 1587416550
transform 0 1 676807 -1 0 604300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4387
timestamp 1587416550
transform 0 1 676807 -1 0 604700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4389
timestamp 1587416550
transform 0 1 676807 -1 0 605100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4388
timestamp 1587416550
transform 0 1 676807 -1 0 604900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4390
timestamp 1587416550
transform 0 1 676807 -1 0 605300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4391
timestamp 1587416550
transform 0 1 676807 -1 0 605500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4393
timestamp 1587416550
transform 0 1 676807 -1 0 605900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4392
timestamp 1587416550
transform 0 1 676807 -1 0 605700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4394
timestamp 1587416550
transform 0 1 676807 -1 0 606100
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad  gpio_pad[1]
timestamp 1587416550
transform 0 1 676807 -1 0 622100
box -143 -414 16134 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3064
timestamp 1587416550
transform 0 -1 207593 1 0 617100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3065
timestamp 1587416550
transform 0 -1 207593 1 0 617300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3066
timestamp 1587416550
transform 0 -1 207593 1 0 617500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3067
timestamp 1587416550
transform 0 -1 207593 1 0 617700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3068
timestamp 1587416550
transform 0 -1 207593 1 0 617900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3069
timestamp 1587416550
transform 0 -1 207593 1 0 618100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3070
timestamp 1587416550
transform 0 -1 207593 1 0 618300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3071
timestamp 1587416550
transform 0 -1 207593 1 0 618500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3072
timestamp 1587416550
transform 0 -1 207593 1 0 618700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3073
timestamp 1587416550
transform 0 -1 207593 1 0 618900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3074
timestamp 1587416550
transform 0 -1 207593 1 0 619100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3075
timestamp 1587416550
transform 0 -1 207593 1 0 619300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3076
timestamp 1587416550
transform 0 -1 207593 1 0 619500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3077
timestamp 1587416550
transform 0 -1 207593 1 0 619700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3078
timestamp 1587416550
transform 0 -1 207593 1 0 619900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3079
timestamp 1587416550
transform 0 -1 207593 1 0 620100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3080
timestamp 1587416550
transform 0 -1 207593 1 0 620300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3081
timestamp 1587416550
transform 0 -1 207593 1 0 620500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3082
timestamp 1587416550
transform 0 -1 207593 1 0 620700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3083
timestamp 1587416550
transform 0 -1 207593 1 0 620900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3084
timestamp 1587416550
transform 0 -1 207593 1 0 621100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3085
timestamp 1587416550
transform 0 -1 207593 1 0 621300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3086
timestamp 1587416550
transform 0 -1 207593 1 0 621500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3087
timestamp 1587416550
transform 0 -1 207593 1 0 621700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3088
timestamp 1587416550
transform 0 -1 207593 1 0 621900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3089
timestamp 1587416550
transform 0 -1 207593 1 0 622100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3090
timestamp 1587416550
transform 0 -1 207593 1 0 622300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3091
timestamp 1587416550
transform 0 -1 207593 1 0 622500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3092
timestamp 1587416550
transform 0 -1 207593 1 0 622700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3093
timestamp 1587416550
transform 0 -1 207593 1 0 622900
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad  flash_io3_pad
timestamp 1587416550
transform 0 -1 207593 1 0 623100
box -143 -414 16134 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3096
timestamp 1587416550
transform 0 -1 207593 1 0 639300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3095
timestamp 1587416550
transform 0 -1 207593 1 0 639100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3098
timestamp 1587416550
transform 0 -1 207593 1 0 639700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3097
timestamp 1587416550
transform 0 -1 207593 1 0 639500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3100
timestamp 1587416550
transform 0 -1 207593 1 0 640100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3099
timestamp 1587416550
transform 0 -1 207593 1 0 639900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3102
timestamp 1587416550
transform 0 -1 207593 1 0 640500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3101
timestamp 1587416550
transform 0 -1 207593 1 0 640300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3103
timestamp 1587416550
transform 0 -1 207593 1 0 640700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3105
timestamp 1587416550
transform 0 -1 207593 1 0 641100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3104
timestamp 1587416550
transform 0 -1 207593 1 0 640900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3107
timestamp 1587416550
transform 0 -1 207593 1 0 641500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3106
timestamp 1587416550
transform 0 -1 207593 1 0 641300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3109
timestamp 1587416550
transform 0 -1 207593 1 0 641900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3108
timestamp 1587416550
transform 0 -1 207593 1 0 641700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3111
timestamp 1587416550
transform 0 -1 207593 1 0 642300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3110
timestamp 1587416550
transform 0 -1 207593 1 0 642100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3112
timestamp 1587416550
transform 0 -1 207593 1 0 642500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3114
timestamp 1587416550
transform 0 -1 207593 1 0 642900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3113
timestamp 1587416550
transform 0 -1 207593 1 0 642700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3116
timestamp 1587416550
transform 0 -1 207593 1 0 643300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3115
timestamp 1587416550
transform 0 -1 207593 1 0 643100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3118
timestamp 1587416550
transform 0 -1 207593 1 0 643700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3117
timestamp 1587416550
transform 0 -1 207593 1 0 643500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3119
timestamp 1587416550
transform 0 -1 207593 1 0 643900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3121
timestamp 1587416550
transform 0 -1 207593 1 0 644300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3120
timestamp 1587416550
transform 0 -1 207593 1 0 644100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3123
timestamp 1587416550
transform 0 -1 207593 1 0 644700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3122
timestamp 1587416550
transform 0 -1 207593 1 0 644500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3125
timestamp 1587416550
transform 0 -1 207593 1 0 645100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3124
timestamp 1587416550
transform 0 -1 207593 1 0 644900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3127
timestamp 1587416550
transform 0 -1 207593 1 0 645500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3126
timestamp 1587416550
transform 0 -1 207593 1 0 645300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3128
timestamp 1587416550
transform 0 -1 207593 1 0 645700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3130
timestamp 1587416550
transform 0 -1 207593 1 0 646100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3129
timestamp 1587416550
transform 0 -1 207593 1 0 645900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3132
timestamp 1587416550
transform 0 -1 207593 1 0 646500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3131
timestamp 1587416550
transform 0 -1 207593 1 0 646300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3134
timestamp 1587416550
transform 0 -1 207593 1 0 646900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3133
timestamp 1587416550
transform 0 -1 207593 1 0 646700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3135
timestamp 1587416550
transform 0 -1 207593 1 0 647100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3137
timestamp 1587416550
transform 0 -1 207593 1 0 647500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3136
timestamp 1587416550
transform 0 -1 207593 1 0 647300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3139
timestamp 1587416550
transform 0 -1 207593 1 0 647900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3138
timestamp 1587416550
transform 0 -1 207593 1 0 647700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3141
timestamp 1587416550
transform 0 -1 207593 1 0 648300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3140
timestamp 1587416550
transform 0 -1 207593 1 0 648100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3143
timestamp 1587416550
transform 0 -1 207593 1 0 648700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3142
timestamp 1587416550
transform 0 -1 207593 1 0 648500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3144
timestamp 1587416550
transform 0 -1 207593 1 0 648900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3146
timestamp 1587416550
transform 0 -1 207593 1 0 649300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3145
timestamp 1587416550
transform 0 -1 207593 1 0 649100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3148
timestamp 1587416550
transform 0 -1 207593 1 0 649700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3147
timestamp 1587416550
transform 0 -1 207593 1 0 649500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3150
timestamp 1587416550
transform 0 -1 207593 1 0 650100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3149
timestamp 1587416550
transform 0 -1 207593 1 0 649900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3151
timestamp 1587416550
transform 0 -1 207593 1 0 650300
box 0 0 200 39593
use sky130_fd_io__top_gpio_ovtv2  ser_rx_pad /usr/share/pdk/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1587416550
transform 0 -1 208000 1 0 650500
box -80 -88 28211 40076
use sky130_ef_io__com_bus_slice_1um  FILLER_4396
timestamp 1587416550
transform 0 1 676807 -1 0 622300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4397
timestamp 1587416550
transform 0 1 676807 -1 0 622500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4399
timestamp 1587416550
transform 0 1 676807 -1 0 622900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4398
timestamp 1587416550
transform 0 1 676807 -1 0 622700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4400
timestamp 1587416550
transform 0 1 676807 -1 0 623100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4401
timestamp 1587416550
transform 0 1 676807 -1 0 623300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4402
timestamp 1587416550
transform 0 1 676807 -1 0 623500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4403
timestamp 1587416550
transform 0 1 676807 -1 0 623700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4404
timestamp 1587416550
transform 0 1 676807 -1 0 623900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4405
timestamp 1587416550
transform 0 1 676807 -1 0 624100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4406
timestamp 1587416550
transform 0 1 676807 -1 0 624300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4407
timestamp 1587416550
transform 0 1 676807 -1 0 624500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4409
timestamp 1587416550
transform 0 1 676807 -1 0 624900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4408
timestamp 1587416550
transform 0 1 676807 -1 0 624700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4410
timestamp 1587416550
transform 0 1 676807 -1 0 625100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4412
timestamp 1587416550
transform 0 1 676807 -1 0 625500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4411
timestamp 1587416550
transform 0 1 676807 -1 0 625300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4413
timestamp 1587416550
transform 0 1 676807 -1 0 625700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4414
timestamp 1587416550
transform 0 1 676807 -1 0 625900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4415
timestamp 1587416550
transform 0 1 676807 -1 0 626100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4416
timestamp 1587416550
transform 0 1 676807 -1 0 626300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4417
timestamp 1587416550
transform 0 1 676807 -1 0 626500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4418
timestamp 1587416550
transform 0 1 676807 -1 0 626700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4419
timestamp 1587416550
transform 0 1 676807 -1 0 626900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4420
timestamp 1587416550
transform 0 1 676807 -1 0 627100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4421
timestamp 1587416550
transform 0 1 676807 -1 0 627300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4422
timestamp 1587416550
transform 0 1 676807 -1 0 627500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4423
timestamp 1587416550
transform 0 1 676807 -1 0 627700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4424
timestamp 1587416550
transform 0 1 676807 -1 0 627900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4425
timestamp 1587416550
transform 0 1 676807 -1 0 628100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4426
timestamp 1587416550
transform 0 1 676807 -1 0 628300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4428
timestamp 1587416550
transform 0 1 676807 -1 0 628700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4427
timestamp 1587416550
transform 0 1 676807 -1 0 628500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4429
timestamp 1587416550
transform 0 1 676807 -1 0 628900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4430
timestamp 1587416550
transform 0 1 676807 -1 0 629100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4431
timestamp 1587416550
transform 0 1 676807 -1 0 629300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4432
timestamp 1587416550
transform 0 1 676807 -1 0 629500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4433
timestamp 1587416550
transform 0 1 676807 -1 0 629700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4434
timestamp 1587416550
transform 0 1 676807 -1 0 629900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4435
timestamp 1587416550
transform 0 1 676807 -1 0 630100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4436
timestamp 1587416550
transform 0 1 676807 -1 0 630300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4437
timestamp 1587416550
transform 0 1 676807 -1 0 630500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4438
timestamp 1587416550
transform 0 1 676807 -1 0 630700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4439
timestamp 1587416550
transform 0 1 676807 -1 0 630900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4440
timestamp 1587416550
transform 0 1 676807 -1 0 631100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4441
timestamp 1587416550
transform 0 1 676807 -1 0 631300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4442
timestamp 1587416550
transform 0 1 676807 -1 0 631500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4443
timestamp 1587416550
transform 0 1 676807 -1 0 631700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4444
timestamp 1587416550
transform 0 1 676807 -1 0 631900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4445
timestamp 1587416550
transform 0 1 676807 -1 0 632100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4446
timestamp 1587416550
transform 0 1 676807 -1 0 632300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4447
timestamp 1587416550
transform 0 1 676807 -1 0 632500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4448
timestamp 1587416550
transform 0 1 676807 -1 0 632700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4449
timestamp 1587416550
transform 0 1 676807 -1 0 632900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4450
timestamp 1587416550
transform 0 1 676807 -1 0 633100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4451
timestamp 1587416550
transform 0 1 676807 -1 0 633300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4452
timestamp 1587416550
transform 0 1 676807 -1 0 633500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4453
timestamp 1587416550
transform 0 1 676807 -1 0 633700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4454
timestamp 1587416550
transform 0 1 676807 -1 0 633900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4455
timestamp 1587416550
transform 0 1 676807 -1 0 634100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4456
timestamp 1587416550
transform 0 1 676807 -1 0 634300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4457
timestamp 1587416550
transform 0 1 676807 -1 0 634500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4458
timestamp 1587416550
transform 0 1 676807 -1 0 634700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4459
timestamp 1587416550
transform 0 1 676807 -1 0 634900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4460
timestamp 1587416550
transform 0 1 676807 -1 0 635100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4461
timestamp 1587416550
transform 0 1 676807 -1 0 635300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4462
timestamp 1587416550
transform 0 1 676807 -1 0 635500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4463
timestamp 1587416550
transform 0 1 676807 -1 0 635700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4464
timestamp 1587416550
transform 0 1 676807 -1 0 635900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4465
timestamp 1587416550
transform 0 1 676807 -1 0 636100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4466
timestamp 1587416550
transform 0 1 676807 -1 0 636300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4467
timestamp 1587416550
transform 0 1 676807 -1 0 636500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4468
timestamp 1587416550
transform 0 1 676807 -1 0 636700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4469
timestamp 1587416550
transform 0 1 676807 -1 0 636900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4470
timestamp 1587416550
transform 0 1 676807 -1 0 637100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4471
timestamp 1587416550
transform 0 1 676807 -1 0 637300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4472
timestamp 1587416550
transform 0 1 676807 -1 0 637500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4473
timestamp 1587416550
transform 0 1 676807 -1 0 637700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4474
timestamp 1587416550
transform 0 1 676807 -1 0 637900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4475
timestamp 1587416550
transform 0 1 676807 -1 0 638100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4476
timestamp 1587416550
transform 0 1 676807 -1 0 638300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4477
timestamp 1587416550
transform 0 1 676807 -1 0 638500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4478
timestamp 1587416550
transform 0 1 676807 -1 0 638700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4479
timestamp 1587416550
transform 0 1 676807 -1 0 638900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4480
timestamp 1587416550
transform 0 1 676807 -1 0 639100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4481
timestamp 1587416550
transform 0 1 676807 -1 0 639300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4482
timestamp 1587416550
transform 0 1 676807 -1 0 639500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4483
timestamp 1587416550
transform 0 1 676807 -1 0 639700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4484
timestamp 1587416550
transform 0 1 676807 -1 0 639900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4485
timestamp 1587416550
transform 0 1 676807 -1 0 640100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4486
timestamp 1587416550
transform 0 1 676807 -1 0 640300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4487
timestamp 1587416550
transform 0 1 676807 -1 0 640500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4488
timestamp 1587416550
transform 0 1 676807 -1 0 640700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4489
timestamp 1587416550
transform 0 1 676807 -1 0 640900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4490
timestamp 1587416550
transform 0 1 676807 -1 0 641100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4491
timestamp 1587416550
transform 0 1 676807 -1 0 641300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4493
timestamp 1587416550
transform 0 1 676807 -1 0 641700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4492
timestamp 1587416550
transform 0 1 676807 -1 0 641500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4494
timestamp 1587416550
transform 0 1 676807 -1 0 641900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4496
timestamp 1587416550
transform 0 1 676807 -1 0 642300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4495
timestamp 1587416550
transform 0 1 676807 -1 0 642100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4497
timestamp 1587416550
transform 0 1 676807 -1 0 642500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4498
timestamp 1587416550
transform 0 1 676807 -1 0 642700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4500
timestamp 1587416550
transform 0 1 676807 -1 0 643100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4499
timestamp 1587416550
transform 0 1 676807 -1 0 642900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4501
timestamp 1587416550
transform 0 1 676807 -1 0 643300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4502
timestamp 1587416550
transform 0 1 676807 -1 0 643500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4504
timestamp 1587416550
transform 0 1 676807 -1 0 643900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4503
timestamp 1587416550
transform 0 1 676807 -1 0 643700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4505
timestamp 1587416550
transform 0 1 676807 -1 0 644100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4507
timestamp 1587416550
transform 0 1 676807 -1 0 644500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4506
timestamp 1587416550
transform 0 1 676807 -1 0 644300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4508
timestamp 1587416550
transform 0 1 676807 -1 0 644700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4509
timestamp 1587416550
transform 0 1 676807 -1 0 644900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4511
timestamp 1587416550
transform 0 1 676807 -1 0 645300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4510
timestamp 1587416550
transform 0 1 676807 -1 0 645100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4512
timestamp 1587416550
transform 0 1 676807 -1 0 645500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4514
timestamp 1587416550
transform 0 1 676807 -1 0 645900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4513
timestamp 1587416550
transform 0 1 676807 -1 0 645700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4515
timestamp 1587416550
transform 0 1 676807 -1 0 646100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4516
timestamp 1587416550
transform 0 1 676807 -1 0 646300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4518
timestamp 1587416550
transform 0 1 676807 -1 0 646700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4517
timestamp 1587416550
transform 0 1 676807 -1 0 646500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4519
timestamp 1587416550
transform 0 1 676807 -1 0 646900
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad  gpio_pad[0]
timestamp 1587416550
transform 0 1 676807 -1 0 662900
box -143 -414 16134 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3154
timestamp 1587416550
transform 0 -1 207593 1 0 678700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3153
timestamp 1587416550
transform 0 -1 207593 1 0 678500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3156
timestamp 1587416550
transform 0 -1 207593 1 0 679100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3155
timestamp 1587416550
transform 0 -1 207593 1 0 678900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3158
timestamp 1587416550
transform 0 -1 207593 1 0 679500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3157
timestamp 1587416550
transform 0 -1 207593 1 0 679300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3159
timestamp 1587416550
transform 0 -1 207593 1 0 679700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3161
timestamp 1587416550
transform 0 -1 207593 1 0 680100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3160
timestamp 1587416550
transform 0 -1 207593 1 0 679900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3163
timestamp 1587416550
transform 0 -1 207593 1 0 680500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3162
timestamp 1587416550
transform 0 -1 207593 1 0 680300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3165
timestamp 1587416550
transform 0 -1 207593 1 0 680900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3164
timestamp 1587416550
transform 0 -1 207593 1 0 680700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3167
timestamp 1587416550
transform 0 -1 207593 1 0 681300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3166
timestamp 1587416550
transform 0 -1 207593 1 0 681100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3168
timestamp 1587416550
transform 0 -1 207593 1 0 681500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3170
timestamp 1587416550
transform 0 -1 207593 1 0 681900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3169
timestamp 1587416550
transform 0 -1 207593 1 0 681700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3172
timestamp 1587416550
transform 0 -1 207593 1 0 682300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3171
timestamp 1587416550
transform 0 -1 207593 1 0 682100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3174
timestamp 1587416550
transform 0 -1 207593 1 0 682700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3173
timestamp 1587416550
transform 0 -1 207593 1 0 682500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3176
timestamp 1587416550
transform 0 -1 207593 1 0 683100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3175
timestamp 1587416550
transform 0 -1 207593 1 0 682900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3177
timestamp 1587416550
transform 0 -1 207593 1 0 683300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3179
timestamp 1587416550
transform 0 -1 207593 1 0 683700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3178
timestamp 1587416550
transform 0 -1 207593 1 0 683500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3181
timestamp 1587416550
transform 0 -1 207593 1 0 684100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3180
timestamp 1587416550
transform 0 -1 207593 1 0 683900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3183
timestamp 1587416550
transform 0 -1 207593 1 0 684500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3182
timestamp 1587416550
transform 0 -1 207593 1 0 684300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3184
timestamp 1587416550
transform 0 -1 207593 1 0 684700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3186
timestamp 1587416550
transform 0 -1 207593 1 0 685100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3185
timestamp 1587416550
transform 0 -1 207593 1 0 684900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3188
timestamp 1587416550
transform 0 -1 207593 1 0 685500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3187
timestamp 1587416550
transform 0 -1 207593 1 0 685300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3190
timestamp 1587416550
transform 0 -1 207593 1 0 685900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3189
timestamp 1587416550
transform 0 -1 207593 1 0 685700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3192
timestamp 1587416550
transform 0 -1 207593 1 0 686300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3191
timestamp 1587416550
transform 0 -1 207593 1 0 686100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3193
timestamp 1587416550
transform 0 -1 207593 1 0 686500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3195
timestamp 1587416550
transform 0 -1 207593 1 0 686900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3194
timestamp 1587416550
transform 0 -1 207593 1 0 686700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3197
timestamp 1587416550
transform 0 -1 207593 1 0 687300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3196
timestamp 1587416550
transform 0 -1 207593 1 0 687100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3199
timestamp 1587416550
transform 0 -1 207593 1 0 687700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3198
timestamp 1587416550
transform 0 -1 207593 1 0 687500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3201
timestamp 1587416550
transform 0 -1 207593 1 0 688100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3200
timestamp 1587416550
transform 0 -1 207593 1 0 687900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3202
timestamp 1587416550
transform 0 -1 207593 1 0 688300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3204
timestamp 1587416550
transform 0 -1 207593 1 0 688700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3203
timestamp 1587416550
transform 0 -1 207593 1 0 688500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3206
timestamp 1587416550
transform 0 -1 207593 1 0 689100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3205
timestamp 1587416550
transform 0 -1 207593 1 0 688900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3208
timestamp 1587416550
transform 0 -1 207593 1 0 689500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3207
timestamp 1587416550
transform 0 -1 207593 1 0 689300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3209
timestamp 1587416550
transform 0 -1 207593 1 0 689700
box 0 0 200 39593
use sky130_fd_io__top_gpio_ovtv2  ser_tx_pad
timestamp 1587416550
transform 0 -1 208000 1 0 689900
box -80 -88 28211 40076
use sky130_fd_sc_hd__conb_1  mask_rev_value[1]
timestamp 1587416520
transform 1 0 228000 0 1 667085
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1587416520
transform 1 0 228276 0 1 667085
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  mask_rev_value[2]
timestamp 1587416520
transform 1 0 248276 0 1 667085
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value[3]
timestamp 1587416520
transform 1 0 268552 0 1 667085
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1587416520
transform 1 0 248552 0 1 667085
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1587416520
transform 1 0 268828 0 1 667085
box -38 -48 130 592
use striVe_spi  housekeeping
timestamp 1587660775
transform 1 0 288828 0 1 667085
box 0 0 32088 32088
use lvlshiftdown  porb_level_shift
timestamp 1583764616
transform 1 0 340916 0 1 667085
box -66 -23 1986 897
use digital_pll  pll
timestamp 1587660775
transform 1 0 362836 0 1 667085
box 0 0 27735 27735
use sky130_ef_io__com_bus_slice_1um  FILLER_4521
timestamp 1587416550
transform 0 1 676807 -1 0 663100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4522
timestamp 1587416550
transform 0 1 676807 -1 0 663300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4524
timestamp 1587416550
transform 0 1 676807 -1 0 663700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4523
timestamp 1587416550
transform 0 1 676807 -1 0 663500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4525
timestamp 1587416550
transform 0 1 676807 -1 0 663900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4526
timestamp 1587416550
transform 0 1 676807 -1 0 664100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4527
timestamp 1587416550
transform 0 1 676807 -1 0 664300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4528
timestamp 1587416550
transform 0 1 676807 -1 0 664500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4529
timestamp 1587416550
transform 0 1 676807 -1 0 664700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4530
timestamp 1587416550
transform 0 1 676807 -1 0 664900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4531
timestamp 1587416550
transform 0 1 676807 -1 0 665100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4532
timestamp 1587416550
transform 0 1 676807 -1 0 665300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4534
timestamp 1587416550
transform 0 1 676807 -1 0 665700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4533
timestamp 1587416550
transform 0 1 676807 -1 0 665500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4535
timestamp 1587416550
transform 0 1 676807 -1 0 665900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4537
timestamp 1587416550
transform 0 1 676807 -1 0 666300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4536
timestamp 1587416550
transform 0 1 676807 -1 0 666100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4538
timestamp 1587416550
transform 0 1 676807 -1 0 666500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4539
timestamp 1587416550
transform 0 1 676807 -1 0 666700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4540
timestamp 1587416550
transform 0 1 676807 -1 0 666900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4541
timestamp 1587416550
transform 0 1 676807 -1 0 667100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4542
timestamp 1587416550
transform 0 1 676807 -1 0 667300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4543
timestamp 1587416550
transform 0 1 676807 -1 0 667500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4544
timestamp 1587416550
transform 0 1 676807 -1 0 667700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4545
timestamp 1587416550
transform 0 1 676807 -1 0 667900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4546
timestamp 1587416550
transform 0 1 676807 -1 0 668100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4547
timestamp 1587416550
transform 0 1 676807 -1 0 668300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4548
timestamp 1587416550
transform 0 1 676807 -1 0 668500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4549
timestamp 1587416550
transform 0 1 676807 -1 0 668700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4550
timestamp 1587416550
transform 0 1 676807 -1 0 668900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4551
timestamp 1587416550
transform 0 1 676807 -1 0 669100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4553
timestamp 1587416550
transform 0 1 676807 -1 0 669500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4552
timestamp 1587416550
transform 0 1 676807 -1 0 669300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4554
timestamp 1587416550
transform 0 1 676807 -1 0 669700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4555
timestamp 1587416550
transform 0 1 676807 -1 0 669900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4556
timestamp 1587416550
transform 0 1 676807 -1 0 670100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4557
timestamp 1587416550
transform 0 1 676807 -1 0 670300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4558
timestamp 1587416550
transform 0 1 676807 -1 0 670500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4559
timestamp 1587416550
transform 0 1 676807 -1 0 670700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4560
timestamp 1587416550
transform 0 1 676807 -1 0 670900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4561
timestamp 1587416550
transform 0 1 676807 -1 0 671100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4562
timestamp 1587416550
transform 0 1 676807 -1 0 671300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4563
timestamp 1587416550
transform 0 1 676807 -1 0 671500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4564
timestamp 1587416550
transform 0 1 676807 -1 0 671700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4565
timestamp 1587416550
transform 0 1 676807 -1 0 671900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4566
timestamp 1587416550
transform 0 1 676807 -1 0 672100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4567
timestamp 1587416550
transform 0 1 676807 -1 0 672300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4568
timestamp 1587416550
transform 0 1 676807 -1 0 672500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4569
timestamp 1587416550
transform 0 1 676807 -1 0 672700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4570
timestamp 1587416550
transform 0 1 676807 -1 0 672900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4571
timestamp 1587416550
transform 0 1 676807 -1 0 673100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4572
timestamp 1587416550
transform 0 1 676807 -1 0 673300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4573
timestamp 1587416550
transform 0 1 676807 -1 0 673500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4574
timestamp 1587416550
transform 0 1 676807 -1 0 673700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4575
timestamp 1587416550
transform 0 1 676807 -1 0 673900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4576
timestamp 1587416550
transform 0 1 676807 -1 0 674100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4577
timestamp 1587416550
transform 0 1 676807 -1 0 674300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4578
timestamp 1587416550
transform 0 1 676807 -1 0 674500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4579
timestamp 1587416550
transform 0 1 676807 -1 0 674700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4580
timestamp 1587416550
transform 0 1 676807 -1 0 674900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4581
timestamp 1587416550
transform 0 1 676807 -1 0 675100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4582
timestamp 1587416550
transform 0 1 676807 -1 0 675300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4583
timestamp 1587416550
transform 0 1 676807 -1 0 675500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4584
timestamp 1587416550
transform 0 1 676807 -1 0 675700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4585
timestamp 1587416550
transform 0 1 676807 -1 0 675900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4586
timestamp 1587416550
transform 0 1 676807 -1 0 676100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4587
timestamp 1587416550
transform 0 1 676807 -1 0 676300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4588
timestamp 1587416550
transform 0 1 676807 -1 0 676500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4589
timestamp 1587416550
transform 0 1 676807 -1 0 676700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4590
timestamp 1587416550
transform 0 1 676807 -1 0 676900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4591
timestamp 1587416550
transform 0 1 676807 -1 0 677100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4592
timestamp 1587416550
transform 0 1 676807 -1 0 677300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4593
timestamp 1587416550
transform 0 1 676807 -1 0 677500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4594
timestamp 1587416550
transform 0 1 676807 -1 0 677700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4595
timestamp 1587416550
transform 0 1 676807 -1 0 677900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4596
timestamp 1587416550
transform 0 1 676807 -1 0 678100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4597
timestamp 1587416550
transform 0 1 676807 -1 0 678300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4598
timestamp 1587416550
transform 0 1 676807 -1 0 678500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4599
timestamp 1587416550
transform 0 1 676807 -1 0 678700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4600
timestamp 1587416550
transform 0 1 676807 -1 0 678900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4601
timestamp 1587416550
transform 0 1 676807 -1 0 679100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4602
timestamp 1587416550
transform 0 1 676807 -1 0 679300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4603
timestamp 1587416550
transform 0 1 676807 -1 0 679500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4604
timestamp 1587416550
transform 0 1 676807 -1 0 679700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4605
timestamp 1587416550
transform 0 1 676807 -1 0 679900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4606
timestamp 1587416550
transform 0 1 676807 -1 0 680100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4607
timestamp 1587416550
transform 0 1 676807 -1 0 680300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4608
timestamp 1587416550
transform 0 1 676807 -1 0 680500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4609
timestamp 1587416550
transform 0 1 676807 -1 0 680700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4610
timestamp 1587416550
transform 0 1 676807 -1 0 680900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4611
timestamp 1587416550
transform 0 1 676807 -1 0 681100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4612
timestamp 1587416550
transform 0 1 676807 -1 0 681300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4613
timestamp 1587416550
transform 0 1 676807 -1 0 681500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4614
timestamp 1587416550
transform 0 1 676807 -1 0 681700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4615
timestamp 1587416550
transform 0 1 676807 -1 0 681900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4616
timestamp 1587416550
transform 0 1 676807 -1 0 682100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4618
timestamp 1587416550
transform 0 1 676807 -1 0 682500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4617
timestamp 1587416550
transform 0 1 676807 -1 0 682300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4619
timestamp 1587416550
transform 0 1 676807 -1 0 682700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4621
timestamp 1587416550
transform 0 1 676807 -1 0 683100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4620
timestamp 1587416550
transform 0 1 676807 -1 0 682900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4622
timestamp 1587416550
transform 0 1 676807 -1 0 683300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4623
timestamp 1587416550
transform 0 1 676807 -1 0 683500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4625
timestamp 1587416550
transform 0 1 676807 -1 0 683900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4624
timestamp 1587416550
transform 0 1 676807 -1 0 683700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4626
timestamp 1587416550
transform 0 1 676807 -1 0 684100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4627
timestamp 1587416550
transform 0 1 676807 -1 0 684300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4629
timestamp 1587416550
transform 0 1 676807 -1 0 684700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4628
timestamp 1587416550
transform 0 1 676807 -1 0 684500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4630
timestamp 1587416550
transform 0 1 676807 -1 0 684900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4632
timestamp 1587416550
transform 0 1 676807 -1 0 685300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4631
timestamp 1587416550
transform 0 1 676807 -1 0 685100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4633
timestamp 1587416550
transform 0 1 676807 -1 0 685500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4634
timestamp 1587416550
transform 0 1 676807 -1 0 685700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4636
timestamp 1587416550
transform 0 1 676807 -1 0 686100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4635
timestamp 1587416550
transform 0 1 676807 -1 0 685900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4637
timestamp 1587416550
transform 0 1 676807 -1 0 686300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4639
timestamp 1587416550
transform 0 1 676807 -1 0 686700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4638
timestamp 1587416550
transform 0 1 676807 -1 0 686500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4640
timestamp 1587416550
transform 0 1 676807 -1 0 686900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4641
timestamp 1587416550
transform 0 1 676807 -1 0 687100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4643
timestamp 1587416550
transform 0 1 676807 -1 0 687500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4642
timestamp 1587416550
transform 0 1 676807 -1 0 687300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4644
timestamp 1587416550
transform 0 1 676807 -1 0 687700
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad  gpio_pad[11]
timestamp 1587416550
transform 0 1 676807 -1 0 703700
box -143 -414 16134 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3211
timestamp 1587416550
transform 0 -1 207593 1 0 717900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3212
timestamp 1587416550
transform 0 -1 207593 1 0 718100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3213
timestamp 1587416550
transform 0 -1 207593 1 0 718300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3214
timestamp 1587416550
transform 0 -1 207593 1 0 718500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3215
timestamp 1587416550
transform 0 -1 207593 1 0 718700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3216
timestamp 1587416550
transform 0 -1 207593 1 0 718900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3217
timestamp 1587416550
transform 0 -1 207593 1 0 719100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3219
timestamp 1587416550
transform 0 -1 207593 1 0 719500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3218
timestamp 1587416550
transform 0 -1 207593 1 0 719300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3221
timestamp 1587416550
transform 0 -1 207593 1 0 719900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3220
timestamp 1587416550
transform 0 -1 207593 1 0 719700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3223
timestamp 1587416550
transform 0 -1 207593 1 0 720300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3222
timestamp 1587416550
transform 0 -1 207593 1 0 720100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3225
timestamp 1587416550
transform 0 -1 207593 1 0 720700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3224
timestamp 1587416550
transform 0 -1 207593 1 0 720500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3227
timestamp 1587416550
transform 0 -1 207593 1 0 721100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3226
timestamp 1587416550
transform 0 -1 207593 1 0 720900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3229
timestamp 1587416550
transform 0 -1 207593 1 0 721500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3228
timestamp 1587416550
transform 0 -1 207593 1 0 721300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3231
timestamp 1587416550
transform 0 -1 207593 1 0 721900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3230
timestamp 1587416550
transform 0 -1 207593 1 0 721700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3233
timestamp 1587416550
transform 0 -1 207593 1 0 722300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3232
timestamp 1587416550
transform 0 -1 207593 1 0 722100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3235
timestamp 1587416550
transform 0 -1 207593 1 0 722700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3234
timestamp 1587416550
transform 0 -1 207593 1 0 722500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3237
timestamp 1587416550
transform 0 -1 207593 1 0 723100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3236
timestamp 1587416550
transform 0 -1 207593 1 0 722900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3239
timestamp 1587416550
transform 0 -1 207593 1 0 723500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3238
timestamp 1587416550
transform 0 -1 207593 1 0 723300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3241
timestamp 1587416550
transform 0 -1 207593 1 0 723900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3240
timestamp 1587416550
transform 0 -1 207593 1 0 723700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3243
timestamp 1587416550
transform 0 -1 207593 1 0 724300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3242
timestamp 1587416550
transform 0 -1 207593 1 0 724100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3245
timestamp 1587416550
transform 0 -1 207593 1 0 724700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3244
timestamp 1587416550
transform 0 -1 207593 1 0 724500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3247
timestamp 1587416550
transform 0 -1 207593 1 0 725100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3246
timestamp 1587416550
transform 0 -1 207593 1 0 724900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3249
timestamp 1587416550
transform 0 -1 207593 1 0 725500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3248
timestamp 1587416550
transform 0 -1 207593 1 0 725300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3251
timestamp 1587416550
transform 0 -1 207593 1 0 725900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3250
timestamp 1587416550
transform 0 -1 207593 1 0 725700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3253
timestamp 1587416550
transform 0 -1 207593 1 0 726300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3252
timestamp 1587416550
transform 0 -1 207593 1 0 726100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3255
timestamp 1587416550
transform 0 -1 207593 1 0 726700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3254
timestamp 1587416550
transform 0 -1 207593 1 0 726500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3257
timestamp 1587416550
transform 0 -1 207593 1 0 727100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3256
timestamp 1587416550
transform 0 -1 207593 1 0 726900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3259
timestamp 1587416550
transform 0 -1 207593 1 0 727500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3258
timestamp 1587416550
transform 0 -1 207593 1 0 727300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3261
timestamp 1587416550
transform 0 -1 207593 1 0 727900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3260
timestamp 1587416550
transform 0 -1 207593 1 0 727700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3263
timestamp 1587416550
transform 0 -1 207593 1 0 728300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3262
timestamp 1587416550
transform 0 -1 207593 1 0 728100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3265
timestamp 1587416550
transform 0 -1 207593 1 0 728700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3264
timestamp 1587416550
transform 0 -1 207593 1 0 728500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3266
timestamp 1587416550
transform 0 -1 207593 1 0 728900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3268
timestamp 1587416550
transform 0 -1 207593 1 0 729300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_3267
timestamp 1587416550
transform 0 -1 207593 1 0 729100
box 0 0 200 39593
use sky130_ef_io__corner_pad  corner[2]
timestamp 1587416550
transform 0 -1 208800 1 0 729500
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_1um  FILLER_5
timestamp 1587416550
transform 1 0 208800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_6
timestamp 1587416550
transform 1 0 209000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_7
timestamp 1587416550
transform 1 0 209200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_8
timestamp 1587416550
transform 1 0 209400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_9
timestamp 1587416550
transform 1 0 209600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_10
timestamp 1587416550
transform 1 0 209800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_11
timestamp 1587416550
transform 1 0 210000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_12
timestamp 1587416550
transform 1 0 210200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_13
timestamp 1587416550
transform 1 0 210400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_14
timestamp 1587416550
transform 1 0 210600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_15
timestamp 1587416550
transform 1 0 210800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_16
timestamp 1587416550
transform 1 0 211000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_17
timestamp 1587416550
transform 1 0 211200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_18
timestamp 1587416550
transform 1 0 211400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_19
timestamp 1587416550
transform 1 0 211600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_20
timestamp 1587416550
transform 1 0 211800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_21
timestamp 1587416550
transform 1 0 212000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_22
timestamp 1587416550
transform 1 0 212200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_23
timestamp 1587416550
transform 1 0 212400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_24
timestamp 1587416550
transform 1 0 212600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_25
timestamp 1587416550
transform 1 0 212800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_26
timestamp 1587416550
transform 1 0 213000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_27
timestamp 1587416550
transform 1 0 213200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_28
timestamp 1587416550
transform 1 0 213400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_29
timestamp 1587416550
transform 1 0 213600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_30
timestamp 1587416550
transform 1 0 213800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_31
timestamp 1587416550
transform 1 0 214000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_32
timestamp 1587416550
transform 1 0 214200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_34
timestamp 1587416550
transform 1 0 214600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_33
timestamp 1587416550
transform 1 0 214400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_35
timestamp 1587416550
transform 1 0 214800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_36
timestamp 1587416550
transform 1 0 215000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_37
timestamp 1587416550
transform 1 0 215200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_38
timestamp 1587416550
transform 1 0 215400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_39
timestamp 1587416550
transform 1 0 215600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_40
timestamp 1587416550
transform 1 0 215800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_41
timestamp 1587416550
transform 1 0 216000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_42
timestamp 1587416550
transform 1 0 216200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_43
timestamp 1587416550
transform 1 0 216400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_44
timestamp 1587416550
transform 1 0 216600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_45
timestamp 1587416550
transform 1 0 216800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_46
timestamp 1587416550
transform 1 0 217000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_47
timestamp 1587416550
transform 1 0 217200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_48
timestamp 1587416550
transform 1 0 217400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_49
timestamp 1587416550
transform 1 0 217600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_50
timestamp 1587416550
transform 1 0 217800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_51
timestamp 1587416550
transform 1 0 218000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_52
timestamp 1587416550
transform 1 0 218200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_53
timestamp 1587416550
transform 1 0 218400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_54
timestamp 1587416550
transform 1 0 218600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_55
timestamp 1587416550
transform 1 0 218800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_56
timestamp 1587416550
transform 1 0 219000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_57
timestamp 1587416550
transform 1 0 219200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_59
timestamp 1587416550
transform 1 0 219600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_58
timestamp 1587416550
transform 1 0 219400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__vddio_hvc_pad  sky130_ef_io__vddio_hvc_pad_1
timestamp 1587416550
transform 1 0 219800 0 1 729907
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_61
timestamp 1587416550
transform 1 0 234800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_62
timestamp 1587416550
transform 1 0 235000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_63
timestamp 1587416550
transform 1 0 235200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_64
timestamp 1587416550
transform 1 0 235400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_65
timestamp 1587416550
transform 1 0 235600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_66
timestamp 1587416550
transform 1 0 235800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_67
timestamp 1587416550
transform 1 0 236000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_68
timestamp 1587416550
transform 1 0 236200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_69
timestamp 1587416550
transform 1 0 236400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_70
timestamp 1587416550
transform 1 0 236600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_71
timestamp 1587416550
transform 1 0 236800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_72
timestamp 1587416550
transform 1 0 237000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_73
timestamp 1587416550
transform 1 0 237200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_74
timestamp 1587416550
transform 1 0 237400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_75
timestamp 1587416550
transform 1 0 237600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_76
timestamp 1587416550
transform 1 0 237800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_77
timestamp 1587416550
transform 1 0 238000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_78
timestamp 1587416550
transform 1 0 238200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_79
timestamp 1587416550
transform 1 0 238400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_80
timestamp 1587416550
transform 1 0 238600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_81
timestamp 1587416550
transform 1 0 238800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_82
timestamp 1587416550
transform 1 0 239000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_83
timestamp 1587416550
transform 1 0 239200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_84
timestamp 1587416550
transform 1 0 239400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_85
timestamp 1587416550
transform 1 0 239600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_86
timestamp 1587416550
transform 1 0 239800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_87
timestamp 1587416550
transform 1 0 240000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_88
timestamp 1587416550
transform 1 0 240200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_89
timestamp 1587416550
transform 1 0 240400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_90
timestamp 1587416550
transform 1 0 240600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_91
timestamp 1587416550
transform 1 0 240800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_92
timestamp 1587416550
transform 1 0 241000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_93
timestamp 1587416550
transform 1 0 241200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_94
timestamp 1587416550
transform 1 0 241400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_95
timestamp 1587416550
transform 1 0 241600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_96
timestamp 1587416550
transform 1 0 241800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_97
timestamp 1587416550
transform 1 0 242000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_98
timestamp 1587416550
transform 1 0 242200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_99
timestamp 1587416550
transform 1 0 242400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_100
timestamp 1587416550
transform 1 0 242600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_101
timestamp 1587416550
transform 1 0 242800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_102
timestamp 1587416550
transform 1 0 243000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_103
timestamp 1587416550
transform 1 0 243200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_104
timestamp 1587416550
transform 1 0 243400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_105
timestamp 1587416550
transform 1 0 243600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_106
timestamp 1587416550
transform 1 0 243800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_107
timestamp 1587416550
transform 1 0 244000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_108
timestamp 1587416550
transform 1 0 244200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_109
timestamp 1587416550
transform 1 0 244400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_110
timestamp 1587416550
transform 1 0 244600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_111
timestamp 1587416550
transform 1 0 244800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_112
timestamp 1587416550
transform 1 0 245000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_113
timestamp 1587416550
transform 1 0 245200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_114
timestamp 1587416550
transform 1 0 245400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_115
timestamp 1587416550
transform 1 0 245600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_116
timestamp 1587416550
transform 1 0 245800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__vdda_lvc_pad  vdd3v3lclamp[0]
timestamp 1587416550
transform 1 0 246000 0 1 729907
box 0 -7 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_119
timestamp 1587416550
transform 1 0 261200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_118
timestamp 1587416550
transform 1 0 261000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_120
timestamp 1587416550
transform 1 0 261400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_121
timestamp 1587416550
transform 1 0 261600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_122
timestamp 1587416550
transform 1 0 261800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_123
timestamp 1587416550
transform 1 0 262000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_124
timestamp 1587416550
transform 1 0 262200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_125
timestamp 1587416550
transform 1 0 262400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_126
timestamp 1587416550
transform 1 0 262600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_127
timestamp 1587416550
transform 1 0 262800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_128
timestamp 1587416550
transform 1 0 263000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_129
timestamp 1587416550
transform 1 0 263200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_130
timestamp 1587416550
transform 1 0 263400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_131
timestamp 1587416550
transform 1 0 263600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_132
timestamp 1587416550
transform 1 0 263800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_133
timestamp 1587416550
transform 1 0 264000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_134
timestamp 1587416550
transform 1 0 264200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_135
timestamp 1587416550
transform 1 0 264400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_136
timestamp 1587416550
transform 1 0 264600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_137
timestamp 1587416550
transform 1 0 264800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_138
timestamp 1587416550
transform 1 0 265000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_139
timestamp 1587416550
transform 1 0 265200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_140
timestamp 1587416550
transform 1 0 265400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_141
timestamp 1587416550
transform 1 0 265600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_142
timestamp 1587416550
transform 1 0 265800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_143
timestamp 1587416550
transform 1 0 266000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_144
timestamp 1587416550
transform 1 0 266200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_145
timestamp 1587416550
transform 1 0 266400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_146
timestamp 1587416550
transform 1 0 266600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_147
timestamp 1587416550
transform 1 0 266800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_148
timestamp 1587416550
transform 1 0 267000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_149
timestamp 1587416550
transform 1 0 267200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_150
timestamp 1587416550
transform 1 0 267400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_151
timestamp 1587416550
transform 1 0 267600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_152
timestamp 1587416550
transform 1 0 267800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_153
timestamp 1587416550
transform 1 0 268000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_154
timestamp 1587416550
transform 1 0 268200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_155
timestamp 1587416550
transform 1 0 268400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_156
timestamp 1587416550
transform 1 0 268600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_157
timestamp 1587416550
transform 1 0 268800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_158
timestamp 1587416550
transform 1 0 269000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_159
timestamp 1587416550
transform 1 0 269200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_160
timestamp 1587416550
transform 1 0 269400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_161
timestamp 1587416550
transform 1 0 269600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_162
timestamp 1587416550
transform 1 0 269800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_163
timestamp 1587416550
transform 1 0 270000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_164
timestamp 1587416550
transform 1 0 270200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_165
timestamp 1587416550
transform 1 0 270400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_166
timestamp 1587416550
transform 1 0 270600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_167
timestamp 1587416550
transform 1 0 270800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_168
timestamp 1587416550
transform 1 0 271000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_169
timestamp 1587416550
transform 1 0 271200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_170
timestamp 1587416550
transform 1 0 271400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_171
timestamp 1587416550
transform 1 0 271600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_172
timestamp 1587416550
transform 1 0 271800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_173
timestamp 1587416550
transform 1 0 272000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__vccd_hvc_pad  vdd1v8hclamp[0]
timestamp 1587416550
transform 1 0 272200 0 1 729907
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_175
timestamp 1587416550
transform 1 0 287200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_176
timestamp 1587416550
transform 1 0 287400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_177
timestamp 1587416550
transform 1 0 287600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_178
timestamp 1587416550
transform 1 0 287800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_179
timestamp 1587416550
transform 1 0 288000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_180
timestamp 1587416550
transform 1 0 288200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_181
timestamp 1587416550
transform 1 0 288400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_182
timestamp 1587416550
transform 1 0 288600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_183
timestamp 1587416550
transform 1 0 288800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_184
timestamp 1587416550
transform 1 0 289000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_185
timestamp 1587416550
transform 1 0 289200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_186
timestamp 1587416550
transform 1 0 289400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_187
timestamp 1587416550
transform 1 0 289600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_188
timestamp 1587416550
transform 1 0 289800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_189
timestamp 1587416550
transform 1 0 290000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_190
timestamp 1587416550
transform 1 0 290200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_191
timestamp 1587416550
transform 1 0 290400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_192
timestamp 1587416550
transform 1 0 290600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_193
timestamp 1587416550
transform 1 0 290800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_194
timestamp 1587416550
transform 1 0 291000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_195
timestamp 1587416550
transform 1 0 291200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_196
timestamp 1587416550
transform 1 0 291400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_197
timestamp 1587416550
transform 1 0 291600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_198
timestamp 1587416550
transform 1 0 291800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_199
timestamp 1587416550
transform 1 0 292000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_200
timestamp 1587416550
transform 1 0 292200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_201
timestamp 1587416550
transform 1 0 292400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_202
timestamp 1587416550
transform 1 0 292600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_203
timestamp 1587416550
transform 1 0 292800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_204
timestamp 1587416550
transform 1 0 293000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_205
timestamp 1587416550
transform 1 0 293200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_206
timestamp 1587416550
transform 1 0 293400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_207
timestamp 1587416550
transform 1 0 293600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_208
timestamp 1587416550
transform 1 0 293800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_209
timestamp 1587416550
transform 1 0 294000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_210
timestamp 1587416550
transform 1 0 294200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_211
timestamp 1587416550
transform 1 0 294400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_212
timestamp 1587416550
transform 1 0 294600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_213
timestamp 1587416550
transform 1 0 294800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_214
timestamp 1587416550
transform 1 0 295000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_215
timestamp 1587416550
transform 1 0 295200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_216
timestamp 1587416550
transform 1 0 295400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_217
timestamp 1587416550
transform 1 0 295600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_218
timestamp 1587416550
transform 1 0 295800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_219
timestamp 1587416550
transform 1 0 296000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_220
timestamp 1587416550
transform 1 0 296200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_221
timestamp 1587416550
transform 1 0 296400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_222
timestamp 1587416550
transform 1 0 296600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_223
timestamp 1587416550
transform 1 0 296800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_224
timestamp 1587416550
transform 1 0 297000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_225
timestamp 1587416550
transform 1 0 297200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_226
timestamp 1587416550
transform 1 0 297400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_227
timestamp 1587416550
transform 1 0 297600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_228
timestamp 1587416550
transform 1 0 297800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_229
timestamp 1587416550
transform 1 0 298000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__vssa_hvc_pad  vsshclamp[0]
timestamp 1587416550
transform 1 0 298200 0 1 729907
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_231
timestamp 1587416550
transform 1 0 313200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_232
timestamp 1587416550
transform 1 0 313400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_233
timestamp 1587416550
transform 1 0 313600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_235
timestamp 1587416550
transform 1 0 314000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_236
timestamp 1587416550
transform 1 0 314200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_234
timestamp 1587416550
transform 1 0 313800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_237
timestamp 1587416550
transform 1 0 314400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_238
timestamp 1587416550
transform 1 0 314600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_240
timestamp 1587416550
transform 1 0 315000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_239
timestamp 1587416550
transform 1 0 314800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_242
timestamp 1587416550
transform 1 0 315400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_243
timestamp 1587416550
transform 1 0 315600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_241
timestamp 1587416550
transform 1 0 315200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_244
timestamp 1587416550
transform 1 0 315800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_245
timestamp 1587416550
transform 1 0 316000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_246
timestamp 1587416550
transform 1 0 316200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_247
timestamp 1587416550
transform 1 0 316400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_248
timestamp 1587416550
transform 1 0 316600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_249
timestamp 1587416550
transform 1 0 316800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_250
timestamp 1587416550
transform 1 0 317000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_251
timestamp 1587416550
transform 1 0 317200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_252
timestamp 1587416550
transform 1 0 317400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_253
timestamp 1587416550
transform 1 0 317600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_254
timestamp 1587416550
transform 1 0 317800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_255
timestamp 1587416550
transform 1 0 318000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_256
timestamp 1587416550
transform 1 0 318200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_257
timestamp 1587416550
transform 1 0 318400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_258
timestamp 1587416550
transform 1 0 318600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_259
timestamp 1587416550
transform 1 0 318800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_260
timestamp 1587416550
transform 1 0 319000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_261
timestamp 1587416550
transform 1 0 319200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_262
timestamp 1587416550
transform 1 0 319400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_263
timestamp 1587416550
transform 1 0 319600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_264
timestamp 1587416550
transform 1 0 319800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_265
timestamp 1587416550
transform 1 0 320000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_266
timestamp 1587416550
transform 1 0 320200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_267
timestamp 1587416550
transform 1 0 320400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_268
timestamp 1587416550
transform 1 0 320600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_269
timestamp 1587416550
transform 1 0 320800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_270
timestamp 1587416550
transform 1 0 321000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_271
timestamp 1587416550
transform 1 0 321200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_272
timestamp 1587416550
transform 1 0 321400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_273
timestamp 1587416550
transform 1 0 321600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_274
timestamp 1587416550
transform 1 0 321800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_275
timestamp 1587416550
transform 1 0 322000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_276
timestamp 1587416550
transform 1 0 322200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_277
timestamp 1587416550
transform 1 0 322400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_278
timestamp 1587416550
transform 1 0 322600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_279
timestamp 1587416550
transform 1 0 322800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_280
timestamp 1587416550
transform 1 0 323000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_282
timestamp 1587416550
transform 1 0 323400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_281
timestamp 1587416550
transform 1 0 323200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_283
timestamp 1587416550
transform 1 0 323600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_285
timestamp 1587416550
transform 1 0 324000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_284
timestamp 1587416550
transform 1 0 323800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_286
timestamp 1587416550
transform 1 0 324200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__vssd_lvc_pad  sky130_ef_io__vssd_lvc_pad_0 /usr/share/pdk/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1587416550
transform 1 0 324400 0 1 729907
box 0 -7 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_288
timestamp 1587416550
transform 1 0 339400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_289
timestamp 1587416550
transform 1 0 339600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_290
timestamp 1587416550
transform 1 0 339800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_291
timestamp 1587416550
transform 1 0 340000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_292
timestamp 1587416550
transform 1 0 340200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_293
timestamp 1587416550
transform 1 0 340400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_294
timestamp 1587416550
transform 1 0 340600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_296
timestamp 1587416550
transform 1 0 341000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_297
timestamp 1587416550
transform 1 0 341200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_295
timestamp 1587416550
transform 1 0 340800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_298
timestamp 1587416550
transform 1 0 341400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_299
timestamp 1587416550
transform 1 0 341600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_301
timestamp 1587416550
transform 1 0 342000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_300
timestamp 1587416550
transform 1 0 341800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_303
timestamp 1587416550
transform 1 0 342400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_302
timestamp 1587416550
transform 1 0 342200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_304
timestamp 1587416550
transform 1 0 342600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_305
timestamp 1587416550
transform 1 0 342800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_306
timestamp 1587416550
transform 1 0 343000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_307
timestamp 1587416550
transform 1 0 343200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_308
timestamp 1587416550
transform 1 0 343400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_309
timestamp 1587416550
transform 1 0 343600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_310
timestamp 1587416550
transform 1 0 343800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_311
timestamp 1587416550
transform 1 0 344000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_312
timestamp 1587416550
transform 1 0 344200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_313
timestamp 1587416550
transform 1 0 344400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_314
timestamp 1587416550
transform 1 0 344600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_315
timestamp 1587416550
transform 1 0 344800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_316
timestamp 1587416550
transform 1 0 345000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_317
timestamp 1587416550
transform 1 0 345200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_318
timestamp 1587416550
transform 1 0 345400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_319
timestamp 1587416550
transform 1 0 345600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_320
timestamp 1587416550
transform 1 0 345800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_321
timestamp 1587416550
transform 1 0 346000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_322
timestamp 1587416550
transform 1 0 346200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_323
timestamp 1587416550
transform 1 0 346400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_324
timestamp 1587416550
transform 1 0 346600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_325
timestamp 1587416550
transform 1 0 346800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_326
timestamp 1587416550
transform 1 0 347000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_327
timestamp 1587416550
transform 1 0 347200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_328
timestamp 1587416550
transform 1 0 347400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_329
timestamp 1587416550
transform 1 0 347600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_330
timestamp 1587416550
transform 1 0 347800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_331
timestamp 1587416550
transform 1 0 348000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_332
timestamp 1587416550
transform 1 0 348200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_333
timestamp 1587416550
transform 1 0 348400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_334
timestamp 1587416550
transform 1 0 348600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_335
timestamp 1587416550
transform 1 0 348800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_336
timestamp 1587416550
transform 1 0 349000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_337
timestamp 1587416550
transform 1 0 349200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_338
timestamp 1587416550
transform 1 0 349400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_339
timestamp 1587416550
transform 1 0 349600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_340
timestamp 1587416550
transform 1 0 349800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_341
timestamp 1587416550
transform 1 0 350000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_342
timestamp 1587416550
transform 1 0 350200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_343
timestamp 1587416550
transform 1 0 350400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_345
timestamp 1587416550
transform 1 0 366600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_346
timestamp 1587416550
transform 1 0 366800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_347
timestamp 1587416550
transform 1 0 367000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_348
timestamp 1587416550
transform 1 0 367200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad  gpio_pad[8]
timestamp 1587416550
transform 1 0 350600 0 1 729907
box -143 -414 16134 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_349
timestamp 1587416550
transform 1 0 367400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_350
timestamp 1587416550
transform 1 0 367600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_351
timestamp 1587416550
transform 1 0 367800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_352
timestamp 1587416550
transform 1 0 368000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_353
timestamp 1587416550
transform 1 0 368200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_354
timestamp 1587416550
transform 1 0 368400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_355
timestamp 1587416550
transform 1 0 368600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_356
timestamp 1587416550
transform 1 0 368800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_357
timestamp 1587416550
transform 1 0 369000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_358
timestamp 1587416550
transform 1 0 369200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_359
timestamp 1587416550
transform 1 0 369400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_360
timestamp 1587416550
transform 1 0 369600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_361
timestamp 1587416550
transform 1 0 369800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_362
timestamp 1587416550
transform 1 0 370000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_363
timestamp 1587416550
transform 1 0 370200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_364
timestamp 1587416550
transform 1 0 370400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_365
timestamp 1587416550
transform 1 0 370600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_366
timestamp 1587416550
transform 1 0 370800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_367
timestamp 1587416550
transform 1 0 371000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_368
timestamp 1587416550
transform 1 0 371200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_369
timestamp 1587416550
transform 1 0 371400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_370
timestamp 1587416550
transform 1 0 371600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_371
timestamp 1587416550
transform 1 0 371800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_372
timestamp 1587416550
transform 1 0 372000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_373
timestamp 1587416550
transform 1 0 372200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_374
timestamp 1587416550
transform 1 0 372400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_375
timestamp 1587416550
transform 1 0 372600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_376
timestamp 1587416550
transform 1 0 372800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_377
timestamp 1587416550
transform 1 0 373000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_378
timestamp 1587416550
transform 1 0 373200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_379
timestamp 1587416550
transform 1 0 373400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_380
timestamp 1587416550
transform 1 0 373600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_381
timestamp 1587416550
transform 1 0 373800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_382
timestamp 1587416550
transform 1 0 374000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_383
timestamp 1587416550
transform 1 0 374200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_384
timestamp 1587416550
transform 1 0 374400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_385
timestamp 1587416550
transform 1 0 374600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_386
timestamp 1587416550
transform 1 0 374800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_387
timestamp 1587416550
transform 1 0 375000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_388
timestamp 1587416550
transform 1 0 375200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_389
timestamp 1587416550
transform 1 0 375400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_390
timestamp 1587416550
transform 1 0 375600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_391
timestamp 1587416550
transform 1 0 375800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_392
timestamp 1587416550
transform 1 0 376000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_393
timestamp 1587416550
transform 1 0 376200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_394
timestamp 1587416550
transform 1 0 376400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_395
timestamp 1587416550
transform 1 0 376600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_396
timestamp 1587416550
transform 1 0 376800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_397
timestamp 1587416550
transform 1 0 377000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_398
timestamp 1587416550
transform 1 0 377200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_399
timestamp 1587416550
transform 1 0 377400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_400
timestamp 1587416550
transform 1 0 377600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_402
timestamp 1587416550
transform 1 0 393800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_403
timestamp 1587416550
transform 1 0 394000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_404
timestamp 1587416550
transform 1 0 394200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_405
timestamp 1587416550
transform 1 0 394400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_406
timestamp 1587416550
transform 1 0 394600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_407
timestamp 1587416550
transform 1 0 394800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_408
timestamp 1587416550
transform 1 0 395000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_409
timestamp 1587416550
transform 1 0 395200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_410
timestamp 1587416550
transform 1 0 395400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_411
timestamp 1587416550
transform 1 0 395600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_412
timestamp 1587416550
transform 1 0 395800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_413
timestamp 1587416550
transform 1 0 396000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_414
timestamp 1587416550
transform 1 0 396200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_415
timestamp 1587416550
transform 1 0 396400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_416
timestamp 1587416550
transform 1 0 396600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_417
timestamp 1587416550
transform 1 0 396800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_418
timestamp 1587416550
transform 1 0 397000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_419
timestamp 1587416550
transform 1 0 397200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_420
timestamp 1587416550
transform 1 0 397400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_421
timestamp 1587416550
transform 1 0 397600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_422
timestamp 1587416550
transform 1 0 397800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_423
timestamp 1587416550
transform 1 0 398000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_424
timestamp 1587416550
transform 1 0 398200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_425
timestamp 1587416550
transform 1 0 398400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_426
timestamp 1587416550
transform 1 0 398600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_427
timestamp 1587416550
transform 1 0 398800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_428
timestamp 1587416550
transform 1 0 399000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_429
timestamp 1587416550
transform 1 0 399200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_431
timestamp 1587416550
transform 1 0 399600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_430
timestamp 1587416550
transform 1 0 399400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_432
timestamp 1587416550
transform 1 0 399800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_433
timestamp 1587416550
transform 1 0 400000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_434
timestamp 1587416550
transform 1 0 400200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_435
timestamp 1587416550
transform 1 0 400400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_436
timestamp 1587416550
transform 1 0 400600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_437
timestamp 1587416550
transform 1 0 400800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_438
timestamp 1587416550
transform 1 0 401000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_439
timestamp 1587416550
transform 1 0 401200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_440
timestamp 1587416550
transform 1 0 401400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_441
timestamp 1587416550
transform 1 0 401600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_443
timestamp 1587416550
transform 1 0 402000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_442
timestamp 1587416550
transform 1 0 401800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_444
timestamp 1587416550
transform 1 0 402200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_445
timestamp 1587416550
transform 1 0 402400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_446
timestamp 1587416550
transform 1 0 402600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_447
timestamp 1587416550
transform 1 0 402800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_448
timestamp 1587416550
transform 1 0 403000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_450
timestamp 1587416550
transform 1 0 403400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_449
timestamp 1587416550
transform 1 0 403200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_451
timestamp 1587416550
transform 1 0 403600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_453
timestamp 1587416550
transform 1 0 404000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_452
timestamp 1587416550
transform 1 0 403800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_454
timestamp 1587416550
transform 1 0 404200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_456
timestamp 1587416550
transform 1 0 404600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_455
timestamp 1587416550
transform 1 0 404400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad  gpio_pad[7]
timestamp 1587416550
transform 1 0 377800 0 1 729907
box -143 -414 16134 39593
use sky130_ef_io__gpiov2_pad  gpio_pad[6]
timestamp 1587416550
transform 1 0 404800 0 1 729907
box -143 -414 16134 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_458
timestamp 1587416550
transform 1 0 420800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_459
timestamp 1587416550
transform 1 0 421000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_460
timestamp 1587416550
transform 1 0 421200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_461
timestamp 1587416550
transform 1 0 421400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_462
timestamp 1587416550
transform 1 0 421600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_463
timestamp 1587416550
transform 1 0 421800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_464
timestamp 1587416550
transform 1 0 422000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_465
timestamp 1587416550
transform 1 0 422200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_466
timestamp 1587416550
transform 1 0 422400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_468
timestamp 1587416550
transform 1 0 422800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_467
timestamp 1587416550
transform 1 0 422600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_469
timestamp 1587416550
transform 1 0 423000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_470
timestamp 1587416550
transform 1 0 423200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_471
timestamp 1587416550
transform 1 0 423400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_472
timestamp 1587416550
transform 1 0 423600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_473
timestamp 1587416550
transform 1 0 423800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_474
timestamp 1587416550
transform 1 0 424000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_475
timestamp 1587416550
transform 1 0 424200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_476
timestamp 1587416550
transform 1 0 424400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_477
timestamp 1587416550
transform 1 0 424600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_478
timestamp 1587416550
transform 1 0 424800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_479
timestamp 1587416550
transform 1 0 425000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_480
timestamp 1587416550
transform 1 0 425200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_481
timestamp 1587416550
transform 1 0 425400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_482
timestamp 1587416550
transform 1 0 425600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_483
timestamp 1587416550
transform 1 0 425800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_484
timestamp 1587416550
transform 1 0 426000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_485
timestamp 1587416550
transform 1 0 426200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_486
timestamp 1587416550
transform 1 0 426400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_487
timestamp 1587416550
transform 1 0 426600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_488
timestamp 1587416550
transform 1 0 426800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_489
timestamp 1587416550
transform 1 0 427000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_490
timestamp 1587416550
transform 1 0 427200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_491
timestamp 1587416550
transform 1 0 427400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_492
timestamp 1587416550
transform 1 0 427600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_493
timestamp 1587416550
transform 1 0 427800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_494
timestamp 1587416550
transform 1 0 428000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_495
timestamp 1587416550
transform 1 0 428200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_496
timestamp 1587416550
transform 1 0 428400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_497
timestamp 1587416550
transform 1 0 428600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_498
timestamp 1587416550
transform 1 0 428800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_499
timestamp 1587416550
transform 1 0 429000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_500
timestamp 1587416550
transform 1 0 429200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_501
timestamp 1587416550
transform 1 0 429400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_502
timestamp 1587416550
transform 1 0 429600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_503
timestamp 1587416550
transform 1 0 429800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_504
timestamp 1587416550
transform 1 0 430000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_505
timestamp 1587416550
transform 1 0 430200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_506
timestamp 1587416550
transform 1 0 430400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_507
timestamp 1587416550
transform 1 0 430600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_508
timestamp 1587416550
transform 1 0 430800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_509
timestamp 1587416550
transform 1 0 431000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_510
timestamp 1587416550
transform 1 0 431200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_511
timestamp 1587416550
transform 1 0 431400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_512
timestamp 1587416550
transform 1 0 431600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_513
timestamp 1587416550
transform 1 0 431800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_515
timestamp 1587416550
transform 1 0 448000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_516
timestamp 1587416550
transform 1 0 448200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_517
timestamp 1587416550
transform 1 0 448400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_518
timestamp 1587416550
transform 1 0 448600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_519
timestamp 1587416550
transform 1 0 448800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad  gpio_pad[5]
timestamp 1587416550
transform 1 0 432000 0 1 729907
box -143 -414 16134 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_520
timestamp 1587416550
transform 1 0 449000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_521
timestamp 1587416550
transform 1 0 449200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_522
timestamp 1587416550
transform 1 0 449400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_523
timestamp 1587416550
transform 1 0 449600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_524
timestamp 1587416550
transform 1 0 449800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_525
timestamp 1587416550
transform 1 0 450000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_526
timestamp 1587416550
transform 1 0 450200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_527
timestamp 1587416550
transform 1 0 450400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_528
timestamp 1587416550
transform 1 0 450600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_529
timestamp 1587416550
transform 1 0 450800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_530
timestamp 1587416550
transform 1 0 451000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_531
timestamp 1587416550
transform 1 0 451200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_532
timestamp 1587416550
transform 1 0 451400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_533
timestamp 1587416550
transform 1 0 451600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_534
timestamp 1587416550
transform 1 0 451800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_535
timestamp 1587416550
transform 1 0 452000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_536
timestamp 1587416550
transform 1 0 452200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_537
timestamp 1587416550
transform 1 0 452400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_538
timestamp 1587416550
transform 1 0 452600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_539
timestamp 1587416550
transform 1 0 452800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_540
timestamp 1587416550
transform 1 0 453000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_541
timestamp 1587416550
transform 1 0 453200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_542
timestamp 1587416550
transform 1 0 453400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_543
timestamp 1587416550
transform 1 0 453600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_544
timestamp 1587416550
transform 1 0 453800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_545
timestamp 1587416550
transform 1 0 454000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_546
timestamp 1587416550
transform 1 0 454200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_547
timestamp 1587416550
transform 1 0 454400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_548
timestamp 1587416550
transform 1 0 454600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_549
timestamp 1587416550
transform 1 0 454800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_550
timestamp 1587416550
transform 1 0 455000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_551
timestamp 1587416550
transform 1 0 455200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_552
timestamp 1587416550
transform 1 0 455400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_553
timestamp 1587416550
transform 1 0 455600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_554
timestamp 1587416550
transform 1 0 455800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_555
timestamp 1587416550
transform 1 0 456000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_556
timestamp 1587416550
transform 1 0 456200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_557
timestamp 1587416550
transform 1 0 456400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_558
timestamp 1587416550
transform 1 0 456600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_559
timestamp 1587416550
transform 1 0 456800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_560
timestamp 1587416550
transform 1 0 457000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_561
timestamp 1587416550
transform 1 0 457200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_562
timestamp 1587416550
transform 1 0 457400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_563
timestamp 1587416550
transform 1 0 457600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_564
timestamp 1587416550
transform 1 0 457800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_565
timestamp 1587416550
transform 1 0 458000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_566
timestamp 1587416550
transform 1 0 458200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_567
timestamp 1587416550
transform 1 0 458400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_568
timestamp 1587416550
transform 1 0 458600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_569
timestamp 1587416550
transform 1 0 458800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_570
timestamp 1587416550
transform 1 0 459000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_572
timestamp 1587416550
transform 1 0 475200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_573
timestamp 1587416550
transform 1 0 475400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_574
timestamp 1587416550
transform 1 0 475600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_575
timestamp 1587416550
transform 1 0 475800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_576
timestamp 1587416550
transform 1 0 476000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_577
timestamp 1587416550
transform 1 0 476200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_578
timestamp 1587416550
transform 1 0 476400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_579
timestamp 1587416550
transform 1 0 476600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_581
timestamp 1587416550
transform 1 0 477000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_580
timestamp 1587416550
transform 1 0 476800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_582
timestamp 1587416550
transform 1 0 477200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_583
timestamp 1587416550
transform 1 0 477400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_584
timestamp 1587416550
transform 1 0 477600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_585
timestamp 1587416550
transform 1 0 477800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_586
timestamp 1587416550
transform 1 0 478000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_587
timestamp 1587416550
transform 1 0 478200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_588
timestamp 1587416550
transform 1 0 478400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_589
timestamp 1587416550
transform 1 0 478600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_590
timestamp 1587416550
transform 1 0 478800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_591
timestamp 1587416550
transform 1 0 479000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_592
timestamp 1587416550
transform 1 0 479200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_593
timestamp 1587416550
transform 1 0 479400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_594
timestamp 1587416550
transform 1 0 479600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_595
timestamp 1587416550
transform 1 0 479800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_596
timestamp 1587416550
transform 1 0 480000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_597
timestamp 1587416550
transform 1 0 480200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_599
timestamp 1587416550
transform 1 0 480600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_598
timestamp 1587416550
transform 1 0 480400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_600
timestamp 1587416550
transform 1 0 480800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_601
timestamp 1587416550
transform 1 0 481000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_602
timestamp 1587416550
transform 1 0 481200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_603
timestamp 1587416550
transform 1 0 481400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_604
timestamp 1587416550
transform 1 0 481600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_605
timestamp 1587416550
transform 1 0 481800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_606
timestamp 1587416550
transform 1 0 482000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_607
timestamp 1587416550
transform 1 0 482200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_608
timestamp 1587416550
transform 1 0 482400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_609
timestamp 1587416550
transform 1 0 482600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_610
timestamp 1587416550
transform 1 0 482800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_611
timestamp 1587416550
transform 1 0 483000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_612
timestamp 1587416550
transform 1 0 483200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_613
timestamp 1587416550
transform 1 0 483400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_614
timestamp 1587416550
transform 1 0 483600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_616
timestamp 1587416550
transform 1 0 484000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_615
timestamp 1587416550
transform 1 0 483800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_617
timestamp 1587416550
transform 1 0 484200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_619
timestamp 1587416550
transform 1 0 484600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_618
timestamp 1587416550
transform 1 0 484400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_620
timestamp 1587416550
transform 1 0 484800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_622
timestamp 1587416550
transform 1 0 485200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_621
timestamp 1587416550
transform 1 0 485000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_623
timestamp 1587416550
transform 1 0 485400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_625
timestamp 1587416550
transform 1 0 485800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_624
timestamp 1587416550
transform 1 0 485600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_626
timestamp 1587416550
transform 1 0 486000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad  gpio_pad[15]
timestamp 1587416550
transform 1 0 459200 0 1 729907
box -143 -414 16134 39593
use sky130_ef_io__gpiov2_pad  gpio_pad[14]
timestamp 1587416550
transform 1 0 486200 0 1 729907
box -143 -414 16134 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_628
timestamp 1587416550
transform 1 0 502200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_629
timestamp 1587416550
transform 1 0 502400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_630
timestamp 1587416550
transform 1 0 502600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_631
timestamp 1587416550
transform 1 0 502800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_633
timestamp 1587416550
transform 1 0 503200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_632
timestamp 1587416550
transform 1 0 503000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_635
timestamp 1587416550
transform 1 0 503600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_636
timestamp 1587416550
transform 1 0 503800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_634
timestamp 1587416550
transform 1 0 503400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_637
timestamp 1587416550
transform 1 0 504000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_638
timestamp 1587416550
transform 1 0 504200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_639
timestamp 1587416550
transform 1 0 504400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_640
timestamp 1587416550
transform 1 0 504600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_642
timestamp 1587416550
transform 1 0 505000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_641
timestamp 1587416550
transform 1 0 504800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_644
timestamp 1587416550
transform 1 0 505400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_643
timestamp 1587416550
transform 1 0 505200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_645
timestamp 1587416550
transform 1 0 505600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_646
timestamp 1587416550
transform 1 0 505800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_647
timestamp 1587416550
transform 1 0 506000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_648
timestamp 1587416550
transform 1 0 506200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_649
timestamp 1587416550
transform 1 0 506400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_650
timestamp 1587416550
transform 1 0 506600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_651
timestamp 1587416550
transform 1 0 506800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_652
timestamp 1587416550
transform 1 0 507000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_653
timestamp 1587416550
transform 1 0 507200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_654
timestamp 1587416550
transform 1 0 507400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_655
timestamp 1587416550
transform 1 0 507600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_656
timestamp 1587416550
transform 1 0 507800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_657
timestamp 1587416550
transform 1 0 508000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_658
timestamp 1587416550
transform 1 0 508200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_659
timestamp 1587416550
transform 1 0 508400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_660
timestamp 1587416550
transform 1 0 508600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_661
timestamp 1587416550
transform 1 0 508800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_662
timestamp 1587416550
transform 1 0 509000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_663
timestamp 1587416550
transform 1 0 509200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_664
timestamp 1587416550
transform 1 0 509400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_665
timestamp 1587416550
transform 1 0 509600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_666
timestamp 1587416550
transform 1 0 509800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_667
timestamp 1587416550
transform 1 0 510000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_668
timestamp 1587416550
transform 1 0 510200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_669
timestamp 1587416550
transform 1 0 510400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_670
timestamp 1587416550
transform 1 0 510600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_671
timestamp 1587416550
transform 1 0 510800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_672
timestamp 1587416550
transform 1 0 511000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_673
timestamp 1587416550
transform 1 0 511200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_674
timestamp 1587416550
transform 1 0 511400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_675
timestamp 1587416550
transform 1 0 511600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_677
timestamp 1587416550
transform 1 0 512000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_676
timestamp 1587416550
transform 1 0 511800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_678
timestamp 1587416550
transform 1 0 512200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_679
timestamp 1587416550
transform 1 0 512400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_680
timestamp 1587416550
transform 1 0 512600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_681
timestamp 1587416550
transform 1 0 512800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_682
timestamp 1587416550
transform 1 0 513000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_683
timestamp 1587416550
transform 1 0 513200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_685
timestamp 1587416550
transform 1 0 529400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_686
timestamp 1587416550
transform 1 0 529600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_687
timestamp 1587416550
transform 1 0 529800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_688
timestamp 1587416550
transform 1 0 530000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_689
timestamp 1587416550
transform 1 0 530200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_690
timestamp 1587416550
transform 1 0 530400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad  gpio_pad[13]
timestamp 1587416550
transform 1 0 513400 0 1 729907
box -143 -414 16134 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_691
timestamp 1587416550
transform 1 0 530600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_692
timestamp 1587416550
transform 1 0 530800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_693
timestamp 1587416550
transform 1 0 531000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_694
timestamp 1587416550
transform 1 0 531200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_695
timestamp 1587416550
transform 1 0 531400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_696
timestamp 1587416550
transform 1 0 531600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_697
timestamp 1587416550
transform 1 0 531800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_698
timestamp 1587416550
transform 1 0 532000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_699
timestamp 1587416550
transform 1 0 532200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_700
timestamp 1587416550
transform 1 0 532400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_701
timestamp 1587416550
transform 1 0 532600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_702
timestamp 1587416550
transform 1 0 532800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_703
timestamp 1587416550
transform 1 0 533000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_704
timestamp 1587416550
transform 1 0 533200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_705
timestamp 1587416550
transform 1 0 533400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_706
timestamp 1587416550
transform 1 0 533600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_707
timestamp 1587416550
transform 1 0 533800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_708
timestamp 1587416550
transform 1 0 534000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_709
timestamp 1587416550
transform 1 0 534200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_710
timestamp 1587416550
transform 1 0 534400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_711
timestamp 1587416550
transform 1 0 534600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_712
timestamp 1587416550
transform 1 0 534800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_713
timestamp 1587416550
transform 1 0 535000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_714
timestamp 1587416550
transform 1 0 535200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_715
timestamp 1587416550
transform 1 0 535400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_716
timestamp 1587416550
transform 1 0 535600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_717
timestamp 1587416550
transform 1 0 535800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_718
timestamp 1587416550
transform 1 0 536000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_719
timestamp 1587416550
transform 1 0 536200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_720
timestamp 1587416550
transform 1 0 536400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_721
timestamp 1587416550
transform 1 0 536600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_722
timestamp 1587416550
transform 1 0 536800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_723
timestamp 1587416550
transform 1 0 537000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_724
timestamp 1587416550
transform 1 0 537200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_725
timestamp 1587416550
transform 1 0 537400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_726
timestamp 1587416550
transform 1 0 537600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_727
timestamp 1587416550
transform 1 0 537800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_728
timestamp 1587416550
transform 1 0 538000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_729
timestamp 1587416550
transform 1 0 538200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_730
timestamp 1587416550
transform 1 0 538400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_731
timestamp 1587416550
transform 1 0 538600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_732
timestamp 1587416550
transform 1 0 538800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_733
timestamp 1587416550
transform 1 0 539000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_734
timestamp 1587416550
transform 1 0 539200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_735
timestamp 1587416550
transform 1 0 539400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_736
timestamp 1587416550
transform 1 0 539600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_737
timestamp 1587416550
transform 1 0 539800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_738
timestamp 1587416550
transform 1 0 540000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_739
timestamp 1587416550
transform 1 0 540200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_740
timestamp 1587416550
transform 1 0 540400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_742
timestamp 1587416550
transform 1 0 556600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_743
timestamp 1587416550
transform 1 0 556800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_744
timestamp 1587416550
transform 1 0 557000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_745
timestamp 1587416550
transform 1 0 557200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_746
timestamp 1587416550
transform 1 0 557400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_747
timestamp 1587416550
transform 1 0 557600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_748
timestamp 1587416550
transform 1 0 557800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_749
timestamp 1587416550
transform 1 0 558000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_750
timestamp 1587416550
transform 1 0 558200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_751
timestamp 1587416550
transform 1 0 558400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_752
timestamp 1587416550
transform 1 0 558600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_753
timestamp 1587416550
transform 1 0 558800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_754
timestamp 1587416550
transform 1 0 559000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_755
timestamp 1587416550
transform 1 0 559200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_756
timestamp 1587416550
transform 1 0 559400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_757
timestamp 1587416550
transform 1 0 559600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_758
timestamp 1587416550
transform 1 0 559800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_759
timestamp 1587416550
transform 1 0 560000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_760
timestamp 1587416550
transform 1 0 560200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_761
timestamp 1587416550
transform 1 0 560400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_762
timestamp 1587416550
transform 1 0 560600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_763
timestamp 1587416550
transform 1 0 560800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_764
timestamp 1587416550
transform 1 0 561000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_765
timestamp 1587416550
transform 1 0 561200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_766
timestamp 1587416550
transform 1 0 561400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_767
timestamp 1587416550
transform 1 0 561600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_768
timestamp 1587416550
transform 1 0 561800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_769
timestamp 1587416550
transform 1 0 562000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_770
timestamp 1587416550
transform 1 0 562200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_771
timestamp 1587416550
transform 1 0 562400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_772
timestamp 1587416550
transform 1 0 562600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_773
timestamp 1587416550
transform 1 0 562800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_774
timestamp 1587416550
transform 1 0 563000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_775
timestamp 1587416550
transform 1 0 563200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_776
timestamp 1587416550
transform 1 0 563400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_777
timestamp 1587416550
transform 1 0 563600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_778
timestamp 1587416550
transform 1 0 563800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_779
timestamp 1587416550
transform 1 0 564000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_780
timestamp 1587416550
transform 1 0 564200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_782
timestamp 1587416550
transform 1 0 564600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_781
timestamp 1587416550
transform 1 0 564400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_783
timestamp 1587416550
transform 1 0 564800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_784
timestamp 1587416550
transform 1 0 565000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_785
timestamp 1587416550
transform 1 0 565200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_787
timestamp 1587416550
transform 1 0 565600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_786
timestamp 1587416550
transform 1 0 565400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_788
timestamp 1587416550
transform 1 0 565800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_790
timestamp 1587416550
transform 1 0 566200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_789
timestamp 1587416550
transform 1 0 566000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_791
timestamp 1587416550
transform 1 0 566400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_793
timestamp 1587416550
transform 1 0 566800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_792
timestamp 1587416550
transform 1 0 566600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_794
timestamp 1587416550
transform 1 0 567000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_796
timestamp 1587416550
transform 1 0 567400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_795
timestamp 1587416550
transform 1 0 567200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_797
timestamp 1587416550
transform 1 0 567600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad  gpio_pad[12]
timestamp 1587416550
transform 1 0 540600 0 1 729907
box -143 -414 16134 39593
use sky130_ef_io__gpiov2_pad  irq_pad
timestamp 1587416550
transform 1 0 567800 0 1 729907
box -143 -414 16134 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_799
timestamp 1587416550
transform 1 0 583800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_800
timestamp 1587416550
transform 1 0 584000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_801
timestamp 1587416550
transform 1 0 584200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_802
timestamp 1587416550
transform 1 0 584400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_804
timestamp 1587416550
transform 1 0 584800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_803
timestamp 1587416550
transform 1 0 584600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_806
timestamp 1587416550
transform 1 0 585200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_807
timestamp 1587416550
transform 1 0 585400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_805
timestamp 1587416550
transform 1 0 585000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_808
timestamp 1587416550
transform 1 0 585600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_809
timestamp 1587416550
transform 1 0 585800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_810
timestamp 1587416550
transform 1 0 586000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_811
timestamp 1587416550
transform 1 0 586200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_813
timestamp 1587416550
transform 1 0 586600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_812
timestamp 1587416550
transform 1 0 586400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_815
timestamp 1587416550
transform 1 0 587000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_814
timestamp 1587416550
transform 1 0 586800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_816
timestamp 1587416550
transform 1 0 587200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_817
timestamp 1587416550
transform 1 0 587400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_818
timestamp 1587416550
transform 1 0 587600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_819
timestamp 1587416550
transform 1 0 587800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_820
timestamp 1587416550
transform 1 0 588000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_821
timestamp 1587416550
transform 1 0 588200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_822
timestamp 1587416550
transform 1 0 588400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_823
timestamp 1587416550
transform 1 0 588600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_824
timestamp 1587416550
transform 1 0 588800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_825
timestamp 1587416550
transform 1 0 589000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_826
timestamp 1587416550
transform 1 0 589200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_827
timestamp 1587416550
transform 1 0 589400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_828
timestamp 1587416550
transform 1 0 589600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_829
timestamp 1587416550
transform 1 0 589800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_830
timestamp 1587416550
transform 1 0 590000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_831
timestamp 1587416550
transform 1 0 590200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_832
timestamp 1587416550
transform 1 0 590400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_833
timestamp 1587416550
transform 1 0 590600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_834
timestamp 1587416550
transform 1 0 590800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_835
timestamp 1587416550
transform 1 0 591000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_836
timestamp 1587416550
transform 1 0 591200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_837
timestamp 1587416550
transform 1 0 591400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_838
timestamp 1587416550
transform 1 0 591600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_839
timestamp 1587416550
transform 1 0 591800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_840
timestamp 1587416550
transform 1 0 592000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_841
timestamp 1587416550
transform 1 0 592200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_842
timestamp 1587416550
transform 1 0 592400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_843
timestamp 1587416550
transform 1 0 592600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_844
timestamp 1587416550
transform 1 0 592800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_845
timestamp 1587416550
transform 1 0 593000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_846
timestamp 1587416550
transform 1 0 593200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_847
timestamp 1587416550
transform 1 0 593400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_848
timestamp 1587416550
transform 1 0 593600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_849
timestamp 1587416550
transform 1 0 593800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_850
timestamp 1587416550
transform 1 0 594000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_851
timestamp 1587416550
transform 1 0 594200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_852
timestamp 1587416550
transform 1 0 594400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_853
timestamp 1587416550
transform 1 0 594600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_855
timestamp 1587416550
transform 1 0 610800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_856
timestamp 1587416550
transform 1 0 611000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_857
timestamp 1587416550
transform 1 0 611200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_858
timestamp 1587416550
transform 1 0 611400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_859
timestamp 1587416550
transform 1 0 611600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_860
timestamp 1587416550
transform 1 0 611800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_861
timestamp 1587416550
transform 1 0 612000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad  SDO_pad
timestamp 1587416550
transform 1 0 594800 0 1 729907
box -143 -414 16134 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_862
timestamp 1587416550
transform 1 0 612200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_863
timestamp 1587416550
transform 1 0 612400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_864
timestamp 1587416550
transform 1 0 612600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_865
timestamp 1587416550
transform 1 0 612800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_866
timestamp 1587416550
transform 1 0 613000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_867
timestamp 1587416550
transform 1 0 613200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_868
timestamp 1587416550
transform 1 0 613400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_869
timestamp 1587416550
transform 1 0 613600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_870
timestamp 1587416550
transform 1 0 613800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_871
timestamp 1587416550
transform 1 0 614000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_872
timestamp 1587416550
transform 1 0 614200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_873
timestamp 1587416550
transform 1 0 614400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_874
timestamp 1587416550
transform 1 0 614600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_875
timestamp 1587416550
transform 1 0 614800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_876
timestamp 1587416550
transform 1 0 615000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_877
timestamp 1587416550
transform 1 0 615200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_878
timestamp 1587416550
transform 1 0 615400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_879
timestamp 1587416550
transform 1 0 615600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_880
timestamp 1587416550
transform 1 0 615800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_881
timestamp 1587416550
transform 1 0 616000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_882
timestamp 1587416550
transform 1 0 616200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_883
timestamp 1587416550
transform 1 0 616400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_884
timestamp 1587416550
transform 1 0 616600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_885
timestamp 1587416550
transform 1 0 616800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_886
timestamp 1587416550
transform 1 0 617000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_887
timestamp 1587416550
transform 1 0 617200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_888
timestamp 1587416550
transform 1 0 617400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_889
timestamp 1587416550
transform 1 0 617600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_890
timestamp 1587416550
transform 1 0 617800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_891
timestamp 1587416550
transform 1 0 618000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_892
timestamp 1587416550
transform 1 0 618200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_893
timestamp 1587416550
transform 1 0 618400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_894
timestamp 1587416550
transform 1 0 618600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_895
timestamp 1587416550
transform 1 0 618800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_896
timestamp 1587416550
transform 1 0 619000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_897
timestamp 1587416550
transform 1 0 619200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_898
timestamp 1587416550
transform 1 0 619400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_899
timestamp 1587416550
transform 1 0 619600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_900
timestamp 1587416550
transform 1 0 619800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_901
timestamp 1587416550
transform 1 0 620000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_902
timestamp 1587416550
transform 1 0 620200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_903
timestamp 1587416550
transform 1 0 620400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_904
timestamp 1587416550
transform 1 0 620600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_905
timestamp 1587416550
transform 1 0 620800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_906
timestamp 1587416550
transform 1 0 621000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_907
timestamp 1587416550
transform 1 0 621200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_908
timestamp 1587416550
transform 1 0 621400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_909
timestamp 1587416550
transform 1 0 621600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_910
timestamp 1587416550
transform 1 0 621800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_912
timestamp 1587416550
transform 1 0 638000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_913
timestamp 1587416550
transform 1 0 638200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_914
timestamp 1587416550
transform 1 0 638400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_915
timestamp 1587416550
transform 1 0 638600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_916
timestamp 1587416550
transform 1 0 638800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_918
timestamp 1587416550
transform 1 0 639200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_917
timestamp 1587416550
transform 1 0 639000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_919
timestamp 1587416550
transform 1 0 639400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_920
timestamp 1587416550
transform 1 0 639600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_921
timestamp 1587416550
transform 1 0 639800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_923
timestamp 1587416550
transform 1 0 640200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_922
timestamp 1587416550
transform 1 0 640000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_924
timestamp 1587416550
transform 1 0 640400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_925
timestamp 1587416550
transform 1 0 640600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_926
timestamp 1587416550
transform 1 0 640800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_927
timestamp 1587416550
transform 1 0 641000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_928
timestamp 1587416550
transform 1 0 641200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_929
timestamp 1587416550
transform 1 0 641400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_930
timestamp 1587416550
transform 1 0 641600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_931
timestamp 1587416550
transform 1 0 641800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_932
timestamp 1587416550
transform 1 0 642000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_933
timestamp 1587416550
transform 1 0 642200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_934
timestamp 1587416550
transform 1 0 642400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_935
timestamp 1587416550
transform 1 0 642600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_936
timestamp 1587416550
transform 1 0 642800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_937
timestamp 1587416550
transform 1 0 643000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_938
timestamp 1587416550
transform 1 0 643200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_939
timestamp 1587416550
transform 1 0 643400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_940
timestamp 1587416550
transform 1 0 643600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_941
timestamp 1587416550
transform 1 0 643800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_942
timestamp 1587416550
transform 1 0 644000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_943
timestamp 1587416550
transform 1 0 644200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_944
timestamp 1587416550
transform 1 0 644400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_945
timestamp 1587416550
transform 1 0 644600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_946
timestamp 1587416550
transform 1 0 644800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_947
timestamp 1587416550
transform 1 0 645000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_948
timestamp 1587416550
transform 1 0 645200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_949
timestamp 1587416550
transform 1 0 645400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_950
timestamp 1587416550
transform 1 0 645600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_951
timestamp 1587416550
transform 1 0 645800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_952
timestamp 1587416550
transform 1 0 646000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_953
timestamp 1587416550
transform 1 0 646200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_954
timestamp 1587416550
transform 1 0 646400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_955
timestamp 1587416550
transform 1 0 646600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_956
timestamp 1587416550
transform 1 0 646800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_957
timestamp 1587416550
transform 1 0 647000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_958
timestamp 1587416550
transform 1 0 647200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_959
timestamp 1587416550
transform 1 0 647400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_960
timestamp 1587416550
transform 1 0 647600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_961
timestamp 1587416550
transform 1 0 647800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_963
timestamp 1587416550
transform 1 0 648200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_962
timestamp 1587416550
transform 1 0 648000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_965
timestamp 1587416550
transform 1 0 648600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_964
timestamp 1587416550
transform 1 0 648400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_966
timestamp 1587416550
transform 1 0 648800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_967
timestamp 1587416550
transform 1 0 649000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad  SDI_pad
timestamp 1587416550
transform 1 0 622000 0 1 729907
box -143 -414 16134 39593
use sky130_ef_io__gpiov2_pad  flash_csb_pad
timestamp 1587416550
transform 1 0 649200 0 1 729907
box -143 -414 16134 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4646
timestamp 1587416550
transform 0 1 676807 -1 0 703900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4647
timestamp 1587416550
transform 0 1 676807 -1 0 704100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4649
timestamp 1587416550
transform 0 1 676807 -1 0 704500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4648
timestamp 1587416550
transform 0 1 676807 -1 0 704300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4650
timestamp 1587416550
transform 0 1 676807 -1 0 704700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4651
timestamp 1587416550
transform 0 1 676807 -1 0 704900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4653
timestamp 1587416550
transform 0 1 676807 -1 0 705300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4652
timestamp 1587416550
transform 0 1 676807 -1 0 705100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4654
timestamp 1587416550
transform 0 1 676807 -1 0 705500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4655
timestamp 1587416550
transform 0 1 676807 -1 0 705700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4656
timestamp 1587416550
transform 0 1 676807 -1 0 705900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4658
timestamp 1587416550
transform 0 1 676807 -1 0 706300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4657
timestamp 1587416550
transform 0 1 676807 -1 0 706100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4659
timestamp 1587416550
transform 0 1 676807 -1 0 706500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4660
timestamp 1587416550
transform 0 1 676807 -1 0 706700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4662
timestamp 1587416550
transform 0 1 676807 -1 0 707100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4661
timestamp 1587416550
transform 0 1 676807 -1 0 706900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4663
timestamp 1587416550
transform 0 1 676807 -1 0 707300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4664
timestamp 1587416550
transform 0 1 676807 -1 0 707500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4666
timestamp 1587416550
transform 0 1 676807 -1 0 707900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4665
timestamp 1587416550
transform 0 1 676807 -1 0 707700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4667
timestamp 1587416550
transform 0 1 676807 -1 0 708100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4668
timestamp 1587416550
transform 0 1 676807 -1 0 708300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4670
timestamp 1587416550
transform 0 1 676807 -1 0 708700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4669
timestamp 1587416550
transform 0 1 676807 -1 0 708500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4671
timestamp 1587416550
transform 0 1 676807 -1 0 708900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4672
timestamp 1587416550
transform 0 1 676807 -1 0 709100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4674
timestamp 1587416550
transform 0 1 676807 -1 0 709500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4673
timestamp 1587416550
transform 0 1 676807 -1 0 709300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4675
timestamp 1587416550
transform 0 1 676807 -1 0 709700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4676
timestamp 1587416550
transform 0 1 676807 -1 0 709900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4678
timestamp 1587416550
transform 0 1 676807 -1 0 710300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4677
timestamp 1587416550
transform 0 1 676807 -1 0 710100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4679
timestamp 1587416550
transform 0 1 676807 -1 0 710500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4680
timestamp 1587416550
transform 0 1 676807 -1 0 710700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4682
timestamp 1587416550
transform 0 1 676807 -1 0 711100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4681
timestamp 1587416550
transform 0 1 676807 -1 0 710900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4683
timestamp 1587416550
transform 0 1 676807 -1 0 711300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4684
timestamp 1587416550
transform 0 1 676807 -1 0 711500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4686
timestamp 1587416550
transform 0 1 676807 -1 0 711900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4685
timestamp 1587416550
transform 0 1 676807 -1 0 711700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4687
timestamp 1587416550
transform 0 1 676807 -1 0 712100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4688
timestamp 1587416550
transform 0 1 676807 -1 0 712300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4689
timestamp 1587416550
transform 0 1 676807 -1 0 712500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4691
timestamp 1587416550
transform 0 1 676807 -1 0 712900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4690
timestamp 1587416550
transform 0 1 676807 -1 0 712700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4692
timestamp 1587416550
transform 0 1 676807 -1 0 713100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4693
timestamp 1587416550
transform 0 1 676807 -1 0 713300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4695
timestamp 1587416550
transform 0 1 676807 -1 0 713700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4694
timestamp 1587416550
transform 0 1 676807 -1 0 713500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4696
timestamp 1587416550
transform 0 1 676807 -1 0 713900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4697
timestamp 1587416550
transform 0 1 676807 -1 0 714100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4699
timestamp 1587416550
transform 0 1 676807 -1 0 714500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4698
timestamp 1587416550
transform 0 1 676807 -1 0 714300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4700
timestamp 1587416550
transform 0 1 676807 -1 0 714700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4701
timestamp 1587416550
transform 0 1 676807 -1 0 714900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4703
timestamp 1587416550
transform 0 1 676807 -1 0 715300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4702
timestamp 1587416550
transform 0 1 676807 -1 0 715100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4704
timestamp 1587416550
transform 0 1 676807 -1 0 715500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4705
timestamp 1587416550
transform 0 1 676807 -1 0 715700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4707
timestamp 1587416550
transform 0 1 676807 -1 0 716100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4706
timestamp 1587416550
transform 0 1 676807 -1 0 715900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4708
timestamp 1587416550
transform 0 1 676807 -1 0 716300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4709
timestamp 1587416550
transform 0 1 676807 -1 0 716500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4711
timestamp 1587416550
transform 0 1 676807 -1 0 716900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4710
timestamp 1587416550
transform 0 1 676807 -1 0 716700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4712
timestamp 1587416550
transform 0 1 676807 -1 0 717100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4713
timestamp 1587416550
transform 0 1 676807 -1 0 717300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4715
timestamp 1587416550
transform 0 1 676807 -1 0 717700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4714
timestamp 1587416550
transform 0 1 676807 -1 0 717500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4716
timestamp 1587416550
transform 0 1 676807 -1 0 717900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4717
timestamp 1587416550
transform 0 1 676807 -1 0 718100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4719
timestamp 1587416550
transform 0 1 676807 -1 0 718500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4718
timestamp 1587416550
transform 0 1 676807 -1 0 718300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4720
timestamp 1587416550
transform 0 1 676807 -1 0 718700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4721
timestamp 1587416550
transform 0 1 676807 -1 0 718900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4722
timestamp 1587416550
transform 0 1 676807 -1 0 719100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4724
timestamp 1587416550
transform 0 1 676807 -1 0 719500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4723
timestamp 1587416550
transform 0 1 676807 -1 0 719300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4726
timestamp 1587416550
transform 0 1 676807 -1 0 719900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4725
timestamp 1587416550
transform 0 1 676807 -1 0 719700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4728
timestamp 1587416550
transform 0 1 676807 -1 0 720300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4727
timestamp 1587416550
transform 0 1 676807 -1 0 720100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4730
timestamp 1587416550
transform 0 1 676807 -1 0 720700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4729
timestamp 1587416550
transform 0 1 676807 -1 0 720500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4732
timestamp 1587416550
transform 0 1 676807 -1 0 721100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4731
timestamp 1587416550
transform 0 1 676807 -1 0 720900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4734
timestamp 1587416550
transform 0 1 676807 -1 0 721500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4733
timestamp 1587416550
transform 0 1 676807 -1 0 721300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4736
timestamp 1587416550
transform 0 1 676807 -1 0 721900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4735
timestamp 1587416550
transform 0 1 676807 -1 0 721700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4739
timestamp 1587416550
transform 0 1 676807 -1 0 722500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4738
timestamp 1587416550
transform 0 1 676807 -1 0 722300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4737
timestamp 1587416550
transform 0 1 676807 -1 0 722100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4741
timestamp 1587416550
transform 0 1 676807 -1 0 722900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4740
timestamp 1587416550
transform 0 1 676807 -1 0 722700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4743
timestamp 1587416550
transform 0 1 676807 -1 0 723300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4742
timestamp 1587416550
transform 0 1 676807 -1 0 723100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4745
timestamp 1587416550
transform 0 1 676807 -1 0 723700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4744
timestamp 1587416550
transform 0 1 676807 -1 0 723500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4747
timestamp 1587416550
transform 0 1 676807 -1 0 724100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4746
timestamp 1587416550
transform 0 1 676807 -1 0 723900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4749
timestamp 1587416550
transform 0 1 676807 -1 0 724500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4748
timestamp 1587416550
transform 0 1 676807 -1 0 724300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4751
timestamp 1587416550
transform 0 1 676807 -1 0 724900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4750
timestamp 1587416550
transform 0 1 676807 -1 0 724700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4753
timestamp 1587416550
transform 0 1 676807 -1 0 725300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4752
timestamp 1587416550
transform 0 1 676807 -1 0 725100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4756
timestamp 1587416550
transform 0 1 676807 -1 0 725900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4755
timestamp 1587416550
transform 0 1 676807 -1 0 725700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4754
timestamp 1587416550
transform 0 1 676807 -1 0 725500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4758
timestamp 1587416550
transform 0 1 676807 -1 0 726300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4757
timestamp 1587416550
transform 0 1 676807 -1 0 726100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4760
timestamp 1587416550
transform 0 1 676807 -1 0 726700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4759
timestamp 1587416550
transform 0 1 676807 -1 0 726500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4762
timestamp 1587416550
transform 0 1 676807 -1 0 727100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4761
timestamp 1587416550
transform 0 1 676807 -1 0 726900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4764
timestamp 1587416550
transform 0 1 676807 -1 0 727500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4763
timestamp 1587416550
transform 0 1 676807 -1 0 727300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4766
timestamp 1587416550
transform 0 1 676807 -1 0 727900
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4765
timestamp 1587416550
transform 0 1 676807 -1 0 727700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4768
timestamp 1587416550
transform 0 1 676807 -1 0 728300
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4767
timestamp 1587416550
transform 0 1 676807 -1 0 728100
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4770
timestamp 1587416550
transform 0 1 676807 -1 0 728700
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_4769
timestamp 1587416550
transform 0 1 676807 -1 0 728500
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_969
timestamp 1587416550
transform 1 0 665200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_970
timestamp 1587416550
transform 1 0 665400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_971
timestamp 1587416550
transform 1 0 665600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_972
timestamp 1587416550
transform 1 0 665800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_973
timestamp 1587416550
transform 1 0 666000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_974
timestamp 1587416550
transform 1 0 666200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_975
timestamp 1587416550
transform 1 0 666400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_976
timestamp 1587416550
transform 1 0 666600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_977
timestamp 1587416550
transform 1 0 666800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_978
timestamp 1587416550
transform 1 0 667000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_979
timestamp 1587416550
transform 1 0 667200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_980
timestamp 1587416550
transform 1 0 667400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_981
timestamp 1587416550
transform 1 0 667600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_982
timestamp 1587416550
transform 1 0 667800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_983
timestamp 1587416550
transform 1 0 668000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_984
timestamp 1587416550
transform 1 0 668200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_985
timestamp 1587416550
transform 1 0 668400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_986
timestamp 1587416550
transform 1 0 668600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_987
timestamp 1587416550
transform 1 0 668800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_988
timestamp 1587416550
transform 1 0 669000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_989
timestamp 1587416550
transform 1 0 669200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_990
timestamp 1587416550
transform 1 0 669400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_991
timestamp 1587416550
transform 1 0 669600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_992
timestamp 1587416550
transform 1 0 669800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_993
timestamp 1587416550
transform 1 0 670000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_994
timestamp 1587416550
transform 1 0 670200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_995
timestamp 1587416550
transform 1 0 670400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_996
timestamp 1587416550
transform 1 0 670600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_997
timestamp 1587416550
transform 1 0 670800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_998
timestamp 1587416550
transform 1 0 671000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_999
timestamp 1587416550
transform 1 0 671200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1000
timestamp 1587416550
transform 1 0 671400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1001
timestamp 1587416550
transform 1 0 671600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1002
timestamp 1587416550
transform 1 0 671800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1003
timestamp 1587416550
transform 1 0 672000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1004
timestamp 1587416550
transform 1 0 672200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1005
timestamp 1587416550
transform 1 0 672400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1006
timestamp 1587416550
transform 1 0 672600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1007
timestamp 1587416550
transform 1 0 672800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1008
timestamp 1587416550
transform 1 0 673000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1009
timestamp 1587416550
transform 1 0 673200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1010
timestamp 1587416550
transform 1 0 673400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1011
timestamp 1587416550
transform 1 0 673600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1012
timestamp 1587416550
transform 1 0 673800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1013
timestamp 1587416550
transform 1 0 674000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1014
timestamp 1587416550
transform 1 0 674200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1015
timestamp 1587416550
transform 1 0 674400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1016
timestamp 1587416550
transform 1 0 674600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1017
timestamp 1587416550
transform 1 0 674800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1018
timestamp 1587416550
transform 1 0 675000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1019
timestamp 1587416550
transform 1 0 675200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1020
timestamp 1587416550
transform 1 0 675400 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1021
timestamp 1587416550
transform 1 0 675600 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1022
timestamp 1587416550
transform 1 0 675800 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1023
timestamp 1587416550
transform 1 0 676000 0 1 729907
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_1024
timestamp 1587416550
transform 1 0 676200 0 1 729907
box 0 0 200 39593
use sky130_ef_io__corner_pad  corner[3]
timestamp 1587416550
transform 1 0 676400 0 1 728700
box 0 0 40000 40800
use advSeal_6um_gen  advSeal_6um_gen_0
timestamp 1584566829
transform 1 0 0 0 1 0
box 0 0 886000 989000
<< labels >>
flabel metal5 s 175734 273638 185752 284112 0 FreeSans 16000 0 0 0 vdd
port 0 nsew
flabel metal5 s 176136 353254 186152 363328 0 FreeSans 16000 0 0 0 vss
port 1 nsew
flabel metal5 s 175906 380556 185408 390630 0 FreeSans 16000 0 0 0 comp_inp
port 2 nsew
flabel metal5 s 175964 409004 185350 414956 0 FreeSans 16000 0 0 0 RSTB
port 3 nsew
flabel metal5 s 175850 434588 185350 444490 0 FreeSans 16000 0 0 0 CSB
port 4 nsew
flabel metal5 s 175734 461604 185694 472078 0 FreeSans 16000 0 0 0 SCK
port 5 nsew
flabel metal5 s 176078 489650 185408 499380 0 FreeSans 16000 0 0 0 xclk
port 6 nsew
flabel metal5 s 176308 516722 185122 526796 0 FreeSans 16000 0 0 0 flash_clk
port 7 nsew
flabel metal5 s 176250 544310 185464 554328 0 FreeSans 16000 0 0 0 flash_io0
port 8 nsew
flabel metal5 s 176078 571440 185580 581572 0 FreeSans 16000 0 0 0 flash_io1
port 9 nsew
flabel metal5 s 176136 599200 185752 608988 0 FreeSans 16000 0 0 0 flash_io2
port 10 nsew
flabel metal5 s 175850 626618 185350 636748 0 FreeSans 16000 0 0 0 flash_io3
port 11 nsew
flabel metal5 s 176536 655006 183462 666168 0 FreeSans 16000 0 0 0 ser_rx
port 12 nsew
flabel metal5 s 176764 694556 183634 705776 0 FreeSans 16000 0 0 0 ser_tx
port 13 nsew
flabel metal5 s 354142 751394 363700 761868 0 FreeSans 16000 0 0 0 gpio[8]
port 14 nsew
flabel metal5 s 381786 751908 390716 761524 0 FreeSans 16000 0 0 0 gpio[7]
port 15 nsew
flabel metal5 s 408058 751850 417732 760894 0 FreeSans 16000 0 0 0 gpio[6]
port 16 nsew
flabel metal5 s 435532 751850 445662 761810 0 FreeSans 16000 0 0 0 gpio[5]
port 17 nsew
flabel metal5 s 462948 751794 472736 761238 0 FreeSans 16000 0 0 0 gpio[15]
port 18 nsew
flabel metal5 s 489620 751850 499752 761524 0 FreeSans 16000 0 0 0 gpio[14]
port 19 nsew
flabel metal5 s 517324 751736 526138 761638 0 FreeSans 16000 0 0 0 gpio[13]
port 20 nsew
flabel metal5 s 544510 751450 553554 761238 0 FreeSans 16000 0 0 0 gpio[12]
port 21 nsew
flabel metal5 s 571640 752022 580798 761466 0 FreeSans 16000 0 0 0 irq
port 22 nsew
flabel metal5 s 598428 752022 607814 761638 0 FreeSans 16000 0 0 0 SDO
port 23 nsew
flabel metal5 s 625328 751794 634486 761066 0 FreeSans 16000 0 0 0 SDI
port 24 nsew
flabel metal5 s 653146 751966 662590 761696 0 FreeSans 16000 0 0 0 flash_csb
port 25 nsew
flabel metal5 s 699050 690206 707864 699822 0 FreeSans 16000 0 0 0 gpio[11]
port 26 nsew
flabel metal5 s 698534 649626 708436 659242 0 FreeSans 16000 0 0 0 gpio[0]
port 27 nsew
flabel metal5 s 698420 608530 708894 619062 0 FreeSans 16000 0 0 0 gpio[1]
port 28 nsew
flabel metal5 s 698362 568236 708722 578080 0 FreeSans 16000 0 0 0 gpio[2]
port 29 nsew
flabel metal5 s 698192 526682 708436 536412 0 FreeSans 16000 0 0 0 gpio[3]
port 30 nsew
flabel metal5 s 699336 486388 708494 495488 0 FreeSans 16000 0 0 0 gpio[4]
port 31 nsew
flabel metal5 s 645590 227334 654978 236950 0 FreeSans 16000 0 0 0 gpio[9]
port 32 nsew
flabel metal5 s 613882 227562 622180 236892 0 FreeSans 16000 0 0 0 gpio[10]
port 33 nsew
flabel metal5 s 580398 227048 589498 237006 0 FreeSans 16000 0 0 0 xi
port 34 nsew
flabel metal5 s 547658 227276 557618 237064 0 FreeSans 16000 0 0 0 xo
port 35 nsew
flabel metal5 s 515606 227048 524364 237122 0 FreeSans 16000 0 0 0 adc0_in
port 36 nsew
flabel metal5 s 483038 227276 492140 237178 0 FreeSans 16000 0 0 0 adc1_in
port 37 nsew
flabel metal5 s 450356 227220 459456 237294 0 FreeSans 16000 0 0 0 adc_high
port 38 nsew
flabel metal5 s 417502 226934 427004 236664 0 FreeSans 16000 0 0 0 adc_low
port 39 nsew
flabel metal5 s 385050 227620 394952 237064 0 FreeSans 16000 0 0 0 comp_inn
port 40 nsew
flabel metal5 s 291182 227048 298794 237464 0 FreeSans 16000 0 0 0 vdd1v8
port 41 nsew
flabel metal5 253032 711304 253032 711304 0 FreeSans 12800 0 0 0 vdd1v8
flabel metal5 226440 654050 226440 654050 0 FreeSans 12800 0 0 0 vss
flabel metal4 239546 277776 239546 277776 0 FreeSans 12800 0 0 0 vss
flabel metal5 226196 268268 226196 268268 0 FreeSans 12800 0 0 0 vdd1v8
flabel metal4 645492 290158 645492 290158 0 FreeSans 12800 0 0 0 vss
flabel metal4 632358 697894 632358 697894 0 FreeSans 12800 0 0 0 vdd1v8
<< end >>
