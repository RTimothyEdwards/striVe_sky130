VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO digital_pll
  CLASS BLOCK ;
  FOREIGN digital_pll ;
  ORIGIN 0.000 0.000 ;
  SIZE 138.675 BY 138.675 ;
  PIN reset
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.920 0.000 82.620 2.100 ;
    END
  END reset
  PIN extclk_sel
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.880 0.000 2.580 2.100 ;
    END
  END extclk_sel
  PIN osc
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 136.515 113.110 138.675 114.610 ;
    END
  END osc
  PIN clockc
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.910 2.160 121.410 ;
    END
  END clockc
  PIN clockp[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 122.400 0.000 123.100 2.100 ;
    END
  END clockp[1]
  PIN clockp[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 136.515 83.190 138.675 84.690 ;
    END
  END clockp[0]
  PIN clockd[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 31.320 136.575 32.020 138.675 ;
    END
  END clockd[3]
  PIN clockd[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.190 2.160 16.690 ;
    END
  END clockd[2]
  PIN clockd[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 136.515 128.070 138.675 129.570 ;
    END
  END clockd[1]
  PIN clockd[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 136.515 53.270 138.675 54.770 ;
    END
  END clockd[0]
  PIN div[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 136.515 68.230 138.675 69.730 ;
    END
  END div[4]
  PIN div[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.080 136.575 11.780 138.675 ;
    END
  END div[3]
  PIN div[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.030 2.160 76.530 ;
    END
  END div[2]
  PIN div[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 132.520 0.000 133.220 2.100 ;
    END
  END div[1]
  PIN div[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.200 136.575 21.900 138.675 ;
    END
  END div[0]
  PIN sel[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 102.160 0.000 102.860 2.100 ;
    END
  END sel[2]
  PIN sel[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 92.040 0.000 92.740 2.100 ;
    END
  END sel[1]
  PIN sel[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 136.515 9.750 138.675 11.250 ;
    END
  END sel[0]
  PIN dco
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.440 0.000 42.140 2.100 ;
    END
  END dco
  PIN ext_trim[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.110 2.160 46.610 ;
    END
  END ext_trim[25]
  PIN ext_trim[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 112.280 0.000 112.980 2.100 ;
    END
  END ext_trim[24]
  PIN ext_trim[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 136.515 98.150 138.675 99.650 ;
    END
  END ext_trim[23]
  PIN ext_trim[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.070 2.160 61.570 ;
    END
  END ext_trim[22]
  PIN ext_trim[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.870 2.160 136.370 ;
    END
  END ext_trim[21]
  PIN ext_trim[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.080 0.000 11.780 2.100 ;
    END
  END ext_trim[20]
  PIN ext_trim[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.200 0.000 21.900 2.100 ;
    END
  END ext_trim[19]
  PIN ext_trim[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.800 0.000 72.500 2.100 ;
    END
  END ext_trim[18]
  PIN ext_trim[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.560 0.000 52.260 2.100 ;
    END
  END ext_trim[17]
  PIN ext_trim[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 131.600 136.575 132.300 138.675 ;
    END
  END ext_trim[16]
  PIN ext_trim[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.680 0.000 62.380 2.100 ;
    END
  END ext_trim[15]
  PIN ext_trim[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.440 136.575 42.140 138.675 ;
    END
  END ext_trim[14]
  PIN ext_trim[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.880 136.575 71.580 138.675 ;
    END
  END ext_trim[13]
  PIN ext_trim[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.990 2.160 91.490 ;
    END
  END ext_trim[12]
  PIN ext_trim[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.320 0.000 32.020 2.100 ;
    END
  END ext_trim[11]
  PIN ext_trim[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.480 136.575 122.180 138.675 ;
    END
  END ext_trim[10]
  PIN ext_trim[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 60.760 136.575 61.460 138.675 ;
    END
  END ext_trim[9]
  PIN ext_trim[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.950 2.160 106.450 ;
    END
  END ext_trim[8]
  PIN ext_trim[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.150 2.160 31.650 ;
    END
  END ext_trim[7]
  PIN ext_trim[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 111.360 136.575 112.060 138.675 ;
    END
  END ext_trim[6]
  PIN ext_trim[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 101.240 136.575 101.940 138.675 ;
    END
  END ext_trim[5]
  PIN ext_trim[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.120 136.575 91.820 138.675 ;
    END
  END ext_trim[4]
  PIN ext_trim[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 136.515 24.710 138.675 26.210 ;
    END
  END ext_trim[3]
  PIN ext_trim[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.000 136.575 81.700 138.675 ;
    END
  END ext_trim[2]
  PIN ext_trim[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 136.515 38.310 138.675 39.810 ;
    END
  END ext_trim[1]
  PIN ext_trim[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.560 136.575 52.260 138.675 ;
    END
  END ext_trim[0]
  PIN vdd
    PORT
      LAYER met4 ;
        RECT 17.520 2.160 19.120 7.280 ;
    END
  END vdd
  PIN vss
    PORT
      LAYER met4 ;
        RECT 94.320 2.000 95.920 4.560 ;
    END
  END vss
  OBS
      LAYER li1 ;
        RECT 2.000 1.915 136.320 135.365 ;
      LAYER met1 ;
        RECT 2.000 1.760 136.320 136.600 ;
      LAYER met2 ;
        RECT 2.090 136.295 10.800 136.695 ;
        RECT 12.060 136.295 20.920 136.695 ;
        RECT 22.180 136.295 31.040 136.695 ;
        RECT 32.300 136.295 41.160 136.695 ;
        RECT 42.420 136.295 51.280 136.695 ;
        RECT 52.540 136.295 60.480 136.695 ;
        RECT 61.740 136.295 70.600 136.695 ;
        RECT 71.860 136.295 80.720 136.695 ;
        RECT 81.980 136.295 90.840 136.695 ;
        RECT 92.100 136.295 100.960 136.695 ;
        RECT 102.220 136.295 111.080 136.695 ;
        RECT 112.340 136.295 121.200 136.695 ;
        RECT 122.460 136.295 131.320 136.695 ;
        RECT 132.580 136.295 132.940 136.695 ;
        RECT 2.090 2.380 132.940 136.295 ;
        RECT 2.860 1.760 10.800 2.380 ;
        RECT 12.060 1.760 20.920 2.380 ;
        RECT 22.180 1.760 31.040 2.380 ;
        RECT 32.300 1.760 41.160 2.380 ;
        RECT 42.420 1.760 51.280 2.380 ;
        RECT 52.540 1.760 61.400 2.380 ;
        RECT 62.660 1.760 71.520 2.380 ;
        RECT 72.780 1.760 81.640 2.380 ;
        RECT 82.900 1.760 91.760 2.380 ;
        RECT 93.020 1.760 101.880 2.380 ;
        RECT 103.140 1.760 112.000 2.380 ;
        RECT 113.260 1.760 122.120 2.380 ;
        RECT 123.380 1.760 132.240 2.380 ;
      LAYER met3 ;
        RECT 2.560 134.470 136.745 135.520 ;
        RECT 1.930 129.970 136.745 134.470 ;
        RECT 1.930 127.670 136.115 129.970 ;
        RECT 1.930 121.810 136.745 127.670 ;
        RECT 2.560 119.510 136.745 121.810 ;
        RECT 1.930 115.010 136.745 119.510 ;
        RECT 1.930 112.710 136.115 115.010 ;
        RECT 1.930 106.850 136.745 112.710 ;
        RECT 2.560 104.550 136.745 106.850 ;
        RECT 1.930 100.050 136.745 104.550 ;
        RECT 1.930 97.750 136.115 100.050 ;
        RECT 1.930 91.890 136.745 97.750 ;
        RECT 2.560 89.590 136.745 91.890 ;
        RECT 1.930 85.090 136.745 89.590 ;
        RECT 1.930 82.790 136.115 85.090 ;
        RECT 1.930 76.930 136.745 82.790 ;
        RECT 2.560 74.630 136.745 76.930 ;
        RECT 1.930 70.130 136.745 74.630 ;
        RECT 1.930 67.830 136.115 70.130 ;
        RECT 1.930 61.970 136.745 67.830 ;
        RECT 2.560 59.670 136.745 61.970 ;
        RECT 1.930 55.170 136.745 59.670 ;
        RECT 1.930 52.870 136.115 55.170 ;
        RECT 1.930 47.010 136.745 52.870 ;
        RECT 2.560 44.710 136.745 47.010 ;
        RECT 1.930 40.210 136.745 44.710 ;
        RECT 1.930 37.910 136.115 40.210 ;
        RECT 1.930 32.050 136.745 37.910 ;
        RECT 2.560 29.750 136.745 32.050 ;
        RECT 1.930 26.610 136.745 29.750 ;
        RECT 1.930 24.310 136.115 26.610 ;
        RECT 1.930 17.090 136.745 24.310 ;
        RECT 2.560 14.790 136.745 17.090 ;
        RECT 1.930 11.650 136.745 14.790 ;
        RECT 1.930 9.350 136.115 11.650 ;
        RECT 1.930 1.760 136.745 9.350 ;
      LAYER met4 ;
        RECT 17.520 7.680 95.920 135.520 ;
        RECT 19.520 4.960 95.920 7.680 ;
        RECT 19.520 1.760 93.920 4.960 ;
      LAYER met5 ;
        RECT 2.000 17.850 136.320 96.040 ;
  END
END digital_pll
END LIBRARY

