magic
tech sky130A
magscale 1 2
timestamp 1586549923
<< checkpaint >>
rect -860 -908 32940 32716
<< locali >>
rect 23613 24455 23647 24761
rect 7237 19627 7271 19865
rect 8249 5551 8283 5721
rect 17357 2287 17391 2389
rect 17817 1675 17851 1845
rect 20209 1675 20243 1913
<< viali >>
rect 27661 30745 27695 30779
rect 19749 30609 19783 30643
rect 20025 30609 20059 30643
rect 27385 30609 27419 30643
rect 4753 30541 4787 30575
rect 5489 30541 5523 30575
rect 17541 30541 17575 30575
rect 28581 30541 28615 30575
rect 29133 30541 29167 30575
rect 5029 30473 5063 30507
rect 5305 30473 5339 30507
rect 17817 30473 17851 30507
rect 18093 30473 18127 30507
rect 28857 30473 28891 30507
rect 29317 30473 29351 30507
rect 18369 30405 18403 30439
rect 7513 30201 7547 30235
rect 28857 30201 28891 30235
rect 4017 30133 4051 30167
rect 4937 30133 4971 30167
rect 9261 30133 9295 30167
rect 3373 30065 3407 30099
rect 8985 30065 9019 30099
rect 12573 30065 12607 30099
rect 19197 30065 19231 30099
rect 20485 30065 20519 30099
rect 23061 30065 23095 30099
rect 24349 30065 24383 30099
rect 25821 30065 25855 30099
rect 28029 30065 28063 30099
rect 29317 30065 29351 30099
rect 3557 29997 3591 30031
rect 4661 29997 4695 30031
rect 6685 29997 6719 30031
rect 11009 29997 11043 30031
rect 12757 29997 12791 30031
rect 16161 29997 16195 30031
rect 16437 29997 16471 30031
rect 18185 29997 18219 30031
rect 23337 29997 23371 30031
rect 26005 29997 26039 30031
rect 28213 29997 28247 30031
rect 28673 29997 28707 30031
rect 29501 29997 29535 30031
rect 1073 29929 1107 29963
rect 13309 29929 13343 29963
rect 24533 29929 24567 29963
rect 1257 29861 1291 29895
rect 13217 29861 13251 29895
rect 20669 29861 20703 29895
rect 24165 29861 24199 29895
rect 3189 29657 3223 29691
rect 3373 29657 3407 29691
rect 4293 29657 4327 29691
rect 5029 29657 5063 29691
rect 7697 29657 7731 29691
rect 9537 29657 9571 29691
rect 16529 29657 16563 29691
rect 16897 29657 16931 29691
rect 19013 29657 19047 29691
rect 20485 29657 20519 29691
rect 23061 29657 23095 29691
rect 23337 29657 23371 29691
rect 23429 29657 23463 29691
rect 23613 29657 23647 29691
rect 26925 29657 26959 29691
rect 27845 29657 27879 29691
rect 4753 29589 4787 29623
rect 17173 29589 17207 29623
rect 981 29521 1015 29555
rect 3833 29521 3867 29555
rect 9445 29521 9479 29555
rect 10273 29521 10307 29555
rect 10549 29521 10583 29555
rect 11745 29521 11779 29555
rect 12021 29521 12055 29555
rect 12573 29521 12607 29555
rect 16437 29521 16471 29555
rect 17357 29521 17391 29555
rect 18461 29521 18495 29555
rect 24073 29521 24107 29555
rect 28581 29521 28615 29555
rect 4109 29453 4143 29487
rect 7237 29453 7271 29487
rect 7605 29453 7639 29487
rect 8157 29453 8191 29487
rect 9997 29453 10031 29487
rect 10733 29453 10767 29487
rect 12297 29453 12331 29487
rect 13033 29453 13067 29487
rect 15977 29453 16011 29487
rect 16713 29453 16747 29487
rect 17909 29453 17943 29487
rect 18185 29453 18219 29487
rect 18369 29453 18403 29487
rect 19565 29453 19599 29487
rect 20117 29453 20151 29487
rect 20577 29453 20611 29487
rect 20853 29453 20887 29487
rect 21405 29453 21439 29487
rect 24165 29453 24199 29487
rect 27017 29453 27051 29487
rect 1257 29385 1291 29419
rect 3005 29385 3039 29419
rect 4017 29385 4051 29419
rect 4937 29385 4971 29419
rect 7881 29385 7915 29419
rect 9077 29385 9111 29419
rect 12757 29385 12791 29419
rect 13309 29385 13343 29419
rect 15057 29385 15091 29419
rect 15793 29385 15827 29419
rect 16253 29385 16287 29419
rect 19841 29385 19875 29419
rect 21129 29385 21163 29419
rect 21589 29385 21623 29419
rect 24441 29385 24475 29419
rect 26189 29385 26223 29419
rect 27293 29385 27327 29419
rect 27569 29385 27603 29419
rect 27937 29385 27971 29419
rect 28213 29385 28247 29419
rect 28857 29385 28891 29419
rect 30605 29385 30639 29419
rect 889 29317 923 29351
rect 3465 29317 3499 29351
rect 3741 29317 3775 29351
rect 5213 29317 5247 29351
rect 9169 29317 9203 29351
rect 12941 29317 12975 29351
rect 15609 29317 15643 29351
rect 19473 29317 19507 29351
rect 23797 29317 23831 29351
rect 26281 29317 26315 29351
rect 26557 29317 26591 29351
rect 28397 29317 28431 29351
rect 1073 29113 1107 29147
rect 3925 29113 3959 29147
rect 16253 29113 16287 29147
rect 18093 29113 18127 29147
rect 24165 29113 24199 29147
rect 24625 29113 24659 29147
rect 29409 29113 29443 29147
rect 29961 29113 29995 29147
rect 4569 29045 4603 29079
rect 24349 29045 24383 29079
rect 3649 28977 3683 29011
rect 5029 28977 5063 29011
rect 5673 28977 5707 29011
rect 6869 28977 6903 29011
rect 8985 28977 9019 29011
rect 9169 28977 9203 29011
rect 10641 28977 10675 29011
rect 11837 28977 11871 29011
rect 13125 28977 13159 29011
rect 15057 28977 15091 29011
rect 15333 28977 15367 29011
rect 15425 28977 15459 29011
rect 16069 28977 16103 29011
rect 17081 28977 17115 29011
rect 17449 28977 17483 29011
rect 18921 28977 18955 29011
rect 20209 28977 20243 29011
rect 23521 28977 23555 29011
rect 26925 28977 26959 29011
rect 29777 28977 29811 29011
rect 4937 28909 4971 28943
rect 5581 28909 5615 28943
rect 12021 28909 12055 28943
rect 13309 28909 13343 28943
rect 14597 28909 14631 28943
rect 15701 28909 15735 28943
rect 17725 28909 17759 28943
rect 20393 28909 20427 28943
rect 23797 28909 23831 28943
rect 27201 28909 27235 28943
rect 28949 28909 28983 28943
rect 5305 28841 5339 28875
rect 8157 28841 8191 28875
rect 16989 28841 17023 28875
rect 1901 28773 1935 28807
rect 2085 28773 2119 28807
rect 3465 28773 3499 28807
rect 4017 28773 4051 28807
rect 4293 28773 4327 28807
rect 6225 28773 6259 28807
rect 6961 28773 6995 28807
rect 9261 28773 9295 28807
rect 9629 28773 9663 28807
rect 10457 28773 10491 28807
rect 18277 28773 18311 28807
rect 19197 28773 19231 28807
rect 24993 28773 25027 28807
rect 29593 28773 29627 28807
rect 1625 28569 1659 28603
rect 4293 28569 4327 28603
rect 5305 28569 5339 28603
rect 5673 28569 5707 28603
rect 6409 28569 6443 28603
rect 6869 28569 6903 28603
rect 9721 28569 9755 28603
rect 12849 28569 12883 28603
rect 13677 28569 13711 28603
rect 14965 28569 14999 28603
rect 15425 28569 15459 28603
rect 16989 28569 17023 28603
rect 17725 28569 17759 28603
rect 23705 28569 23739 28603
rect 24533 28569 24567 28603
rect 27201 28569 27235 28603
rect 27569 28569 27603 28603
rect 28213 28569 28247 28603
rect 29961 28569 29995 28603
rect 2177 28501 2211 28535
rect 5489 28501 5523 28535
rect 7973 28501 8007 28535
rect 8433 28501 8467 28535
rect 9629 28501 9663 28535
rect 12021 28501 12055 28535
rect 13953 28501 13987 28535
rect 17173 28501 17207 28535
rect 17633 28501 17667 28535
rect 23981 28501 24015 28535
rect 27293 28501 27327 28535
rect 1533 28433 1567 28467
rect 3097 28433 3131 28467
rect 4937 28433 4971 28467
rect 8249 28433 8283 28467
rect 9353 28433 9387 28467
rect 13217 28433 13251 28467
rect 13769 28433 13803 28467
rect 14505 28433 14539 28467
rect 16161 28433 16195 28467
rect 17449 28433 17483 28467
rect 18369 28433 18403 28467
rect 20117 28433 20151 28467
rect 21865 28433 21899 28467
rect 25085 28433 25119 28467
rect 25913 28433 25947 28467
rect 28765 28433 28799 28467
rect 1901 28365 1935 28399
rect 2177 28365 2211 28399
rect 2821 28365 2855 28399
rect 3557 28365 3591 28399
rect 4477 28365 4511 28399
rect 4661 28365 4695 28399
rect 5029 28365 5063 28399
rect 6317 28365 6351 28399
rect 7053 28365 7087 28399
rect 7605 28365 7639 28399
rect 8433 28365 8467 28399
rect 9077 28365 9111 28399
rect 9905 28365 9939 28399
rect 10089 28365 10123 28399
rect 10457 28365 10491 28399
rect 13033 28365 13067 28399
rect 14781 28365 14815 28399
rect 15793 28365 15827 28399
rect 18093 28365 18127 28399
rect 21589 28365 21623 28399
rect 22417 28365 22451 28399
rect 22785 28365 22819 28399
rect 22969 28365 23003 28399
rect 24993 28365 25027 28399
rect 25821 28365 25855 28399
rect 28029 28365 28063 28399
rect 28673 28365 28707 28399
rect 29501 28365 29535 28399
rect 29593 28365 29627 28399
rect 6133 28297 6167 28331
rect 10273 28297 10307 28331
rect 11101 28297 11135 28331
rect 15609 28297 15643 28331
rect 16437 28297 16471 28331
rect 20393 28297 20427 28331
rect 22233 28297 22267 28331
rect 23245 28297 23279 28331
rect 23521 28297 23555 28331
rect 24809 28297 24843 28331
rect 1349 28229 1383 28263
rect 3465 28229 3499 28263
rect 3925 28229 3959 28263
rect 5857 28229 5891 28263
rect 7697 28229 7731 28263
rect 10549 28229 10583 28263
rect 11009 28229 11043 28263
rect 11837 28229 11871 28263
rect 14689 28229 14723 28263
rect 15241 28229 15275 28263
rect 16345 28229 16379 28263
rect 18001 28229 18035 28263
rect 20209 28229 20243 28263
rect 27017 28229 27051 28263
rect 28397 28229 28431 28263
rect 29777 28229 29811 28263
rect 2729 28025 2763 28059
rect 4293 28025 4327 28059
rect 4477 28025 4511 28059
rect 4753 28025 4787 28059
rect 8157 28025 8191 28059
rect 9261 28025 9295 28059
rect 10365 28025 10399 28059
rect 15885 28025 15919 28059
rect 18921 28025 18955 28059
rect 19197 28025 19231 28059
rect 23061 28025 23095 28059
rect 24993 28025 25027 28059
rect 28673 28025 28707 28059
rect 3925 27957 3959 27991
rect 15149 27957 15183 27991
rect 18185 27957 18219 27991
rect 20577 27957 20611 27991
rect 24625 27957 24659 27991
rect 27201 27957 27235 27991
rect 1901 27889 1935 27923
rect 2085 27889 2119 27923
rect 3373 27889 3407 27923
rect 3557 27889 3591 27923
rect 5673 27889 5707 27923
rect 9261 27889 9295 27923
rect 9445 27889 9479 27923
rect 10549 27889 10583 27923
rect 15333 27889 15367 27923
rect 16805 27889 16839 27923
rect 20209 27889 20243 27923
rect 22417 27889 22451 27923
rect 24349 27889 24383 27923
rect 27937 27889 27971 27923
rect 28029 27889 28063 27923
rect 29685 27889 29719 27923
rect 2453 27821 2487 27855
rect 4109 27821 4143 27855
rect 4845 27821 4879 27855
rect 5397 27821 5431 27855
rect 5857 27821 5891 27855
rect 10825 27821 10859 27855
rect 12573 27821 12607 27855
rect 22601 27821 22635 27855
rect 27109 27821 27143 27855
rect 30053 27821 30087 27855
rect 7513 27753 7547 27787
rect 7329 27685 7363 27719
rect 15425 27685 15459 27719
rect 16621 27685 16655 27719
rect 2177 27481 2211 27515
rect 3925 27481 3959 27515
rect 5397 27481 5431 27515
rect 6961 27481 6995 27515
rect 9445 27481 9479 27515
rect 10365 27481 10399 27515
rect 10825 27481 10859 27515
rect 11009 27481 11043 27515
rect 14781 27481 14815 27515
rect 15977 27481 16011 27515
rect 20945 27481 20979 27515
rect 25085 27481 25119 27515
rect 27201 27481 27235 27515
rect 27569 27481 27603 27515
rect 29961 27481 29995 27515
rect 2361 27413 2395 27447
rect 5029 27413 5063 27447
rect 5305 27413 5339 27447
rect 7053 27413 7087 27447
rect 7237 27413 7271 27447
rect 7605 27413 7639 27447
rect 14965 27413 14999 27447
rect 15517 27413 15551 27447
rect 16621 27413 16655 27447
rect 27477 27413 27511 27447
rect 1349 27345 1383 27379
rect 3189 27345 3223 27379
rect 4937 27345 4971 27379
rect 9353 27345 9387 27379
rect 10641 27345 10675 27379
rect 11377 27345 11411 27379
rect 12665 27345 12699 27379
rect 20485 27345 20519 27379
rect 22969 27345 23003 27379
rect 1165 27277 1199 27311
rect 2545 27277 2579 27311
rect 2913 27277 2947 27311
rect 3097 27277 3131 27311
rect 7881 27277 7915 27311
rect 7973 27277 8007 27311
rect 8709 27277 8743 27311
rect 8893 27277 8927 27311
rect 9629 27277 9663 27311
rect 11561 27277 11595 27311
rect 12205 27277 12239 27311
rect 12573 27277 12607 27311
rect 15149 27277 15183 27311
rect 19933 27277 19967 27311
rect 1993 27209 2027 27243
rect 3649 27209 3683 27243
rect 6777 27209 6811 27243
rect 11193 27209 11227 27243
rect 11745 27209 11779 27243
rect 19749 27209 19783 27243
rect 20209 27209 20243 27243
rect 22325 27209 22359 27243
rect 22601 27209 22635 27243
rect 23245 27209 23279 27243
rect 24993 27209 25027 27243
rect 1073 27141 1107 27175
rect 1717 27141 1751 27175
rect 3557 27141 3591 27175
rect 15333 27141 15367 27175
rect 15701 27141 15735 27175
rect 16713 27141 16747 27175
rect 20669 27141 20703 27175
rect 22233 27141 22267 27175
rect 22785 27141 22819 27175
rect 27109 27141 27143 27175
rect 29685 27141 29719 27175
rect 2729 26937 2763 26971
rect 7513 26937 7547 26971
rect 8709 26937 8743 26971
rect 11837 26937 11871 26971
rect 23061 26937 23095 26971
rect 24441 26937 24475 26971
rect 9261 26869 9295 26903
rect 26097 26869 26131 26903
rect 3373 26801 3407 26835
rect 6593 26801 6627 26835
rect 9813 26801 9847 26835
rect 9997 26801 10031 26835
rect 10089 26801 10123 26835
rect 10641 26801 10675 26835
rect 14873 26801 14907 26835
rect 15149 26801 15183 26835
rect 16437 26801 16471 26835
rect 16529 26801 16563 26835
rect 21221 26801 21255 26835
rect 25821 26801 25855 26835
rect 28581 26801 28615 26835
rect 6961 26733 6995 26767
rect 10365 26733 10399 26767
rect 15333 26733 15367 26767
rect 21405 26733 21439 26767
rect 797 26665 831 26699
rect 6869 26665 6903 26699
rect 14965 26665 14999 26699
rect 981 26597 1015 26631
rect 3465 26597 3499 26631
rect 6758 26597 6792 26631
rect 7237 26597 7271 26631
rect 14689 26597 14723 26631
rect 16713 26597 16747 26631
rect 28765 26597 28799 26631
rect 5673 26393 5707 26427
rect 6409 26393 6443 26427
rect 7329 26393 7363 26427
rect 8157 26393 8191 26427
rect 8709 26393 8743 26427
rect 10273 26393 10307 26427
rect 12481 26393 12515 26427
rect 14137 26393 14171 26427
rect 16437 26393 16471 26427
rect 16621 26393 16655 26427
rect 16805 26393 16839 26427
rect 21405 26393 21439 26427
rect 21773 26393 21807 26427
rect 24625 26393 24659 26427
rect 24993 26393 25027 26427
rect 26097 26393 26131 26427
rect 28581 26393 28615 26427
rect 28765 26393 28799 26427
rect 6961 26325 6995 26359
rect 10181 26325 10215 26359
rect 20669 26325 20703 26359
rect 2729 26257 2763 26291
rect 7145 26257 7179 26291
rect 8525 26257 8559 26291
rect 9997 26257 10031 26291
rect 13953 26257 13987 26291
rect 14321 26257 14355 26291
rect 26925 26257 26959 26291
rect 27569 26257 27603 26291
rect 705 26189 739 26223
rect 4293 26189 4327 26223
rect 5949 26189 5983 26223
rect 6133 26189 6167 26223
rect 6225 26189 6259 26223
rect 6777 26189 6811 26223
rect 9261 26189 9295 26223
rect 9353 26189 9387 26223
rect 9629 26189 9663 26223
rect 9813 26189 9847 26223
rect 11745 26189 11779 26223
rect 14873 26189 14907 26223
rect 15057 26189 15091 26223
rect 15425 26189 15459 26223
rect 15517 26189 15551 26223
rect 17725 26189 17759 26223
rect 18461 26189 18495 26223
rect 20761 26189 20795 26223
rect 24901 26189 24935 26223
rect 27201 26189 27235 26223
rect 27661 26189 27695 26223
rect 29409 26189 29443 26223
rect 981 26121 1015 26155
rect 4845 26121 4879 26155
rect 12021 26121 12055 26155
rect 12297 26121 12331 26155
rect 18001 26121 18035 26155
rect 21037 26121 21071 26155
rect 21497 26121 21531 26155
rect 24717 26121 24751 26155
rect 25545 26121 25579 26155
rect 27017 26121 27051 26155
rect 27845 26121 27879 26155
rect 29685 26121 29719 26155
rect 29961 26121 29995 26155
rect 3373 26053 3407 26087
rect 3557 26053 3591 26087
rect 4569 26053 4603 26087
rect 4937 26053 4971 26087
rect 8249 26053 8283 26087
rect 14689 26053 14723 26087
rect 15793 26053 15827 26087
rect 18277 26053 18311 26087
rect 25453 26053 25487 26087
rect 25913 26053 25947 26087
rect 30145 26053 30179 26087
rect 1809 25849 1843 25883
rect 8709 25849 8743 25883
rect 9537 25849 9571 25883
rect 14689 25849 14723 25883
rect 15149 25849 15183 25883
rect 15333 25849 15367 25883
rect 23797 25849 23831 25883
rect 6041 25781 6075 25815
rect 6685 25781 6719 25815
rect 16161 25781 16195 25815
rect 18369 25781 18403 25815
rect 27293 25781 27327 25815
rect 4017 25713 4051 25747
rect 4385 25713 4419 25747
rect 5765 25713 5799 25747
rect 9261 25713 9295 25747
rect 14965 25713 14999 25747
rect 17817 25713 17851 25747
rect 18277 25713 18311 25747
rect 20209 25713 20243 25747
rect 21589 25713 21623 25747
rect 24533 25713 24567 25747
rect 26741 25713 26775 25747
rect 26925 25713 26959 25747
rect 28121 25713 28155 25747
rect 889 25645 923 25679
rect 3465 25645 3499 25679
rect 3925 25645 3959 25679
rect 4293 25645 4327 25679
rect 6869 25645 6903 25679
rect 16529 25645 16563 25679
rect 17725 25645 17759 25679
rect 20393 25645 20427 25679
rect 21865 25645 21899 25679
rect 23613 25645 23647 25679
rect 28397 25645 28431 25679
rect 28673 25645 28707 25679
rect 16621 25577 16655 25611
rect 17449 25577 17483 25611
rect 797 25509 831 25543
rect 9629 25509 9663 25543
rect 16299 25509 16333 25543
rect 16437 25509 16471 25543
rect 17541 25509 17575 25543
rect 24625 25509 24659 25543
rect 3465 25305 3499 25339
rect 4937 25305 4971 25339
rect 5673 25305 5707 25339
rect 12481 25305 12515 25339
rect 12849 25305 12883 25339
rect 16253 25305 16287 25339
rect 20209 25305 20243 25339
rect 21313 25305 21347 25339
rect 22233 25305 22267 25339
rect 22509 25305 22543 25339
rect 22693 25305 22727 25339
rect 23337 25305 23371 25339
rect 23981 25305 24015 25339
rect 24993 25305 25027 25339
rect 26465 25305 26499 25339
rect 26833 25305 26867 25339
rect 27201 25305 27235 25339
rect 1625 25237 1659 25271
rect 2085 25237 2119 25271
rect 3281 25237 3315 25271
rect 13217 25237 13251 25271
rect 16345 25237 16379 25271
rect 16805 25237 16839 25271
rect 21037 25237 21071 25271
rect 23613 25237 23647 25271
rect 4385 25169 4419 25203
rect 11009 25169 11043 25203
rect 16621 25169 16655 25203
rect 20025 25169 20059 25203
rect 20485 25169 20519 25203
rect 21865 25169 21899 25203
rect 24441 25169 24475 25203
rect 28029 25169 28063 25203
rect 28581 25169 28615 25203
rect 1441 25101 1475 25135
rect 2177 25101 2211 25135
rect 2361 25101 2395 25135
rect 2637 25101 2671 25135
rect 2729 25101 2763 25135
rect 4109 25101 4143 25135
rect 6133 25101 6167 25135
rect 6685 25101 6719 25135
rect 10365 25101 10399 25135
rect 12481 25101 12515 25135
rect 17357 25101 17391 25135
rect 20301 25101 20335 25135
rect 20853 25101 20887 25135
rect 21405 25101 21439 25135
rect 21589 25101 21623 25135
rect 24349 25101 24383 25135
rect 24717 25101 24751 25135
rect 24901 25101 24935 25135
rect 25821 25101 25855 25135
rect 26925 25101 26959 25135
rect 1257 25033 1291 25067
rect 3925 25033 3959 25067
rect 4753 25033 4787 25067
rect 6409 25033 6443 25067
rect 6869 25033 6903 25067
rect 10641 25033 10675 25067
rect 13493 25033 13527 25067
rect 17633 25033 17667 25067
rect 19381 25033 19415 25067
rect 22325 25033 22359 25067
rect 25177 25033 25211 25067
rect 26097 25033 26131 25067
rect 28213 25033 28247 25067
rect 28857 25033 28891 25067
rect 30605 25033 30639 25067
rect 3557 24965 3591 24999
rect 3833 24965 3867 24999
rect 4569 24965 4603 24999
rect 5857 24965 5891 24999
rect 11193 24965 11227 24999
rect 12665 24965 12699 24999
rect 13309 24965 13343 24999
rect 14965 24965 14999 24999
rect 15977 24965 16011 24999
rect 16989 24965 17023 24999
rect 17173 24965 17207 24999
rect 23153 24965 23187 24999
rect 26557 24965 26591 24999
rect 27845 24965 27879 24999
rect 28305 24965 28339 24999
rect 1809 24761 1843 24795
rect 3373 24761 3407 24795
rect 18185 24761 18219 24795
rect 23613 24761 23647 24795
rect 28765 24761 28799 24795
rect 17173 24693 17207 24727
rect 4477 24625 4511 24659
rect 4661 24625 4695 24659
rect 7605 24625 7639 24659
rect 9261 24625 9295 24659
rect 15609 24625 15643 24659
rect 15793 24625 15827 24659
rect 17909 24625 17943 24659
rect 20945 24625 20979 24659
rect 3649 24557 3683 24591
rect 4201 24557 4235 24591
rect 7053 24557 7087 24591
rect 7789 24557 7823 24591
rect 16161 24557 16195 24591
rect 17081 24557 17115 24591
rect 18001 24557 18035 24591
rect 21221 24557 21255 24591
rect 22969 24557 23003 24591
rect 26189 24693 26223 24727
rect 25913 24625 25947 24659
rect 27201 24625 27235 24659
rect 27569 24625 27603 24659
rect 28213 24625 28247 24659
rect 29593 24625 29627 24659
rect 28489 24557 28523 24591
rect 29777 24557 29811 24591
rect 28397 24489 28431 24523
rect 2177 24421 2211 24455
rect 9537 24421 9571 24455
rect 13309 24421 13343 24455
rect 18461 24421 18495 24455
rect 23613 24421 23647 24455
rect 23705 24421 23739 24455
rect 4201 24217 4235 24251
rect 9537 24217 9571 24251
rect 10457 24217 10491 24251
rect 12389 24217 12423 24251
rect 15701 24217 15735 24251
rect 16069 24217 16103 24251
rect 17357 24217 17391 24251
rect 17725 24217 17759 24251
rect 21313 24217 21347 24251
rect 21589 24217 21623 24251
rect 25913 24217 25947 24251
rect 26097 24217 26131 24251
rect 27385 24217 27419 24251
rect 28029 24217 28063 24251
rect 29777 24217 29811 24251
rect 29869 24217 29903 24251
rect 1993 24149 2027 24183
rect 2453 24149 2487 24183
rect 3741 24149 3775 24183
rect 17081 24149 17115 24183
rect 17633 24149 17667 24183
rect 21037 24149 21071 24183
rect 27293 24149 27327 24183
rect 29409 24149 29443 24183
rect 1809 24081 1843 24115
rect 3005 24081 3039 24115
rect 3925 24081 3959 24115
rect 6869 24081 6903 24115
rect 8985 24081 9019 24115
rect 9261 24081 9295 24115
rect 9997 24081 10031 24115
rect 10641 24081 10675 24115
rect 15885 24081 15919 24115
rect 2637 24013 2671 24047
rect 2729 24013 2763 24047
rect 3097 24013 3131 24047
rect 6501 24013 6535 24047
rect 6961 24013 6995 24047
rect 9813 24013 9847 24047
rect 11745 24013 11779 24047
rect 13217 24013 13251 24047
rect 19289 24013 19323 24047
rect 19841 24013 19875 24047
rect 28857 24013 28891 24047
rect 29225 24013 29259 24047
rect 29501 24013 29535 24047
rect 1625 23945 1659 23979
rect 6685 23945 6719 23979
rect 7237 23945 7271 23979
rect 12021 23945 12055 23979
rect 12941 23945 12975 23979
rect 13493 23945 13527 23979
rect 15241 23945 15275 23979
rect 19565 23945 19599 23979
rect 21221 23945 21255 23979
rect 27569 23945 27603 23979
rect 27845 23945 27879 23979
rect 4109 23877 4143 23911
rect 12573 23877 12607 23911
rect 13125 23877 13159 23911
rect 20025 23877 20059 23911
rect 2177 23673 2211 23707
rect 7697 23673 7731 23707
rect 7789 23673 7823 23707
rect 13217 23673 13251 23707
rect 24257 23673 24291 23707
rect 29593 23605 29627 23639
rect 1165 23537 1199 23571
rect 3373 23537 3407 23571
rect 6869 23537 6903 23571
rect 9077 23537 9111 23571
rect 11101 23537 11135 23571
rect 11561 23537 11595 23571
rect 18645 23537 18679 23571
rect 21589 23537 21623 23571
rect 22969 23537 23003 23571
rect 23153 23537 23187 23571
rect 27385 23537 27419 23571
rect 27569 23537 27603 23571
rect 28305 23537 28339 23571
rect 28489 23537 28523 23571
rect 29777 23537 29811 23571
rect 981 23469 1015 23503
rect 1441 23469 1475 23503
rect 7053 23469 7087 23503
rect 9353 23469 9387 23503
rect 10917 23469 10951 23503
rect 11469 23469 11503 23503
rect 18553 23469 18587 23503
rect 30145 23469 30179 23503
rect 11929 23401 11963 23435
rect 12297 23401 12331 23435
rect 26833 23401 26867 23435
rect 27201 23401 27235 23435
rect 797 23333 831 23367
rect 3649 23333 3683 23367
rect 6225 23333 6259 23367
rect 12389 23333 12423 23367
rect 18829 23333 18863 23367
rect 21681 23333 21715 23367
rect 23245 23333 23279 23367
rect 24073 23333 24107 23367
rect 3097 23129 3131 23163
rect 3833 23129 3867 23163
rect 5765 23129 5799 23163
rect 7697 23129 7731 23163
rect 10641 23129 10675 23163
rect 12481 23129 12515 23163
rect 14965 23129 14999 23163
rect 18001 23129 18035 23163
rect 18553 23129 18587 23163
rect 21313 23129 21347 23163
rect 23613 23129 23647 23163
rect 24257 23129 24291 23163
rect 25821 23129 25855 23163
rect 26925 23129 26959 23163
rect 27753 23129 27787 23163
rect 29961 23129 29995 23163
rect 30421 23129 30455 23163
rect 5949 23061 5983 23095
rect 6501 23061 6535 23095
rect 11285 23061 11319 23095
rect 27477 23061 27511 23095
rect 27661 23061 27695 23095
rect 29685 23061 29719 23095
rect 30145 23061 30179 23095
rect 981 22993 1015 23027
rect 2729 22993 2763 23027
rect 3373 22993 3407 23027
rect 4201 22993 4235 23027
rect 6317 22993 6351 23027
rect 7053 22993 7087 23027
rect 11101 22993 11135 23027
rect 11929 22993 11963 23027
rect 13125 22993 13159 23027
rect 18645 22993 18679 23027
rect 21497 22993 21531 23027
rect 21865 22993 21899 23027
rect 23245 22993 23279 23027
rect 23889 22993 23923 23027
rect 24441 22993 24475 23027
rect 24901 22993 24935 23027
rect 26189 22993 26223 23027
rect 27109 22993 27143 23027
rect 705 22925 739 22959
rect 3741 22925 3775 22959
rect 5581 22925 5615 22959
rect 6501 22925 6535 22959
rect 7329 22925 7363 22959
rect 12021 22925 12055 22959
rect 12665 22925 12699 22959
rect 12849 22925 12883 22959
rect 13217 22925 13251 22959
rect 14689 22925 14723 22959
rect 14781 22925 14815 22959
rect 21589 22925 21623 22959
rect 22141 22925 22175 22959
rect 22325 22925 22359 22959
rect 23337 22925 23371 22959
rect 24625 22925 24659 22959
rect 24993 22925 25027 22959
rect 26005 22925 26039 22959
rect 26557 22925 26591 22959
rect 3557 22857 3591 22891
rect 4385 22857 4419 22891
rect 9169 22857 9203 22891
rect 14321 22857 14355 22891
rect 18185 22857 18219 22891
rect 18921 22857 18955 22891
rect 20669 22857 20703 22891
rect 3281 22789 3315 22823
rect 9353 22789 9387 22823
rect 10825 22789 10859 22823
rect 11009 22789 11043 22823
rect 18277 22789 18311 22823
rect 22969 22789 23003 22823
rect 27201 22789 27235 22823
rect 30237 22789 30271 22823
rect 797 22585 831 22619
rect 1257 22585 1291 22619
rect 6133 22585 6167 22619
rect 6501 22585 6535 22619
rect 12297 22585 12331 22619
rect 18829 22585 18863 22619
rect 19105 22585 19139 22619
rect 24073 22585 24107 22619
rect 22049 22517 22083 22551
rect 3925 22449 3959 22483
rect 4109 22449 4143 22483
rect 4569 22449 4603 22483
rect 5029 22449 5063 22483
rect 7421 22449 7455 22483
rect 9997 22449 10031 22483
rect 13033 22449 13067 22483
rect 14689 22449 14723 22483
rect 16345 22449 16379 22483
rect 22509 22449 22543 22483
rect 22693 22449 22727 22483
rect 22969 22449 23003 22483
rect 23153 22449 23187 22483
rect 26373 22449 26407 22483
rect 26557 22449 26591 22483
rect 27017 22449 27051 22483
rect 27477 22449 27511 22483
rect 28581 22449 28615 22483
rect 28673 22449 28707 22483
rect 7605 22381 7639 22415
rect 10365 22381 10399 22415
rect 11745 22381 11779 22415
rect 13493 22381 13527 22415
rect 14873 22381 14907 22415
rect 23429 22381 23463 22415
rect 3373 22313 3407 22347
rect 3741 22313 3775 22347
rect 6869 22313 6903 22347
rect 25821 22313 25855 22347
rect 25913 22313 25947 22347
rect 889 22245 923 22279
rect 1349 22245 1383 22279
rect 6317 22245 6351 22279
rect 13033 22245 13067 22279
rect 16621 22245 16655 22279
rect 17449 22245 17483 22279
rect 18737 22245 18771 22279
rect 28857 22245 28891 22279
rect 2361 22041 2395 22075
rect 2913 22041 2947 22075
rect 3281 22041 3315 22075
rect 3649 22041 3683 22075
rect 5029 22041 5063 22075
rect 5949 22041 5983 22075
rect 8157 22041 8191 22075
rect 10457 22041 10491 22075
rect 16897 22041 16931 22075
rect 21773 22041 21807 22075
rect 22233 22041 22267 22075
rect 25361 22041 25395 22075
rect 28581 22041 28615 22075
rect 28765 22041 28799 22075
rect 28949 22041 28983 22075
rect 4937 21973 4971 22007
rect 6501 21973 6535 22007
rect 10089 21973 10123 22007
rect 13217 21973 13251 22007
rect 16621 21973 16655 22007
rect 17173 21973 17207 22007
rect 21957 21973 21991 22007
rect 25545 21973 25579 22007
rect 25821 21973 25855 22007
rect 27293 21973 27327 22007
rect 4293 21905 4327 21939
rect 5397 21905 5431 21939
rect 13401 21905 13435 21939
rect 15425 21905 15459 21939
rect 18093 21905 18127 21939
rect 22141 21905 22175 21939
rect 25729 21905 25763 21939
rect 26281 21905 26315 21939
rect 26925 21905 26959 21939
rect 2545 21837 2579 21871
rect 2637 21837 2671 21871
rect 3833 21837 3867 21871
rect 4017 21837 4051 21871
rect 4661 21837 4695 21871
rect 5765 21837 5799 21871
rect 6133 21837 6167 21871
rect 6685 21837 6719 21871
rect 7145 21837 7179 21871
rect 7421 21837 7455 21871
rect 7789 21837 7823 21871
rect 10549 21837 10583 21871
rect 17357 21837 17391 21871
rect 17541 21837 17575 21871
rect 17633 21837 17667 21871
rect 19105 21837 19139 21871
rect 19565 21837 19599 21871
rect 22417 21837 22451 21871
rect 26373 21837 26407 21871
rect 26557 21837 26591 21871
rect 10273 21769 10307 21803
rect 13125 21769 13159 21803
rect 13677 21769 13711 21803
rect 18185 21769 18219 21803
rect 18921 21769 18955 21803
rect 19841 21769 19875 21803
rect 3373 21701 3407 21735
rect 4569 21701 4603 21735
rect 5581 21701 5615 21735
rect 12665 21701 12699 21735
rect 12941 21701 12975 21735
rect 15517 21701 15551 21735
rect 16345 21701 16379 21735
rect 18737 21701 18771 21735
rect 19197 21701 19231 21735
rect 22693 21701 22727 21735
rect 26005 21701 26039 21735
rect 27109 21701 27143 21735
rect 3465 21497 3499 21531
rect 7513 21497 7547 21531
rect 13401 21497 13435 21531
rect 14781 21497 14815 21531
rect 16989 21497 17023 21531
rect 23429 21497 23463 21531
rect 3649 21429 3683 21463
rect 21773 21429 21807 21463
rect 1165 21361 1199 21395
rect 4385 21361 4419 21395
rect 4753 21361 4787 21395
rect 6593 21361 6627 21395
rect 11009 21361 11043 21395
rect 11193 21361 11227 21395
rect 11469 21361 11503 21395
rect 12849 21361 12883 21395
rect 17541 21361 17575 21395
rect 17725 21361 17759 21395
rect 17909 21361 17943 21395
rect 18369 21361 18403 21395
rect 22325 21361 22359 21395
rect 22417 21361 22451 21395
rect 22601 21361 22635 21395
rect 23245 21361 23279 21395
rect 24257 21361 24291 21395
rect 27017 21361 27051 21395
rect 27569 21361 27603 21395
rect 27753 21361 27787 21395
rect 28489 21361 28523 21395
rect 28673 21361 28707 21395
rect 981 21293 1015 21327
rect 1441 21293 1475 21327
rect 3741 21293 3775 21327
rect 4477 21293 4511 21327
rect 4661 21293 4695 21327
rect 5765 21293 5799 21327
rect 6317 21293 6351 21327
rect 6777 21293 6811 21327
rect 10549 21293 10583 21327
rect 11653 21293 11687 21327
rect 11929 21293 11963 21327
rect 13033 21293 13067 21327
rect 17081 21293 17115 21327
rect 18461 21293 18495 21327
rect 22877 21293 22911 21327
rect 24533 21293 24567 21327
rect 25821 21293 25855 21327
rect 27109 21225 27143 21259
rect 797 21157 831 21191
rect 6961 21157 6995 21191
rect 8801 21157 8835 21191
rect 29041 21157 29075 21191
rect 3373 20953 3407 20987
rect 3649 20953 3683 20987
rect 4017 20953 4051 20987
rect 4753 20953 4787 20987
rect 5213 20953 5247 20987
rect 5857 20953 5891 20987
rect 6593 20953 6627 20987
rect 10733 20953 10767 20987
rect 11101 20953 11135 20987
rect 12849 20953 12883 20987
rect 13033 20953 13067 20987
rect 16253 20953 16287 20987
rect 16437 20953 16471 20987
rect 16805 20953 16839 20987
rect 17173 20953 17207 20987
rect 21957 20953 21991 20987
rect 22141 20953 22175 20987
rect 22509 20953 22543 20987
rect 23245 20953 23279 20987
rect 24257 20953 24291 20987
rect 24533 20953 24567 20987
rect 26833 20953 26867 20987
rect 27109 20953 27143 20987
rect 27661 20953 27695 20987
rect 28029 20953 28063 20987
rect 5397 20885 5431 20919
rect 5673 20885 5707 20919
rect 9537 20885 9571 20919
rect 21497 20885 21531 20919
rect 22785 20885 22819 20919
rect 27845 20885 27879 20919
rect 2729 20817 2763 20851
rect 3833 20817 3867 20851
rect 4201 20817 4235 20851
rect 6409 20817 6443 20851
rect 7237 20817 7271 20851
rect 8433 20817 8467 20851
rect 11745 20817 11779 20851
rect 12389 20817 12423 20851
rect 17633 20817 17667 20851
rect 20025 20817 20059 20851
rect 20669 20817 20703 20851
rect 21681 20817 21715 20851
rect 23889 20817 23923 20851
rect 27385 20817 27419 20851
rect 28581 20817 28615 20851
rect 705 20749 739 20783
rect 4293 20749 4327 20783
rect 4661 20749 4695 20783
rect 6225 20749 6259 20783
rect 7329 20749 7363 20783
rect 7697 20749 7731 20783
rect 7881 20749 7915 20783
rect 8709 20749 8743 20783
rect 9077 20749 9111 20783
rect 9537 20749 9571 20783
rect 10641 20749 10675 20783
rect 11837 20749 11871 20783
rect 12573 20749 12607 20783
rect 16989 20749 17023 20783
rect 17357 20749 17391 20783
rect 20393 20749 20427 20783
rect 21865 20749 21899 20783
rect 23429 20749 23463 20783
rect 23613 20749 23647 20783
rect 23981 20749 24015 20783
rect 24993 20749 25027 20783
rect 25637 20749 25671 20783
rect 27293 20749 27327 20783
rect 981 20681 1015 20715
rect 4477 20681 4511 20715
rect 11285 20681 11319 20715
rect 12297 20681 12331 20715
rect 19381 20681 19415 20715
rect 20209 20681 20243 20715
rect 20853 20681 20887 20715
rect 22325 20681 22359 20715
rect 25269 20681 25303 20715
rect 25821 20681 25855 20715
rect 28857 20681 28891 20715
rect 30605 20681 30639 20715
rect 6961 20613 6995 20647
rect 8525 20613 8559 20647
rect 10365 20613 10399 20647
rect 11009 20613 11043 20647
rect 11561 20613 11595 20647
rect 16529 20613 16563 20647
rect 21129 20613 21163 20647
rect 28121 20613 28155 20647
rect 28305 20613 28339 20647
rect 1257 20409 1291 20443
rect 2085 20409 2119 20443
rect 5949 20409 5983 20443
rect 8709 20409 8743 20443
rect 9537 20409 9571 20443
rect 17357 20409 17391 20443
rect 23061 20409 23095 20443
rect 1349 20341 1383 20375
rect 7789 20341 7823 20375
rect 14689 20341 14723 20375
rect 16805 20341 16839 20375
rect 17633 20341 17667 20375
rect 18093 20341 18127 20375
rect 20945 20341 20979 20375
rect 23153 20341 23187 20375
rect 3373 20273 3407 20307
rect 5857 20273 5891 20307
rect 7053 20273 7087 20307
rect 7200 20273 7234 20307
rect 9261 20273 9295 20307
rect 9445 20273 9479 20307
rect 11009 20273 11043 20307
rect 11653 20273 11687 20307
rect 16529 20273 16563 20307
rect 17081 20273 17115 20307
rect 17817 20273 17851 20307
rect 21589 20273 21623 20307
rect 21957 20273 21991 20307
rect 27385 20273 27419 20307
rect 27661 20273 27695 20307
rect 27845 20273 27879 20307
rect 28121 20273 28155 20307
rect 28374 20273 28408 20307
rect 7421 20205 7455 20239
rect 11101 20205 11135 20239
rect 11745 20205 11779 20239
rect 21497 20205 21531 20239
rect 22049 20205 22083 20239
rect 28673 20205 28707 20239
rect 981 20137 1015 20171
rect 7329 20137 7363 20171
rect 12021 20137 12055 20171
rect 14965 20137 14999 20171
rect 797 20069 831 20103
rect 3465 20069 3499 20103
rect 6777 20069 6811 20103
rect 7973 20069 8007 20103
rect 9905 20069 9939 20103
rect 12113 20069 12147 20103
rect 20301 20069 20335 20103
rect 1165 19865 1199 19899
rect 1257 19865 1291 19899
rect 3465 19865 3499 19899
rect 6501 19865 6535 19899
rect 7237 19865 7271 19899
rect 9261 19865 9295 19899
rect 9813 19865 9847 19899
rect 10917 19865 10951 19899
rect 12205 19865 12239 19899
rect 14689 19865 14723 19899
rect 14873 19865 14907 19899
rect 16713 19865 16747 19899
rect 17909 19865 17943 19899
rect 19749 19865 19783 19899
rect 20301 19865 20335 19899
rect 23705 19865 23739 19899
rect 27201 19865 27235 19899
rect 27661 19865 27695 19899
rect 1901 19797 1935 19831
rect 2361 19797 2395 19831
rect 7145 19797 7179 19831
rect 1533 19729 1567 19763
rect 1717 19661 1751 19695
rect 2361 19661 2395 19695
rect 2637 19661 2671 19695
rect 2913 19661 2947 19695
rect 3189 19661 3223 19695
rect 6869 19661 6903 19695
rect 7421 19797 7455 19831
rect 8893 19797 8927 19831
rect 11193 19797 11227 19831
rect 18001 19797 18035 19831
rect 20025 19797 20059 19831
rect 21589 19797 21623 19831
rect 27753 19797 27787 19831
rect 28029 19797 28063 19831
rect 8433 19729 8467 19763
rect 10457 19729 10491 19763
rect 12573 19729 12607 19763
rect 20761 19729 20795 19763
rect 22693 19729 22727 19763
rect 23429 19729 23463 19763
rect 28857 19729 28891 19763
rect 29409 19729 29443 19763
rect 7973 19661 8007 19695
rect 8157 19661 8191 19695
rect 8525 19661 8559 19695
rect 9353 19661 9387 19695
rect 9997 19661 10031 19695
rect 10181 19661 10215 19695
rect 10549 19661 10583 19695
rect 11101 19661 11135 19695
rect 11745 19661 11779 19695
rect 11929 19661 11963 19695
rect 12021 19661 12055 19695
rect 13309 19661 13343 19695
rect 13769 19661 13803 19695
rect 20853 19661 20887 19695
rect 21221 19661 21255 19695
rect 21313 19661 21347 19695
rect 23153 19661 23187 19695
rect 28673 19661 28707 19695
rect 29225 19661 29259 19695
rect 3649 19593 3683 19627
rect 6777 19593 6811 19627
rect 7237 19593 7271 19627
rect 11377 19593 11411 19627
rect 13677 19593 13711 19627
rect 13953 19593 13987 19627
rect 21681 19593 21715 19627
rect 22969 19593 23003 19627
rect 28121 19593 28155 19627
rect 7789 19525 7823 19559
rect 8985 19525 9019 19559
rect 16621 19525 16655 19559
rect 19841 19525 19875 19559
rect 23797 19525 23831 19559
rect 27385 19525 27419 19559
rect 1993 19321 2027 19355
rect 7053 19321 7087 19355
rect 7605 19321 7639 19355
rect 9261 19321 9295 19355
rect 9629 19321 9663 19355
rect 10825 19321 10859 19355
rect 11929 19321 11963 19355
rect 12205 19321 12239 19355
rect 20301 19321 20335 19355
rect 20945 19321 20979 19355
rect 21405 19321 21439 19355
rect 23337 19321 23371 19355
rect 3649 19253 3683 19287
rect 6593 19253 6627 19287
rect 7697 19253 7731 19287
rect 9721 19253 9755 19287
rect 11837 19253 11871 19287
rect 16897 19253 16931 19287
rect 28949 19253 28983 19287
rect 3373 19185 3407 19219
rect 5029 19185 5063 19219
rect 6317 19185 6351 19219
rect 7881 19185 7915 19219
rect 10549 19185 10583 19219
rect 11561 19185 11595 19219
rect 12941 19185 12975 19219
rect 13125 19185 13159 19219
rect 14873 19185 14907 19219
rect 16161 19185 16195 19219
rect 16621 19185 16655 19219
rect 21957 19185 21991 19219
rect 23245 19185 23279 19219
rect 27937 19185 27971 19219
rect 29133 19185 29167 19219
rect 30513 19185 30547 19219
rect 5305 19117 5339 19151
rect 13493 19117 13527 19151
rect 15057 19117 15091 19151
rect 22141 19117 22175 19151
rect 27109 19117 27143 19151
rect 27661 19117 27695 19151
rect 28121 19117 28155 19151
rect 28581 19117 28615 19151
rect 29501 19117 29535 19151
rect 10365 18981 10399 19015
rect 21129 18981 21163 19015
rect 23889 18981 23923 19015
rect 3373 18777 3407 18811
rect 5305 18777 5339 18811
rect 6317 18777 6351 18811
rect 6501 18777 6535 18811
rect 10365 18777 10399 18811
rect 11285 18777 11319 18811
rect 11561 18777 11595 18811
rect 12297 18777 12331 18811
rect 12481 18777 12515 18811
rect 12849 18777 12883 18811
rect 13861 18777 13895 18811
rect 14965 18777 14999 18811
rect 15149 18777 15183 18811
rect 16161 18777 16195 18811
rect 16621 18777 16655 18811
rect 23245 18777 23279 18811
rect 23521 18777 23555 18811
rect 25913 18777 25947 18811
rect 26741 18777 26775 18811
rect 26925 18777 26959 18811
rect 27109 18777 27143 18811
rect 28857 18777 28891 18811
rect 29777 18777 29811 18811
rect 30421 18777 30455 18811
rect 3557 18709 3591 18743
rect 23153 18709 23187 18743
rect 27661 18709 27695 18743
rect 27937 18709 27971 18743
rect 29225 18709 29259 18743
rect 9261 18641 9295 18675
rect 9905 18641 9939 18675
rect 11929 18641 11963 18675
rect 12757 18641 12791 18675
rect 18001 18641 18035 18675
rect 24165 18641 24199 18675
rect 28581 18641 28615 18675
rect 29593 18641 29627 18675
rect 9077 18573 9111 18607
rect 9629 18573 9663 18607
rect 10457 18573 10491 18607
rect 11745 18573 11779 18607
rect 13033 18573 13067 18607
rect 13493 18573 13527 18607
rect 17541 18573 17575 18607
rect 18185 18573 18219 18607
rect 22049 18573 22083 18607
rect 23797 18573 23831 18607
rect 27477 18573 27511 18607
rect 28673 18573 28707 18607
rect 13401 18505 13435 18539
rect 13677 18505 13711 18539
rect 17357 18505 17391 18539
rect 17909 18505 17943 18539
rect 27569 18505 27603 18539
rect 5029 18437 5063 18471
rect 16437 18437 16471 18471
rect 17173 18437 17207 18471
rect 22141 18437 22175 18471
rect 23705 18437 23739 18471
rect 28121 18437 28155 18471
rect 28305 18437 28339 18471
rect 29409 18437 29443 18471
rect 6409 18165 6443 18199
rect 14597 18165 14631 18199
rect 26649 18165 26683 18199
rect 28305 18165 28339 18199
rect 4845 18097 4879 18131
rect 4992 18097 5026 18131
rect 6556 18097 6590 18131
rect 12849 18097 12883 18131
rect 12941 18097 12975 18131
rect 13125 18097 13159 18131
rect 14781 18097 14815 18131
rect 15149 18097 15183 18131
rect 16621 18097 16655 18131
rect 17081 18097 17115 18131
rect 18829 18097 18863 18131
rect 19013 18097 19047 18131
rect 26833 18097 26867 18131
rect 28029 18097 28063 18131
rect 5213 18029 5247 18063
rect 6777 18029 6811 18063
rect 13585 18029 13619 18063
rect 17173 18029 17207 18063
rect 20393 18029 20427 18063
rect 20761 18029 20795 18063
rect 22141 18029 22175 18063
rect 30053 18029 30087 18063
rect 5121 17961 5155 17995
rect 5305 17893 5339 17927
rect 6685 17893 6719 17927
rect 7053 17893 7087 17927
rect 17909 17893 17943 17927
rect 18829 17893 18863 17927
rect 19289 17893 19323 17927
rect 23797 17893 23831 17927
rect 24073 17893 24107 17927
rect 26925 17893 26959 17927
rect 3557 17689 3591 17723
rect 4293 17689 4327 17723
rect 5581 17689 5615 17723
rect 6501 17689 6535 17723
rect 6685 17689 6719 17723
rect 6777 17689 6811 17723
rect 6961 17689 6995 17723
rect 9077 17689 9111 17723
rect 12757 17689 12791 17723
rect 12849 17689 12883 17723
rect 13861 17689 13895 17723
rect 15425 17689 15459 17723
rect 17081 17689 17115 17723
rect 20301 17689 20335 17723
rect 21589 17689 21623 17723
rect 26373 17689 26407 17723
rect 28121 17689 28155 17723
rect 4661 17621 4695 17655
rect 9261 17621 9295 17655
rect 12573 17621 12607 17655
rect 13125 17621 13159 17655
rect 14321 17621 14355 17655
rect 14505 17621 14539 17655
rect 19933 17621 19967 17655
rect 20669 17621 20703 17655
rect 26741 17621 26775 17655
rect 28765 17621 28799 17655
rect 5397 17553 5431 17587
rect 8341 17553 8375 17587
rect 18185 17553 18219 17587
rect 23981 17553 24015 17587
rect 24349 17553 24383 17587
rect 25729 17553 25763 17587
rect 26557 17553 26591 17587
rect 28305 17553 28339 17587
rect 1809 17485 1843 17519
rect 3281 17485 3315 17519
rect 4753 17485 4787 17519
rect 5673 17485 5707 17519
rect 8433 17485 8467 17519
rect 13033 17485 13067 17519
rect 13309 17485 13343 17519
rect 14781 17485 14815 17519
rect 15241 17485 15275 17519
rect 17817 17485 17851 17519
rect 20853 17485 20887 17519
rect 20945 17485 20979 17519
rect 21681 17485 21715 17519
rect 27109 17485 27143 17519
rect 27569 17485 27603 17519
rect 1625 17417 1659 17451
rect 2545 17417 2579 17451
rect 3373 17417 3407 17451
rect 3649 17417 3683 17451
rect 5029 17417 5063 17451
rect 8249 17417 8283 17451
rect 8893 17417 8927 17451
rect 12389 17417 12423 17451
rect 13769 17417 13803 17451
rect 14597 17417 14631 17451
rect 16805 17417 16839 17451
rect 20117 17417 20151 17451
rect 21405 17417 21439 17451
rect 23797 17417 23831 17451
rect 26925 17417 26959 17451
rect 27845 17417 27879 17451
rect 1533 17349 1567 17383
rect 1901 17349 1935 17383
rect 2361 17349 2395 17383
rect 4385 17349 4419 17383
rect 7237 17349 7271 17383
rect 14137 17349 14171 17383
rect 14873 17349 14907 17383
rect 15609 17349 15643 17383
rect 16621 17349 16655 17383
rect 17541 17349 17575 17383
rect 17725 17349 17759 17383
rect 20393 17349 20427 17383
rect 21865 17349 21899 17383
rect 23429 17349 23463 17383
rect 23613 17349 23647 17383
rect 27201 17349 27235 17383
rect 28581 17349 28615 17383
rect 1257 17145 1291 17179
rect 12941 17145 12975 17179
rect 18185 17145 18219 17179
rect 20485 17145 20519 17179
rect 27017 17145 27051 17179
rect 4937 17077 4971 17111
rect 13033 17077 13067 17111
rect 14689 17077 14723 17111
rect 27845 17077 27879 17111
rect 1625 17009 1659 17043
rect 2085 17009 2119 17043
rect 4201 17009 4235 17043
rect 5213 17009 5247 17043
rect 5305 17009 5339 17043
rect 5489 17009 5523 17043
rect 6869 17009 6903 17043
rect 9077 17009 9111 17043
rect 9721 17009 9755 17043
rect 13217 17009 13251 17043
rect 15977 17009 16011 17043
rect 16437 17009 16471 17043
rect 18737 17009 18771 17043
rect 19105 17009 19139 17043
rect 20853 17009 20887 17043
rect 21221 17009 21255 17043
rect 22969 17009 23003 17043
rect 23337 17009 23371 17043
rect 27753 17009 27787 17043
rect 27937 17009 27971 17043
rect 1717 16941 1751 16975
rect 3373 16941 3407 16975
rect 3925 16941 3959 16975
rect 4385 16941 4419 16975
rect 5765 16941 5799 16975
rect 6777 16941 6811 16975
rect 7329 16941 7363 16975
rect 9813 16941 9847 16975
rect 16529 16941 16563 16975
rect 18553 16941 18587 16975
rect 19013 16941 19047 16975
rect 20669 16941 20703 16975
rect 21129 16941 21163 16975
rect 22877 16941 22911 16975
rect 23429 16941 23463 16975
rect 9261 16873 9295 16907
rect 17817 16873 17851 16907
rect 22417 16873 22451 16907
rect 1073 16805 1107 16839
rect 8525 16805 8559 16839
rect 14781 16805 14815 16839
rect 17541 16805 17575 16839
rect 19381 16805 19415 16839
rect 24073 16805 24107 16839
rect 28121 16805 28155 16839
rect 3925 16601 3959 16635
rect 4109 16601 4143 16635
rect 4293 16601 4327 16635
rect 4477 16601 4511 16635
rect 5213 16601 5247 16635
rect 5581 16601 5615 16635
rect 5765 16601 5799 16635
rect 7421 16601 7455 16635
rect 7605 16601 7639 16635
rect 15333 16601 15367 16635
rect 15977 16601 16011 16635
rect 16437 16601 16471 16635
rect 18277 16601 18311 16635
rect 20301 16601 20335 16635
rect 20485 16601 20519 16635
rect 20853 16601 20887 16635
rect 22509 16601 22543 16635
rect 23245 16601 23279 16635
rect 23705 16601 23739 16635
rect 24257 16601 24291 16635
rect 26925 16601 26959 16635
rect 27845 16601 27879 16635
rect 28213 16601 28247 16635
rect 3557 16533 3591 16567
rect 5489 16533 5523 16567
rect 12205 16533 12239 16567
rect 18093 16533 18127 16567
rect 20945 16533 20979 16567
rect 23797 16533 23831 16567
rect 27753 16533 27787 16567
rect 889 16465 923 16499
rect 2453 16465 2487 16499
rect 3373 16465 3407 16499
rect 8341 16465 8375 16499
rect 10457 16465 10491 16499
rect 14505 16465 14539 16499
rect 14965 16465 14999 16499
rect 16161 16465 16195 16499
rect 19289 16465 19323 16499
rect 22417 16465 22451 16499
rect 23429 16465 23463 16499
rect 24901 16465 24935 16499
rect 25913 16465 25947 16499
rect 1625 16397 1659 16431
rect 1809 16397 1843 16431
rect 1993 16397 2027 16431
rect 2545 16397 2579 16431
rect 3189 16397 3223 16431
rect 3741 16397 3775 16431
rect 7237 16397 7271 16431
rect 7789 16397 7823 16431
rect 8433 16397 8467 16431
rect 11745 16397 11779 16431
rect 14229 16397 14263 16431
rect 14781 16397 14815 16431
rect 17173 16397 17207 16431
rect 17449 16397 17483 16431
rect 17725 16397 17759 16431
rect 19381 16397 19415 16431
rect 19749 16397 19783 16431
rect 19841 16397 19875 16431
rect 24441 16397 24475 16431
rect 24625 16397 24659 16431
rect 24993 16397 25027 16431
rect 26281 16397 26315 16431
rect 26465 16397 26499 16431
rect 29961 16397 29995 16431
rect 30329 16397 30363 16431
rect 1165 16329 1199 16363
rect 2729 16329 2763 16363
rect 3005 16329 3039 16363
rect 6685 16329 6719 16363
rect 7329 16329 7363 16363
rect 8157 16329 8191 16363
rect 8709 16329 8743 16363
rect 12113 16329 12147 16363
rect 12389 16329 12423 16363
rect 18737 16329 18771 16363
rect 22693 16329 22727 16363
rect 23061 16329 23095 16363
rect 25729 16329 25763 16363
rect 981 16261 1015 16295
rect 6777 16261 6811 16295
rect 15149 16261 15183 16295
rect 18553 16261 18587 16295
rect 20577 16261 20611 16295
rect 26097 16261 26131 16295
rect 28029 16261 28063 16295
rect 29961 16261 29995 16295
rect 30145 16261 30179 16295
rect 1717 16057 1751 16091
rect 9261 16057 9295 16091
rect 18369 16057 18403 16091
rect 19289 16057 19323 16091
rect 24257 16057 24291 16091
rect 26741 16057 26775 16091
rect 1625 15989 1659 16023
rect 8433 15989 8467 16023
rect 9077 15989 9111 16023
rect 12481 15989 12515 16023
rect 16069 15989 16103 16023
rect 18461 15989 18495 16023
rect 23981 15989 24015 16023
rect 27569 15989 27603 16023
rect 1165 15921 1199 15955
rect 1993 15921 2027 15955
rect 3373 15921 3407 15955
rect 3557 15921 3591 15955
rect 5949 15921 5983 15955
rect 6317 15921 6351 15955
rect 6501 15921 6535 15955
rect 7605 15921 7639 15955
rect 7789 15921 7823 15955
rect 10733 15921 10767 15955
rect 11929 15921 11963 15955
rect 12113 15921 12147 15955
rect 15517 15921 15551 15955
rect 15701 15921 15735 15955
rect 19473 15921 19507 15955
rect 28213 15921 28247 15955
rect 28581 15921 28615 15955
rect 1441 15853 1475 15887
rect 2269 15853 2303 15887
rect 5857 15853 5891 15887
rect 7881 15853 7915 15887
rect 18093 15853 18127 15887
rect 19105 15853 19139 15887
rect 21865 15853 21899 15887
rect 22233 15853 22267 15887
rect 28121 15853 28155 15887
rect 28673 15853 28707 15887
rect 9353 15785 9387 15819
rect 3649 15717 3683 15751
rect 4753 15717 4787 15751
rect 5397 15717 5431 15751
rect 9537 15717 9571 15751
rect 11009 15717 11043 15751
rect 18921 15717 18955 15751
rect 24073 15717 24107 15751
rect 26557 15717 26591 15751
rect 1073 15513 1107 15547
rect 1993 15513 2027 15547
rect 2913 15513 2947 15547
rect 3465 15513 3499 15547
rect 4937 15513 4971 15547
rect 5765 15513 5799 15547
rect 6225 15513 6259 15547
rect 6961 15513 6995 15547
rect 7973 15513 8007 15547
rect 10733 15513 10767 15547
rect 11009 15513 11043 15547
rect 11469 15513 11503 15547
rect 12573 15513 12607 15547
rect 14873 15513 14907 15547
rect 15977 15513 16011 15547
rect 22141 15513 22175 15547
rect 22417 15513 22451 15547
rect 23981 15513 24015 15547
rect 24533 15513 24567 15547
rect 26557 15513 26591 15547
rect 28029 15513 28063 15547
rect 28857 15513 28891 15547
rect 3925 15445 3959 15479
rect 4109 15445 4143 15479
rect 5857 15445 5891 15479
rect 6869 15445 6903 15479
rect 12389 15445 12423 15479
rect 24165 15445 24199 15479
rect 26189 15445 26223 15479
rect 28305 15445 28339 15479
rect 4477 15377 4511 15411
rect 7237 15377 7271 15411
rect 8249 15377 8283 15411
rect 12757 15377 12791 15411
rect 18829 15377 18863 15411
rect 20577 15377 20611 15411
rect 23797 15377 23831 15411
rect 27569 15377 27603 15411
rect 28581 15377 28615 15411
rect 29225 15377 29259 15411
rect 2269 15309 2303 15343
rect 3373 15309 3407 15343
rect 4661 15309 4695 15343
rect 4845 15309 4879 15343
rect 8341 15309 8375 15343
rect 8709 15309 8743 15343
rect 8801 15309 8835 15343
rect 11745 15309 11779 15343
rect 11929 15309 11963 15343
rect 19197 15309 19231 15343
rect 24717 15309 24751 15343
rect 24901 15309 24935 15343
rect 25269 15309 25303 15343
rect 25453 15309 25487 15343
rect 26005 15309 26039 15343
rect 27109 15309 27143 15343
rect 27201 15309 27235 15343
rect 27477 15309 27511 15343
rect 27753 15309 27787 15343
rect 28673 15309 28707 15343
rect 29409 15309 29443 15343
rect 3097 15241 3131 15275
rect 3189 15241 3223 15275
rect 4201 15241 4235 15275
rect 7329 15241 7363 15275
rect 7513 15241 7547 15275
rect 11377 15241 11411 15275
rect 12297 15241 12331 15275
rect 14137 15241 14171 15275
rect 14505 15241 14539 15275
rect 14689 15241 14723 15275
rect 18461 15241 18495 15275
rect 21865 15241 21899 15275
rect 28121 15241 28155 15275
rect 5305 15173 5339 15207
rect 5489 15173 5523 15207
rect 15517 15173 15551 15207
rect 15701 15173 15735 15207
rect 18737 15173 18771 15207
rect 22233 15173 22267 15207
rect 26281 15173 26315 15207
rect 797 14969 831 15003
rect 3373 14969 3407 15003
rect 5581 14969 5615 15003
rect 7789 14969 7823 15003
rect 7973 14969 8007 15003
rect 8157 14969 8191 15003
rect 12113 14969 12147 15003
rect 19289 14969 19323 15003
rect 28581 14969 28615 15003
rect 6317 14901 6351 14935
rect 11377 14901 11411 14935
rect 14689 14901 14723 14935
rect 18829 14901 18863 14935
rect 27753 14901 27787 14935
rect 4477 14833 4511 14867
rect 4753 14833 4787 14867
rect 4845 14833 4879 14867
rect 6501 14833 6535 14867
rect 11561 14833 11595 14867
rect 23429 14833 23463 14867
rect 26373 14833 26407 14867
rect 27017 14833 27051 14867
rect 27109 14833 27143 14867
rect 27385 14833 27419 14867
rect 27477 14833 27511 14867
rect 4017 14765 4051 14799
rect 5121 14765 5155 14799
rect 5397 14765 5431 14799
rect 11929 14765 11963 14799
rect 23705 14765 23739 14799
rect 981 14629 1015 14663
rect 6593 14629 6627 14663
rect 14965 14629 14999 14663
rect 19197 14629 19231 14663
rect 24257 14629 24291 14663
rect 4017 14425 4051 14459
rect 4477 14425 4511 14459
rect 6501 14425 6535 14459
rect 6685 14425 6719 14459
rect 11101 14425 11135 14459
rect 11193 14425 11227 14459
rect 11469 14425 11503 14459
rect 12389 14425 12423 14459
rect 15333 14425 15367 14459
rect 16713 14425 16747 14459
rect 18737 14425 18771 14459
rect 19381 14425 19415 14459
rect 26097 14425 26131 14459
rect 26925 14425 26959 14459
rect 27569 14425 27603 14459
rect 3741 14357 3775 14391
rect 4937 14357 4971 14391
rect 5489 14357 5523 14391
rect 16529 14357 16563 14391
rect 2729 14289 2763 14323
rect 3925 14289 3959 14323
rect 4293 14289 4327 14323
rect 12573 14289 12607 14323
rect 15793 14289 15827 14323
rect 16437 14289 16471 14323
rect 18093 14289 18127 14323
rect 18553 14289 18587 14323
rect 19565 14289 19599 14323
rect 26649 14289 26683 14323
rect 27293 14289 27327 14323
rect 705 14221 739 14255
rect 4569 14221 4603 14255
rect 5121 14221 5155 14255
rect 5397 14221 5431 14255
rect 7605 14221 7639 14255
rect 8341 14221 8375 14255
rect 11745 14221 11779 14255
rect 11929 14221 11963 14255
rect 14505 14221 14539 14255
rect 16069 14221 16103 14255
rect 17817 14221 17851 14255
rect 18369 14221 18403 14255
rect 19749 14221 19783 14255
rect 20117 14221 20151 14255
rect 20301 14221 20335 14255
rect 23245 14221 23279 14255
rect 26741 14221 26775 14255
rect 981 14153 1015 14187
rect 7881 14153 7915 14187
rect 8249 14153 8283 14187
rect 14321 14153 14355 14187
rect 15885 14153 15919 14187
rect 23061 14153 23095 14187
rect 23521 14153 23555 14187
rect 24073 14153 24107 14187
rect 25913 14153 25947 14187
rect 6317 14085 6351 14119
rect 12021 14085 12055 14119
rect 14229 14085 14263 14119
rect 14597 14085 14631 14119
rect 15057 14085 15091 14119
rect 15241 14085 15275 14119
rect 18921 14085 18955 14119
rect 23797 14085 23831 14119
rect 24257 14085 24291 14119
rect 26189 14085 26223 14119
rect 26373 14085 26407 14119
rect 797 13881 831 13915
rect 14689 13881 14723 13915
rect 19749 13881 19783 13915
rect 21681 13881 21715 13915
rect 24809 13881 24843 13915
rect 26465 13881 26499 13915
rect 26741 13881 26775 13915
rect 11837 13813 11871 13847
rect 15241 13813 15275 13847
rect 15609 13813 15643 13847
rect 19197 13813 19231 13847
rect 12849 13745 12883 13779
rect 13033 13745 13067 13779
rect 18645 13745 18679 13779
rect 18737 13745 18771 13779
rect 22049 13745 22083 13779
rect 22417 13745 22451 13779
rect 23429 13745 23463 13779
rect 25821 13745 25855 13779
rect 25913 13745 25947 13779
rect 3373 13677 3407 13711
rect 3649 13677 3683 13711
rect 5397 13677 5431 13711
rect 15333 13677 15367 13711
rect 17357 13677 17391 13711
rect 21865 13677 21899 13711
rect 22325 13677 22359 13711
rect 23705 13677 23739 13711
rect 28397 13677 28431 13711
rect 28765 13677 28799 13711
rect 30145 13677 30179 13711
rect 981 13541 1015 13575
rect 12021 13541 12055 13575
rect 13125 13541 13159 13575
rect 18461 13541 18495 13575
rect 19289 13541 19323 13575
rect 24625 13541 24659 13575
rect 26097 13541 26131 13575
rect 3649 13337 3683 13371
rect 13125 13337 13159 13371
rect 13401 13337 13435 13371
rect 14689 13337 14723 13371
rect 15425 13337 15459 13371
rect 16529 13337 16563 13371
rect 18461 13337 18495 13371
rect 18645 13337 18679 13371
rect 19105 13337 19139 13371
rect 20117 13337 20151 13371
rect 21681 13337 21715 13371
rect 22141 13337 22175 13371
rect 23521 13337 23555 13371
rect 24257 13337 24291 13371
rect 24809 13337 24843 13371
rect 25821 13337 25855 13371
rect 26189 13337 26223 13371
rect 28949 13337 28983 13371
rect 3925 13269 3959 13303
rect 13217 13269 13251 13303
rect 14965 13269 14999 13303
rect 18829 13269 18863 13303
rect 19289 13269 19323 13303
rect 21497 13269 21531 13303
rect 3465 13201 3499 13235
rect 11193 13201 11227 13235
rect 12481 13201 12515 13235
rect 14873 13201 14907 13235
rect 23153 13201 23187 13235
rect 12389 13133 12423 13167
rect 12757 13133 12791 13167
rect 12849 13133 12883 13167
rect 13861 13133 13895 13167
rect 14229 13133 14263 13167
rect 15609 13133 15643 13167
rect 15793 13133 15827 13167
rect 16161 13133 16195 13167
rect 16345 13133 16379 13167
rect 17541 13133 17575 13167
rect 18001 13133 18035 13167
rect 19749 13133 19783 13167
rect 19933 13133 19967 13167
rect 21957 13133 21991 13167
rect 22509 13133 22543 13167
rect 22785 13133 22819 13167
rect 22969 13133 23003 13167
rect 23705 13133 23739 13167
rect 24993 13133 25027 13167
rect 25177 13133 25211 13167
rect 25545 13133 25579 13167
rect 25729 13133 25763 13167
rect 3833 13065 3867 13099
rect 11377 13065 11411 13099
rect 11745 13065 11779 13099
rect 17357 13065 17391 13099
rect 18185 13065 18219 13099
rect 19841 13065 19875 13099
rect 29133 13065 29167 13099
rect 11469 12997 11503 13031
rect 13677 12997 13711 13031
rect 14045 12997 14079 13031
rect 14505 12997 14539 13031
rect 17173 12997 17207 13031
rect 17633 12997 17667 13031
rect 19473 12997 19507 13031
rect 20485 12997 20519 13031
rect 21773 12997 21807 13031
rect 23981 12997 24015 13031
rect 24441 12997 24475 13031
rect 26097 12997 26131 13031
rect 28581 12997 28615 13031
rect 28857 12997 28891 13031
rect 15885 12793 15919 12827
rect 26925 12793 26959 12827
rect 8065 12725 8099 12759
rect 11929 12725 11963 12759
rect 12113 12725 12147 12759
rect 12757 12725 12791 12759
rect 15609 12725 15643 12759
rect 18737 12725 18771 12759
rect 1165 12657 1199 12691
rect 3373 12657 3407 12691
rect 4661 12657 4695 12691
rect 12941 12657 12975 12691
rect 14597 12657 14631 12691
rect 14781 12657 14815 12691
rect 14873 12657 14907 12691
rect 15333 12657 15367 12691
rect 16897 12657 16931 12691
rect 17265 12657 17299 12691
rect 18921 12657 18955 12691
rect 21773 12657 21807 12691
rect 24349 12657 24383 12691
rect 24717 12657 24751 12691
rect 24901 12657 24935 12691
rect 27109 12657 27143 12691
rect 1441 12589 1475 12623
rect 3557 12589 3591 12623
rect 4845 12589 4879 12623
rect 5949 12589 5983 12623
rect 6317 12589 6351 12623
rect 9905 12589 9939 12623
rect 10181 12589 10215 12623
rect 13309 12589 13343 12623
rect 15517 12589 15551 12623
rect 16989 12589 17023 12623
rect 17357 12589 17391 12623
rect 24165 12589 24199 12623
rect 28397 12589 28431 12623
rect 28765 12589 28799 12623
rect 30145 12589 30179 12623
rect 8249 12453 8283 12487
rect 16345 12453 16379 12487
rect 19013 12453 19047 12487
rect 20669 12453 20703 12487
rect 21773 12453 21807 12487
rect 23613 12453 23647 12487
rect 23981 12453 24015 12487
rect 1717 12249 1751 12283
rect 3649 12249 3683 12283
rect 4661 12249 4695 12283
rect 6409 12249 6443 12283
rect 10825 12249 10859 12283
rect 12941 12249 12975 12283
rect 13125 12249 13159 12283
rect 13309 12249 13343 12283
rect 14781 12249 14815 12283
rect 15241 12249 15275 12283
rect 15609 12249 15643 12283
rect 16161 12249 16195 12283
rect 16621 12249 16655 12283
rect 17081 12249 17115 12283
rect 18461 12249 18495 12283
rect 19197 12249 19231 12283
rect 21957 12249 21991 12283
rect 23061 12249 23095 12283
rect 27569 12249 27603 12283
rect 27845 12249 27879 12283
rect 28857 12249 28891 12283
rect 3465 12181 3499 12215
rect 10641 12181 10675 12215
rect 12757 12181 12791 12215
rect 14597 12181 14631 12215
rect 18553 12181 18587 12215
rect 23153 12181 23187 12215
rect 29869 12181 29903 12215
rect 1257 12113 1291 12147
rect 1533 12113 1567 12147
rect 3005 12113 3039 12147
rect 5581 12113 5615 12147
rect 5765 12113 5799 12147
rect 8157 12113 8191 12147
rect 8525 12113 8559 12147
rect 9905 12113 9939 12147
rect 10457 12113 10491 12147
rect 15701 12113 15735 12147
rect 16897 12113 16931 12147
rect 19749 12113 19783 12147
rect 20577 12113 20611 12147
rect 25269 12113 25303 12147
rect 27017 12113 27051 12147
rect 28029 12113 28063 12147
rect 28213 12113 28247 12147
rect 2729 12045 2763 12079
rect 3741 12045 3775 12079
rect 5213 12045 5247 12079
rect 6593 12045 6627 12079
rect 6777 12045 6811 12079
rect 7145 12045 7179 12079
rect 7329 12045 7363 12079
rect 12389 12045 12423 12079
rect 15885 12045 15919 12079
rect 15977 12045 16011 12079
rect 18737 12045 18771 12079
rect 18921 12045 18955 12079
rect 19105 12045 19139 12079
rect 21129 12045 21163 12079
rect 21313 12045 21347 12079
rect 21681 12045 21715 12079
rect 21865 12045 21899 12079
rect 23521 12045 23555 12079
rect 23889 12045 23923 12079
rect 26465 12045 26499 12079
rect 27293 12045 27327 12079
rect 29041 12045 29075 12079
rect 29225 12045 29259 12079
rect 29593 12045 29627 12079
rect 29777 12045 29811 12079
rect 5397 11977 5431 12011
rect 16713 11977 16747 12011
rect 20393 11977 20427 12011
rect 20669 11977 20703 12011
rect 22233 11977 22267 12011
rect 26741 11977 26775 12011
rect 28305 11977 28339 12011
rect 1993 11909 2027 11943
rect 2545 11909 2579 11943
rect 4845 11909 4879 11943
rect 5949 11909 5983 11943
rect 7789 11909 7823 11943
rect 8065 11909 8099 11943
rect 12113 11909 12147 11943
rect 12297 11909 12331 11943
rect 14965 11909 14999 11943
rect 19565 11909 19599 11943
rect 20117 11909 20151 11943
rect 23337 11909 23371 11943
rect 27385 11909 27419 11943
rect 6041 11705 6075 11739
rect 6317 11705 6351 11739
rect 8157 11705 8191 11739
rect 10273 11705 10307 11739
rect 16345 11705 16379 11739
rect 16437 11705 16471 11739
rect 17725 11705 17759 11739
rect 18921 11705 18955 11739
rect 23061 11705 23095 11739
rect 23705 11705 23739 11739
rect 23889 11705 23923 11739
rect 24165 11705 24199 11739
rect 28673 11705 28707 11739
rect 8985 11637 9019 11671
rect 28857 11637 28891 11671
rect 29317 11637 29351 11671
rect 1257 11569 1291 11603
rect 9629 11569 9663 11603
rect 9997 11569 10031 11603
rect 12573 11569 12607 11603
rect 17633 11569 17667 11603
rect 21313 11569 21347 11603
rect 29961 11569 29995 11603
rect 30329 11569 30363 11603
rect 6777 11501 6811 11535
rect 9721 11501 9755 11535
rect 9905 11501 9939 11535
rect 12481 11501 12515 11535
rect 20945 11501 20979 11535
rect 23521 11501 23555 11535
rect 26373 11501 26407 11535
rect 26741 11501 26775 11535
rect 28121 11501 28155 11535
rect 28949 11501 28983 11535
rect 29777 11501 29811 11535
rect 30237 11501 30271 11535
rect 6593 11433 6627 11467
rect 20669 11433 20703 11467
rect 29133 11433 29167 11467
rect 1441 11365 1475 11399
rect 6225 11365 6259 11399
rect 12757 11365 12791 11399
rect 24349 11365 24383 11399
rect 1349 11161 1383 11195
rect 8985 11161 9019 11195
rect 9169 11161 9203 11195
rect 12205 11161 12239 11195
rect 12757 11161 12791 11195
rect 15425 11161 15459 11195
rect 15609 11161 15643 11195
rect 17541 11161 17575 11195
rect 19841 11161 19875 11195
rect 20393 11161 20427 11195
rect 21313 11161 21347 11195
rect 21497 11161 21531 11195
rect 25821 11161 25855 11195
rect 26741 11161 26775 11195
rect 29501 11161 29535 11195
rect 29869 11161 29903 11195
rect 30053 11161 30087 11195
rect 8709 11093 8743 11127
rect 12389 11093 12423 11127
rect 17725 11093 17759 11127
rect 18461 11093 18495 11127
rect 20853 11093 20887 11127
rect 21221 11093 21255 11127
rect 25913 11093 25947 11127
rect 26097 11093 26131 11127
rect 6501 11025 6535 11059
rect 8893 11025 8927 11059
rect 13217 11025 13251 11059
rect 18645 11025 18679 11059
rect 27385 11025 27419 11059
rect 2453 10957 2487 10991
rect 3189 10957 3223 10991
rect 6133 10957 6167 10991
rect 9445 10957 9479 10991
rect 9905 10957 9939 10991
rect 12021 10957 12055 10991
rect 13309 10957 13343 10991
rect 13677 10957 13711 10991
rect 13769 10957 13803 10991
rect 14689 10957 14723 10991
rect 14873 10957 14907 10991
rect 17817 10957 17851 10991
rect 17909 10957 17943 10991
rect 20301 10957 20335 10991
rect 26925 10957 26959 10991
rect 27109 10957 27143 10991
rect 27477 10957 27511 10991
rect 29685 10957 29719 10991
rect 2729 10889 2763 10923
rect 9813 10889 9847 10923
rect 15241 10889 15275 10923
rect 18369 10889 18403 10923
rect 20025 10889 20059 10923
rect 20117 10889 20151 10923
rect 26281 10889 26315 10923
rect 1441 10821 1475 10855
rect 3005 10821 3039 10855
rect 5673 10821 5707 10855
rect 5949 10821 5983 10855
rect 8249 10821 8283 10855
rect 10181 10821 10215 10855
rect 12481 10821 12515 10855
rect 14597 10821 14631 10855
rect 20945 10821 20979 10855
rect 25637 10821 25671 10855
rect 29317 10821 29351 10855
rect 12665 10617 12699 10651
rect 13125 10617 13159 10651
rect 19381 10617 19415 10651
rect 26557 10617 26591 10651
rect 26925 10617 26959 10651
rect 28765 10617 28799 10651
rect 6869 10549 6903 10583
rect 12941 10549 12975 10583
rect 13677 10549 13711 10583
rect 16253 10549 16287 10583
rect 17909 10549 17943 10583
rect 26649 10549 26683 10583
rect 2177 10481 2211 10515
rect 3833 10481 3867 10515
rect 7513 10481 7547 10515
rect 7881 10481 7915 10515
rect 12573 10481 12607 10515
rect 13585 10481 13619 10515
rect 14597 10481 14631 10515
rect 14781 10481 14815 10515
rect 16345 10481 16379 10515
rect 18737 10481 18771 10515
rect 19105 10481 19139 10515
rect 26097 10481 26131 10515
rect 3741 10413 3775 10447
rect 7605 10413 7639 10447
rect 7789 10413 7823 10447
rect 18553 10413 18587 10447
rect 19013 10413 19047 10447
rect 22969 10413 23003 10447
rect 27017 10413 27051 10447
rect 4017 10277 4051 10311
rect 6225 10277 6259 10311
rect 8985 10277 9019 10311
rect 14873 10277 14907 10311
rect 16069 10277 16103 10311
rect 16529 10277 16563 10311
rect 17449 10277 17483 10311
rect 18369 10277 18403 10311
rect 23153 10277 23187 10311
rect 25913 10277 25947 10311
rect 28673 10277 28707 10311
rect 1993 10073 2027 10107
rect 4477 10073 4511 10107
rect 4569 10073 4603 10107
rect 7053 10073 7087 10107
rect 7513 10073 7547 10107
rect 8709 10073 8743 10107
rect 13585 10073 13619 10107
rect 14137 10073 14171 10107
rect 14505 10073 14539 10107
rect 15241 10073 15275 10107
rect 16069 10073 16103 10107
rect 16253 10073 16287 10107
rect 16621 10073 16655 10107
rect 17633 10073 17667 10107
rect 18369 10073 18403 10107
rect 18921 10073 18955 10107
rect 22785 10073 22819 10107
rect 25637 10073 25671 10107
rect 28673 10073 28707 10107
rect 7329 10005 7363 10039
rect 16529 10005 16563 10039
rect 2085 9937 2119 9971
rect 4109 9937 4143 9971
rect 4201 9937 4235 9971
rect 7605 9937 7639 9971
rect 8801 9937 8835 9971
rect 13401 9937 13435 9971
rect 17081 9937 17115 9971
rect 19381 9937 19415 9971
rect 22325 9937 22359 9971
rect 26557 9937 26591 9971
rect 28397 9937 28431 9971
rect 8433 9869 8467 9903
rect 14321 9869 14355 9903
rect 14781 9869 14815 9903
rect 15425 9869 15459 9903
rect 16897 9869 16931 9903
rect 17357 9869 17391 9903
rect 17541 9869 17575 9903
rect 19013 9869 19047 9903
rect 23429 9869 23463 9903
rect 23613 9869 23647 9903
rect 23981 9869 24015 9903
rect 24165 9869 24199 9903
rect 25729 9869 25763 9903
rect 26189 9869 26223 9903
rect 28029 9869 28063 9903
rect 29225 9869 29259 9903
rect 29317 9869 29351 9903
rect 29593 9869 29627 9903
rect 29777 9869 29811 9903
rect 1809 9801 1843 9835
rect 2361 9801 2395 9835
rect 8341 9801 8375 9835
rect 9077 9801 9111 9835
rect 10825 9801 10859 9835
rect 14597 9801 14631 9835
rect 15149 9801 15183 9835
rect 18185 9801 18219 9835
rect 18737 9801 18771 9835
rect 22601 9801 22635 9835
rect 22969 9801 23003 9835
rect 25269 9801 25303 9835
rect 6869 9733 6903 9767
rect 18461 9733 18495 9767
rect 21129 9733 21163 9767
rect 25361 9733 25395 9767
rect 25821 9733 25855 9767
rect 28213 9733 28247 9767
rect 2085 9529 2119 9563
rect 8985 9529 9019 9563
rect 11837 9529 11871 9563
rect 14689 9529 14723 9563
rect 18645 9529 18679 9563
rect 18829 9529 18863 9563
rect 19105 9529 19139 9563
rect 24625 9529 24659 9563
rect 24809 9529 24843 9563
rect 25913 9529 25947 9563
rect 3373 9461 3407 9495
rect 5489 9461 5523 9495
rect 9353 9461 9387 9495
rect 15885 9461 15919 9495
rect 26097 9461 26131 9495
rect 28397 9461 28431 9495
rect 1165 9393 1199 9427
rect 1717 9393 1751 9427
rect 3833 9393 3867 9427
rect 4017 9393 4051 9427
rect 4201 9393 4235 9427
rect 5673 9393 5707 9427
rect 9997 9393 10031 9427
rect 10365 9393 10399 9427
rect 16069 9393 16103 9427
rect 18001 9393 18035 9427
rect 18369 9393 18403 9427
rect 19289 9393 19323 9427
rect 22509 9393 22543 9427
rect 22877 9393 22911 9427
rect 26649 9393 26683 9427
rect 26741 9393 26775 9427
rect 27017 9393 27051 9427
rect 27477 9393 27511 9427
rect 28857 9393 28891 9427
rect 29041 9393 29075 9427
rect 29225 9393 29259 9427
rect 981 9325 1015 9359
rect 1441 9325 1475 9359
rect 6041 9325 6075 9359
rect 9813 9325 9847 9359
rect 10273 9325 10307 9359
rect 18093 9325 18127 9359
rect 18461 9325 18495 9359
rect 27201 9325 27235 9359
rect 29501 9325 29535 9359
rect 29777 9325 29811 9359
rect 797 9189 831 9223
rect 6225 9189 6259 9223
rect 12021 9189 12055 9223
rect 16161 9189 16195 9223
rect 17449 9189 17483 9223
rect 3189 8985 3223 9019
rect 4477 8985 4511 9019
rect 5489 8985 5523 9019
rect 9537 8985 9571 9019
rect 15517 8985 15551 9019
rect 15977 8985 16011 9019
rect 16253 8985 16287 9019
rect 16989 8985 17023 9019
rect 19105 8985 19139 9019
rect 22785 8985 22819 9019
rect 22969 8985 23003 9019
rect 24717 8985 24751 9019
rect 26373 8985 26407 9019
rect 28305 8985 28339 9019
rect 28673 8985 28707 9019
rect 29501 8985 29535 9019
rect 30053 8985 30087 9019
rect 5213 8917 5247 8951
rect 9905 8917 9939 8951
rect 11193 8917 11227 8951
rect 18829 8917 18863 8951
rect 23153 8917 23187 8951
rect 23797 8917 23831 8951
rect 24349 8917 24383 8951
rect 26189 8917 26223 8951
rect 29041 8917 29075 8951
rect 29869 8917 29903 8951
rect 705 8849 739 8883
rect 2729 8849 2763 8883
rect 3373 8849 3407 8883
rect 3557 8849 3591 8883
rect 4201 8849 4235 8883
rect 5673 8849 5707 8883
rect 6501 8849 6535 8883
rect 7973 8849 8007 8883
rect 9353 8849 9387 8883
rect 10181 8849 10215 8883
rect 12665 8849 12699 8883
rect 16805 8849 16839 8883
rect 22601 8849 22635 8883
rect 25177 8849 25211 8883
rect 3649 8781 3683 8815
rect 6133 8781 6167 8815
rect 12205 8781 12239 8815
rect 12389 8781 12423 8815
rect 12757 8781 12791 8815
rect 14781 8781 14815 8815
rect 15241 8781 15275 8815
rect 16069 8781 16103 8815
rect 17541 8781 17575 8815
rect 18277 8781 18311 8815
rect 18553 8781 18587 8815
rect 19657 8781 19691 8815
rect 19749 8781 19783 8815
rect 20025 8781 20059 8815
rect 20209 8781 20243 8815
rect 24165 8781 24199 8815
rect 25085 8781 25119 8815
rect 25453 8781 25487 8815
rect 25637 8781 25671 8815
rect 27109 8781 27143 8815
rect 27201 8781 27235 8815
rect 27477 8781 27511 8815
rect 27661 8781 27695 8815
rect 28029 8781 28063 8815
rect 29317 8781 29351 8815
rect 981 8713 1015 8747
rect 2913 8713 2947 8747
rect 4109 8713 4143 8747
rect 11377 8713 11411 8747
rect 11745 8713 11779 8747
rect 14597 8713 14631 8747
rect 17357 8713 17391 8747
rect 17817 8713 17851 8747
rect 18185 8713 18219 8747
rect 18645 8713 18679 8747
rect 23981 8713 24015 8747
rect 26465 8713 26499 8747
rect 28121 8713 28155 8747
rect 29225 8713 29259 8747
rect 3097 8645 3131 8679
rect 5397 8645 5431 8679
rect 5949 8645 5983 8679
rect 9721 8645 9755 8679
rect 11469 8645 11503 8679
rect 14505 8645 14539 8679
rect 14873 8645 14907 8679
rect 17173 8645 17207 8679
rect 25729 8645 25763 8679
rect 25913 8645 25947 8679
rect 28765 8645 28799 8679
rect 889 8441 923 8475
rect 1257 8441 1291 8475
rect 3925 8441 3959 8475
rect 17449 8441 17483 8475
rect 26373 8441 26407 8475
rect 27109 8441 27143 8475
rect 28397 8441 28431 8475
rect 29409 8441 29443 8475
rect 30053 8441 30087 8475
rect 3741 8373 3775 8407
rect 5305 8373 5339 8407
rect 17541 8373 17575 8407
rect 19105 8373 19139 8407
rect 24717 8373 24751 8407
rect 27201 8373 27235 8407
rect 1901 8305 1935 8339
rect 2269 8305 2303 8339
rect 2361 8305 2395 8339
rect 3649 8305 3683 8339
rect 5489 8305 5523 8339
rect 7513 8305 7547 8339
rect 7881 8305 7915 8339
rect 7973 8305 8007 8339
rect 10825 8305 10859 8339
rect 11193 8305 11227 8339
rect 20945 8305 20979 8339
rect 21221 8305 21255 8339
rect 21773 8305 21807 8339
rect 22877 8305 22911 8339
rect 24441 8305 24475 8339
rect 26649 8305 26683 8339
rect 28673 8305 28707 8339
rect 29225 8305 29259 8339
rect 29961 8305 29995 8339
rect 5857 8237 5891 8271
rect 6869 8237 6903 8271
rect 7329 8237 7363 8271
rect 12573 8237 12607 8271
rect 21497 8237 21531 8271
rect 22785 8237 22819 8271
rect 28857 8237 28891 8271
rect 797 8169 831 8203
rect 1717 8169 1751 8203
rect 21681 8169 21715 8203
rect 26189 8169 26223 8203
rect 26925 8169 26959 8203
rect 6225 8101 6259 8135
rect 23061 8101 23095 8135
rect 25085 8101 25119 8135
rect 26557 8101 26591 8135
rect 1901 7897 1935 7931
rect 2361 7897 2395 7931
rect 3373 7897 3407 7931
rect 3649 7897 3683 7931
rect 5305 7897 5339 7931
rect 5765 7897 5799 7931
rect 6225 7897 6259 7931
rect 6409 7897 6443 7931
rect 6593 7897 6627 7931
rect 11193 7897 11227 7931
rect 14321 7897 14355 7931
rect 17357 7897 17391 7931
rect 17817 7897 17851 7931
rect 20853 7897 20887 7931
rect 21405 7897 21439 7931
rect 22417 7897 22451 7931
rect 24257 7897 24291 7931
rect 28305 7897 28339 7931
rect 29225 7897 29259 7931
rect 29961 7897 29995 7931
rect 30145 7897 30179 7931
rect 11377 7829 11411 7863
rect 18185 7829 18219 7863
rect 20945 7829 20979 7863
rect 22785 7829 22819 7863
rect 23521 7829 23555 7863
rect 23797 7829 23831 7863
rect 2177 7761 2211 7795
rect 7421 7761 7455 7795
rect 8801 7761 8835 7795
rect 10917 7761 10951 7795
rect 15609 7761 15643 7795
rect 23245 7761 23279 7795
rect 25085 7761 25119 7795
rect 889 7693 923 7727
rect 1165 7693 1199 7727
rect 7053 7693 7087 7727
rect 13677 7693 13711 7727
rect 15057 7693 15091 7727
rect 17081 7693 17115 7727
rect 17633 7693 17667 7727
rect 21221 7693 21255 7727
rect 22601 7693 22635 7727
rect 22969 7693 23003 7727
rect 24993 7693 25027 7727
rect 25361 7693 25395 7727
rect 25545 7693 25579 7727
rect 28581 7693 28615 7727
rect 29317 7693 29351 7727
rect 1073 7625 1107 7659
rect 1441 7625 1475 7659
rect 11009 7625 11043 7659
rect 13953 7625 13987 7659
rect 15333 7625 15367 7659
rect 17541 7625 17575 7659
rect 24073 7625 24107 7659
rect 24349 7625 24383 7659
rect 28857 7625 28891 7659
rect 1809 7557 1843 7591
rect 5489 7557 5523 7591
rect 6777 7557 6811 7591
rect 6961 7557 6995 7591
rect 14413 7557 14447 7591
rect 15793 7557 15827 7591
rect 16897 7557 16931 7591
rect 20577 7557 20611 7591
rect 28121 7557 28155 7591
rect 6961 7353 6995 7387
rect 7237 7353 7271 7387
rect 7513 7353 7547 7387
rect 23061 7353 23095 7387
rect 24349 7353 24383 7387
rect 24533 7353 24567 7387
rect 24717 7353 24751 7387
rect 24901 7353 24935 7387
rect 5857 7285 5891 7319
rect 7145 7285 7179 7319
rect 18737 7285 18771 7319
rect 23613 7285 23647 7319
rect 3557 7217 3591 7251
rect 5305 7217 5339 7251
rect 5489 7217 5523 7251
rect 12297 7217 12331 7251
rect 14873 7217 14907 7251
rect 15057 7217 15091 7251
rect 18001 7217 18035 7251
rect 18185 7217 18219 7251
rect 18277 7217 18311 7251
rect 23337 7217 23371 7251
rect 26741 7217 26775 7251
rect 28857 7217 28891 7251
rect 29225 7217 29259 7251
rect 29317 7217 29351 7251
rect 3833 7149 3867 7183
rect 26649 7149 26683 7183
rect 28673 7149 28707 7183
rect 7789 7013 7823 7047
rect 12297 7013 12331 7047
rect 15149 7013 15183 7047
rect 20301 7013 20335 7047
rect 20577 7013 20611 7047
rect 26925 7013 26959 7047
rect 28489 7013 28523 7047
rect 3557 6809 3591 6843
rect 3833 6809 3867 6843
rect 5305 6809 5339 6843
rect 5765 6809 5799 6843
rect 7329 6809 7363 6843
rect 7973 6809 8007 6843
rect 11377 6809 11411 6843
rect 12021 6809 12055 6843
rect 12389 6809 12423 6843
rect 12757 6809 12791 6843
rect 14597 6809 14631 6843
rect 15425 6809 15459 6843
rect 18185 6809 18219 6843
rect 18645 6809 18679 6843
rect 23337 6809 23371 6843
rect 27569 6809 27603 6843
rect 28305 6809 28339 6843
rect 7145 6741 7179 6775
rect 7513 6741 7547 6775
rect 11561 6741 11595 6775
rect 18001 6741 18035 6775
rect 19841 6741 19875 6775
rect 23613 6741 23647 6775
rect 26373 6741 26407 6775
rect 26833 6741 26867 6775
rect 27017 6741 27051 6775
rect 27845 6741 27879 6775
rect 8157 6673 8191 6707
rect 13309 6673 13343 6707
rect 13861 6673 13895 6707
rect 19565 6673 19599 6707
rect 20761 6673 20795 6707
rect 27385 6673 27419 6707
rect 29317 6673 29351 6707
rect 29501 6673 29535 6707
rect 3005 6605 3039 6639
rect 4477 6605 4511 6639
rect 8341 6605 8375 6639
rect 8709 6605 8743 6639
rect 8801 6605 8835 6639
rect 11929 6605 11963 6639
rect 13125 6605 13159 6639
rect 13677 6605 13711 6639
rect 15333 6605 15367 6639
rect 15793 6605 15827 6639
rect 19013 6605 19047 6639
rect 19289 6605 19323 6639
rect 20945 6605 20979 6639
rect 21267 6605 21301 6639
rect 21497 6605 21531 6639
rect 24257 6605 24291 6639
rect 24625 6605 24659 6639
rect 26649 6605 26683 6639
rect 29225 6605 29259 6639
rect 29593 6605 29627 6639
rect 29869 6605 29903 6639
rect 3281 6537 3315 6571
rect 4753 6537 4787 6571
rect 5029 6537 5063 6571
rect 5581 6537 5615 6571
rect 11745 6537 11779 6571
rect 12573 6537 12607 6571
rect 14781 6537 14815 6571
rect 15149 6537 15183 6571
rect 18921 6537 18955 6571
rect 20025 6537 20059 6571
rect 20301 6537 20335 6571
rect 28029 6537 28063 6571
rect 2913 6469 2947 6503
rect 3925 6469 3959 6503
rect 4293 6469 4327 6503
rect 14873 6469 14907 6503
rect 16069 6469 16103 6503
rect 18461 6469 18495 6503
rect 20209 6469 20243 6503
rect 23889 6469 23923 6503
rect 24165 6469 24199 6503
rect 28213 6469 28247 6503
rect 28857 6469 28891 6503
rect 889 6265 923 6299
rect 7789 6265 7823 6299
rect 11837 6265 11871 6299
rect 15241 6265 15275 6299
rect 24257 6265 24291 6299
rect 29225 6265 29259 6299
rect 1165 6197 1199 6231
rect 29133 6197 29167 6231
rect 1993 6129 2027 6163
rect 3649 6129 3683 6163
rect 6777 6129 6811 6163
rect 9445 6129 9479 6163
rect 13217 6129 13251 6163
rect 15793 6129 15827 6163
rect 18277 6129 18311 6163
rect 20209 6129 20243 6163
rect 20577 6129 20611 6163
rect 27385 6129 27419 6163
rect 27753 6129 27787 6163
rect 28397 6129 28431 6163
rect 797 6061 831 6095
rect 1901 6061 1935 6095
rect 2453 6061 2487 6095
rect 2545 6061 2579 6095
rect 3925 6061 3959 6095
rect 5673 6061 5707 6095
rect 6961 6061 6995 6095
rect 9077 6061 9111 6095
rect 10825 6061 10859 6095
rect 13493 6061 13527 6095
rect 16069 6061 16103 6095
rect 21957 6061 21991 6095
rect 28305 6061 28339 6095
rect 27753 5993 27787 6027
rect 12021 5925 12055 5959
rect 18553 5925 18587 5959
rect 28857 5925 28891 5959
rect 2913 5721 2947 5755
rect 3097 5721 3131 5755
rect 3925 5721 3959 5755
rect 7053 5721 7087 5755
rect 7513 5721 7547 5755
rect 8157 5721 8191 5755
rect 8249 5721 8283 5755
rect 13217 5721 13251 5755
rect 13769 5721 13803 5755
rect 14137 5721 14171 5755
rect 15793 5721 15827 5755
rect 15977 5721 16011 5755
rect 18277 5721 18311 5755
rect 19841 5721 19875 5755
rect 20117 5721 20151 5755
rect 23889 5721 23923 5755
rect 24257 5721 24291 5755
rect 24717 5721 24751 5755
rect 26465 5721 26499 5755
rect 27569 5721 27603 5755
rect 705 5585 739 5619
rect 2729 5585 2763 5619
rect 3557 5585 3591 5619
rect 4017 5585 4051 5619
rect 8433 5653 8467 5687
rect 8617 5653 8651 5687
rect 11469 5653 11503 5687
rect 20393 5653 20427 5687
rect 22141 5653 22175 5687
rect 28029 5653 28063 5687
rect 28213 5653 28247 5687
rect 9905 5585 9939 5619
rect 11193 5585 11227 5619
rect 13861 5585 13895 5619
rect 14505 5585 14539 5619
rect 20301 5585 20335 5619
rect 21773 5585 21807 5619
rect 23981 5585 24015 5619
rect 25913 5585 25947 5619
rect 27845 5585 27879 5619
rect 3373 5517 3407 5551
rect 4477 5517 4511 5551
rect 4661 5517 4695 5551
rect 4845 5517 4879 5551
rect 6869 5517 6903 5551
rect 7421 5517 7455 5551
rect 8249 5517 8283 5551
rect 8985 5517 9019 5551
rect 9261 5517 9295 5551
rect 10089 5517 10123 5551
rect 10457 5517 10491 5551
rect 10549 5517 10583 5551
rect 12205 5517 12239 5551
rect 12389 5517 12423 5551
rect 12757 5517 12791 5551
rect 12849 5517 12883 5551
rect 13953 5517 13987 5551
rect 14689 5517 14723 5551
rect 15609 5517 15643 5551
rect 18737 5517 18771 5551
rect 19289 5517 19323 5551
rect 21313 5517 21347 5551
rect 21497 5517 21531 5551
rect 21865 5517 21899 5551
rect 24073 5517 24107 5551
rect 25637 5517 25671 5551
rect 26189 5517 26223 5551
rect 26925 5517 26959 5551
rect 27661 5517 27695 5551
rect 28581 5517 28615 5551
rect 981 5449 1015 5483
rect 3741 5449 3775 5483
rect 7237 5449 7271 5483
rect 7881 5449 7915 5483
rect 8801 5449 8835 5483
rect 9445 5449 9479 5483
rect 11377 5449 11411 5483
rect 11745 5449 11779 5483
rect 19013 5449 19047 5483
rect 19565 5449 19599 5483
rect 26833 5449 26867 5483
rect 27201 5449 27235 5483
rect 28857 5449 28891 5483
rect 29317 5449 29351 5483
rect 6593 5381 6627 5415
rect 9169 5381 9203 5415
rect 13493 5381 13527 5415
rect 15241 5381 15275 5415
rect 15425 5381 15459 5415
rect 16253 5381 16287 5415
rect 18553 5381 18587 5415
rect 20669 5381 20703 5415
rect 20945 5381 20979 5415
rect 24809 5381 24843 5415
rect 29133 5381 29167 5415
rect 889 5177 923 5211
rect 1165 5177 1199 5211
rect 3741 5177 3775 5211
rect 9537 5177 9571 5211
rect 9721 5177 9755 5211
rect 20945 5177 20979 5211
rect 27661 5177 27695 5211
rect 30513 5177 30547 5211
rect 797 5109 831 5143
rect 4109 5109 4143 5143
rect 7881 5109 7915 5143
rect 16989 5109 17023 5143
rect 21221 5109 21255 5143
rect 21681 5109 21715 5143
rect 23429 5109 23463 5143
rect 1441 5041 1475 5075
rect 1901 5041 1935 5075
rect 2269 5041 2303 5075
rect 4661 5041 4695 5075
rect 7329 5041 7363 5075
rect 7513 5041 7547 5075
rect 8985 5041 9019 5075
rect 10917 5041 10951 5075
rect 15425 5041 15459 5075
rect 15609 5041 15643 5075
rect 15885 5041 15919 5075
rect 16161 5041 16195 5075
rect 16354 5041 16388 5075
rect 18369 5041 18403 5075
rect 18737 5041 18771 5075
rect 21405 5041 21439 5075
rect 24257 5041 24291 5075
rect 27109 5041 27143 5075
rect 28397 5041 28431 5075
rect 2361 4973 2395 5007
rect 4201 4973 4235 5007
rect 4569 4973 4603 5007
rect 9169 4973 9203 5007
rect 10549 4973 10583 5007
rect 12297 4973 12331 5007
rect 17909 4973 17943 5007
rect 18829 4973 18863 5007
rect 24441 4973 24475 5007
rect 27293 4973 27327 5007
rect 28765 4973 28799 5007
rect 3833 4905 3867 4939
rect 4845 4837 4879 4871
rect 9997 4837 10031 4871
rect 21037 4837 21071 4871
rect 1625 4633 1659 4667
rect 1901 4633 1935 4667
rect 2085 4633 2119 4667
rect 4753 4633 4787 4667
rect 4937 4633 4971 4667
rect 7513 4633 7547 4667
rect 7789 4633 7823 4667
rect 8801 4633 8835 4667
rect 9537 4633 9571 4667
rect 10733 4633 10767 4667
rect 10917 4633 10951 4667
rect 15333 4633 15367 4667
rect 15885 4633 15919 4667
rect 16437 4633 16471 4667
rect 16621 4633 16655 4667
rect 16897 4633 16931 4667
rect 17449 4633 17483 4667
rect 21773 4633 21807 4667
rect 24257 4633 24291 4667
rect 27109 4633 27143 4667
rect 28949 4633 28983 4667
rect 4661 4565 4695 4599
rect 9813 4565 9847 4599
rect 14597 4565 14631 4599
rect 14689 4565 14723 4599
rect 15425 4565 15459 4599
rect 16253 4565 16287 4599
rect 17633 4565 17667 4599
rect 18185 4565 18219 4599
rect 19197 4565 19231 4599
rect 21589 4565 21623 4599
rect 10641 4497 10675 4531
rect 13677 4497 13711 4531
rect 19013 4497 19047 4531
rect 21957 4497 21991 4531
rect 6317 4429 6351 4463
rect 8893 4429 8927 4463
rect 13769 4429 13803 4463
rect 15149 4429 15183 4463
rect 15701 4429 15735 4463
rect 18369 4429 18403 4463
rect 18553 4429 18587 4463
rect 18737 4429 18771 4463
rect 29133 4429 29167 4463
rect 6133 4361 6167 4395
rect 6777 4361 6811 4395
rect 9169 4361 9203 4395
rect 9721 4361 9755 4395
rect 14229 4361 14263 4395
rect 14965 4361 14999 4395
rect 15609 4361 15643 4395
rect 17173 4361 17207 4395
rect 28765 4361 28799 4395
rect 1533 4293 1567 4327
rect 5949 4293 5983 4327
rect 6409 4293 6443 4327
rect 7053 4293 7087 4327
rect 7421 4293 7455 4327
rect 11193 4293 11227 4327
rect 13493 4293 13527 4327
rect 14413 4293 14447 4327
rect 17817 4293 17851 4327
rect 21497 4293 21531 4327
rect 24441 4293 24475 4327
rect 27293 4293 27327 4327
rect 28673 4293 28707 4327
rect 1257 4089 1291 4123
rect 13861 4089 13895 4123
rect 15609 4089 15643 4123
rect 18737 4089 18771 4123
rect 24901 4089 24935 4123
rect 25177 4089 25211 4123
rect 28213 4089 28247 4123
rect 7513 4021 7547 4055
rect 12297 4021 12331 4055
rect 17265 4021 17299 4055
rect 18553 4021 18587 4055
rect 26373 4021 26407 4055
rect 3465 3953 3499 3987
rect 5581 3953 5615 3987
rect 5765 3953 5799 3987
rect 5949 3953 5983 3987
rect 6961 3953 6995 3987
rect 7145 3953 7179 3987
rect 10917 3953 10951 3987
rect 11653 3953 11687 3987
rect 12021 3953 12055 3987
rect 14597 3953 14631 3987
rect 15885 3953 15919 3987
rect 17909 3953 17943 3987
rect 18277 3953 18311 3987
rect 21681 3953 21715 3987
rect 22049 3953 22083 3987
rect 23705 3953 23739 3987
rect 24073 3953 24107 3987
rect 24257 3953 24291 3987
rect 25821 3953 25855 3987
rect 25913 3953 25947 3987
rect 28397 3953 28431 3987
rect 3373 3885 3407 3919
rect 11745 3885 11779 3919
rect 11929 3885 11963 3919
rect 14781 3885 14815 3919
rect 15425 3885 15459 3919
rect 17817 3885 17851 3919
rect 18369 3885 18403 3919
rect 21497 3885 21531 3919
rect 21957 3885 21991 3919
rect 23797 3885 23831 3919
rect 28765 3885 28799 3919
rect 5397 3817 5431 3851
rect 9445 3817 9479 3851
rect 15977 3817 16011 3851
rect 2361 3749 2395 3783
rect 3649 3749 3683 3783
rect 11285 3749 11319 3783
rect 18921 3749 18955 3783
rect 21313 3749 21347 3783
rect 23337 3749 23371 3783
rect 30513 3749 30547 3783
rect 1257 3545 1291 3579
rect 3649 3545 3683 3579
rect 4017 3545 4051 3579
rect 5397 3545 5431 3579
rect 5489 3545 5523 3579
rect 6409 3545 6443 3579
rect 6961 3545 6995 3579
rect 7145 3545 7179 3579
rect 7421 3545 7455 3579
rect 11285 3545 11319 3579
rect 15057 3545 15091 3579
rect 15885 3545 15919 3579
rect 16069 3545 16103 3579
rect 16805 3545 16839 3579
rect 18185 3545 18219 3579
rect 19841 3545 19875 3579
rect 20393 3545 20427 3579
rect 21037 3545 21071 3579
rect 21313 3545 21347 3579
rect 21681 3545 21715 3579
rect 23337 3545 23371 3579
rect 27661 3545 27695 3579
rect 27845 3545 27879 3579
rect 28857 3545 28891 3579
rect 5213 3477 5247 3511
rect 10733 3477 10767 3511
rect 13217 3477 13251 3511
rect 17081 3477 17115 3511
rect 18001 3477 18035 3511
rect 24441 3477 24475 3511
rect 24901 3477 24935 3511
rect 25269 3477 25303 3511
rect 30237 3477 30271 3511
rect 4201 3409 4235 3443
rect 4937 3409 4971 3443
rect 8893 3409 8927 3443
rect 10089 3409 10123 3443
rect 10917 3409 10951 3443
rect 14505 3409 14539 3443
rect 15241 3409 15275 3443
rect 18645 3409 18679 3443
rect 19197 3409 19231 3443
rect 19933 3409 19967 3443
rect 21497 3409 21531 3443
rect 23613 3409 23647 3443
rect 29041 3409 29075 3443
rect 29869 3409 29903 3443
rect 2729 3341 2763 3375
rect 2913 3341 2947 3375
rect 3097 3341 3131 3375
rect 4334 3341 4368 3375
rect 5949 3341 5983 3375
rect 6133 3341 6167 3375
rect 6225 3341 6259 3375
rect 9997 3341 10031 3375
rect 10365 3341 10399 3375
rect 10457 3341 10491 3375
rect 12205 3341 12239 3375
rect 12389 3341 12423 3375
rect 12757 3341 12791 3375
rect 12941 3341 12975 3375
rect 14413 3341 14447 3375
rect 14781 3341 14815 3375
rect 14965 3341 14999 3375
rect 16989 3341 17023 3375
rect 18759 3341 18793 3375
rect 19105 3341 19139 3375
rect 20117 3341 20151 3375
rect 20209 3341 20243 3375
rect 24625 3341 24659 3375
rect 25545 3341 25579 3375
rect 25637 3341 25671 3375
rect 26097 3341 26131 3375
rect 26557 3341 26591 3375
rect 29225 3341 29259 3375
rect 29593 3341 29627 3375
rect 29777 3341 29811 3375
rect 1993 3273 2027 3307
rect 2269 3273 2303 3307
rect 4753 3273 4787 3307
rect 9077 3273 9111 3307
rect 9353 3273 9387 3307
rect 11561 3273 11595 3307
rect 13493 3273 13527 3307
rect 13769 3273 13803 3307
rect 19381 3273 19415 3307
rect 20761 3273 20795 3307
rect 21865 3273 21899 3307
rect 28029 3273 28063 3307
rect 28213 3273 28247 3307
rect 2177 3205 2211 3239
rect 3373 3205 3407 3239
rect 3925 3205 3959 3239
rect 5673 3205 5707 3239
rect 6777 3205 6811 3239
rect 9261 3205 9295 3239
rect 11101 3205 11135 3239
rect 11837 3205 11871 3239
rect 13585 3205 13619 3239
rect 17357 3205 17391 3239
rect 17541 3205 17575 3239
rect 17725 3205 17759 3239
rect 23153 3205 23187 3239
rect 23429 3205 23463 3239
rect 23889 3205 23923 3239
rect 24809 3205 24843 3239
rect 28305 3205 28339 3239
rect 30053 3205 30087 3239
rect 1073 3001 1107 3035
rect 2361 3001 2395 3035
rect 3373 3001 3407 3035
rect 5213 3001 5247 3035
rect 8157 3001 8191 3035
rect 9445 3001 9479 3035
rect 11837 3001 11871 3035
rect 12205 3001 12239 3035
rect 13769 3001 13803 3035
rect 18093 3001 18127 3035
rect 18277 3001 18311 3035
rect 23521 3001 23555 3035
rect 26189 3001 26223 3035
rect 5765 2933 5799 2967
rect 7513 2933 7547 2967
rect 11745 2933 11779 2967
rect 12113 2933 12147 2967
rect 13125 2933 13159 2967
rect 15517 2933 15551 2967
rect 17081 2933 17115 2967
rect 17633 2933 17667 2967
rect 18645 2933 18679 2967
rect 21405 2933 21439 2967
rect 23153 2933 23187 2967
rect 26097 2933 26131 2967
rect 4109 2865 4143 2899
rect 4477 2865 4511 2899
rect 4569 2865 4603 2899
rect 13309 2865 13343 2899
rect 15701 2865 15735 2899
rect 16897 2865 16931 2899
rect 17173 2865 17207 2899
rect 18737 2865 18771 2899
rect 21129 2865 21163 2899
rect 24993 2865 25027 2899
rect 28029 2865 28063 2899
rect 5489 2797 5523 2831
rect 9721 2797 9755 2831
rect 9997 2797 10031 2831
rect 16069 2797 16103 2831
rect 26373 2797 26407 2831
rect 28397 2797 28431 2831
rect 29777 2797 29811 2831
rect 3925 2729 3959 2763
rect 17909 2729 17943 2763
rect 19289 2729 19323 2763
rect 1257 2661 1291 2695
rect 13401 2661 13435 2695
rect 18461 2661 18495 2695
rect 18921 2661 18955 2695
rect 19473 2661 19507 2695
rect 25821 2661 25855 2695
rect 3373 2457 3407 2491
rect 4385 2457 4419 2491
rect 5673 2457 5707 2491
rect 6133 2457 6167 2491
rect 6961 2457 6995 2491
rect 10733 2457 10767 2491
rect 12481 2457 12515 2491
rect 15701 2457 15735 2491
rect 15977 2457 16011 2491
rect 16621 2457 16655 2491
rect 21221 2457 21255 2491
rect 21497 2457 21531 2491
rect 25821 2457 25855 2491
rect 28673 2457 28707 2491
rect 3741 2389 3775 2423
rect 5489 2389 5523 2423
rect 10549 2389 10583 2423
rect 16805 2389 16839 2423
rect 17357 2389 17391 2423
rect 18461 2389 18495 2423
rect 21681 2389 21715 2423
rect 22969 2389 23003 2423
rect 28029 2389 28063 2423
rect 1257 2321 1291 2355
rect 3557 2321 3591 2355
rect 4569 2321 4603 2355
rect 5949 2321 5983 2355
rect 6685 2321 6719 2355
rect 9813 2321 9847 2355
rect 12665 2321 12699 2355
rect 13401 2321 13435 2355
rect 16897 2321 16931 2355
rect 18185 2321 18219 2355
rect 19013 2321 19047 2355
rect 21313 2321 21347 2355
rect 23797 2321 23831 2355
rect 25545 2321 25579 2355
rect 26833 2321 26867 2355
rect 981 2253 1015 2287
rect 3189 2253 3223 2287
rect 3833 2253 3867 2287
rect 6409 2253 6443 2287
rect 7145 2253 7179 2287
rect 8065 2253 8099 2287
rect 8433 2253 8467 2287
rect 10917 2253 10951 2287
rect 13125 2253 13159 2287
rect 17357 2253 17391 2287
rect 17449 2253 17483 2287
rect 17909 2253 17943 2287
rect 18645 2253 18679 2287
rect 23521 2253 23555 2287
rect 27017 2253 27051 2287
rect 27385 2253 27419 2287
rect 27569 2253 27603 2287
rect 28765 2253 28799 2287
rect 3005 2185 3039 2219
rect 4109 2185 4143 2219
rect 10273 2185 10307 2219
rect 15149 2185 15183 2219
rect 15609 2185 15643 2219
rect 18369 2185 18403 2219
rect 23153 2185 23187 2219
rect 26097 2185 26131 2219
rect 26373 2185 26407 2219
rect 28305 2185 28339 2219
rect 889 2117 923 2151
rect 7697 2117 7731 2151
rect 7973 2117 8007 2151
rect 12757 2117 12791 2151
rect 13033 2117 13067 2151
rect 17173 2117 17207 2151
rect 17541 2117 17575 2151
rect 20761 2117 20795 2151
rect 23337 2117 23371 2151
rect 26281 2117 26315 2151
rect 1257 1913 1291 1947
rect 8157 1913 8191 1947
rect 13217 1913 13251 1947
rect 16989 1913 17023 1947
rect 18369 1913 18403 1947
rect 19381 1913 19415 1947
rect 20209 1913 20243 1947
rect 26465 1913 26499 1947
rect 4201 1845 4235 1879
rect 5949 1845 5983 1879
rect 13309 1845 13343 1879
rect 13493 1845 13527 1879
rect 17817 1845 17851 1879
rect 18001 1845 18035 1879
rect 1165 1777 1199 1811
rect 6777 1777 6811 1811
rect 9721 1777 9755 1811
rect 3925 1709 3959 1743
rect 6961 1709 6995 1743
rect 9997 1709 10031 1743
rect 11745 1709 11779 1743
rect 18553 1777 18587 1811
rect 18737 1777 18771 1811
rect 19105 1777 19139 1811
rect 19013 1709 19047 1743
rect 17817 1641 17851 1675
rect 20301 1777 20335 1811
rect 23889 1777 23923 1811
rect 24257 1777 24291 1811
rect 24441 1777 24475 1811
rect 27845 1777 27879 1811
rect 20669 1709 20703 1743
rect 22049 1709 22083 1743
rect 23705 1709 23739 1743
rect 27477 1709 27511 1743
rect 20209 1641 20243 1675
rect 2177 1573 2211 1607
rect 12757 1573 12791 1607
rect 15149 1573 15183 1607
rect 16713 1573 16747 1607
rect 23521 1573 23555 1607
rect 26005 1573 26039 1607
rect 29593 1573 29627 1607
rect 1073 1369 1107 1403
rect 4109 1369 4143 1403
rect 4385 1369 4419 1403
rect 6777 1369 6811 1403
rect 9813 1369 9847 1403
rect 10089 1369 10123 1403
rect 10365 1369 10399 1403
rect 18185 1369 18219 1403
rect 18461 1369 18495 1403
rect 18737 1369 18771 1403
rect 18921 1369 18955 1403
rect 19473 1369 19507 1403
rect 20853 1369 20887 1403
rect 21129 1369 21163 1403
rect 22417 1369 22451 1403
rect 27477 1369 27511 1403
rect 27845 1369 27879 1403
rect 28029 1369 28063 1403
rect 4017 1301 4051 1335
rect 9997 1301 10031 1335
rect 18369 1301 18403 1335
rect 22601 1301 22635 1335
rect 23245 1301 23279 1335
rect 27753 1301 27787 1335
rect 4569 1233 4603 1267
rect 6961 1233 6995 1267
rect 18001 1233 18035 1267
rect 19657 1233 19691 1267
rect 20577 1233 20611 1267
rect 22785 1233 22819 1267
rect 23705 1233 23739 1267
rect 25453 1233 25487 1267
rect 3557 1165 3591 1199
rect 19841 1165 19875 1199
rect 20209 1165 20243 1199
rect 20301 1165 20335 1199
rect 20669 1165 20703 1199
rect 23429 1165 23463 1199
rect 3741 1097 3775 1131
rect 19105 1097 19139 1131
rect 2085 1029 2119 1063
rect 12573 1029 12607 1063
rect 15057 1029 15091 1063
rect 16621 1029 16655 1063
rect 23061 1029 23095 1063
rect 25821 1029 25855 1063
rect 19473 825 19507 859
rect 23705 825 23739 859
rect 23889 825 23923 859
rect 19289 757 19323 791
rect 23981 757 24015 791
rect 23429 485 23463 519
<< metal1 >>
rect 400 31434 31680 31456
rect 400 31382 18870 31434
rect 18922 31382 18934 31434
rect 18986 31382 18998 31434
rect 19050 31382 19062 31434
rect 19114 31382 19126 31434
rect 19178 31382 31680 31434
rect 400 31360 31680 31382
rect 400 30890 31680 30912
rect 400 30838 3510 30890
rect 3562 30838 3574 30890
rect 3626 30838 3638 30890
rect 3690 30838 3702 30890
rect 3754 30838 3766 30890
rect 3818 30838 31680 30890
rect 400 30816 31680 30838
rect 27462 30776 27468 30788
rect 27388 30748 27468 30776
rect 2622 30668 2628 30720
rect 2680 30708 2686 30720
rect 8602 30708 8608 30720
rect 2680 30680 8608 30708
rect 2680 30668 2686 30680
rect 8602 30668 8608 30680
rect 8660 30668 8666 30720
rect 1150 30600 1156 30652
rect 1208 30640 1214 30652
rect 13386 30640 13392 30652
rect 1208 30612 13392 30640
rect 1208 30600 1214 30612
rect 13386 30600 13392 30612
rect 13444 30600 13450 30652
rect 19274 30600 19280 30652
rect 19332 30640 19338 30652
rect 27388 30649 27416 30748
rect 27462 30736 27468 30748
rect 27520 30776 27526 30788
rect 27649 30779 27707 30785
rect 27649 30776 27661 30779
rect 27520 30748 27661 30776
rect 27520 30736 27526 30748
rect 27649 30745 27661 30748
rect 27695 30745 27707 30779
rect 27649 30739 27707 30745
rect 19737 30643 19795 30649
rect 19737 30640 19749 30643
rect 19332 30612 19749 30640
rect 19332 30600 19338 30612
rect 19737 30609 19749 30612
rect 19783 30640 19795 30643
rect 20013 30643 20071 30649
rect 20013 30640 20025 30643
rect 19783 30612 20025 30640
rect 19783 30609 19795 30612
rect 19737 30603 19795 30609
rect 20013 30609 20025 30612
rect 20059 30609 20071 30643
rect 20013 30603 20071 30609
rect 27373 30643 27431 30649
rect 27373 30609 27385 30643
rect 27419 30609 27431 30643
rect 27373 30603 27431 30609
rect 4002 30532 4008 30584
rect 4060 30572 4066 30584
rect 4741 30575 4799 30581
rect 4741 30572 4753 30575
rect 4060 30544 4753 30572
rect 4060 30532 4066 30544
rect 4741 30541 4753 30544
rect 4787 30572 4799 30575
rect 5477 30575 5535 30581
rect 5477 30572 5489 30575
rect 4787 30544 5489 30572
rect 4787 30541 4799 30544
rect 4741 30535 4799 30541
rect 5477 30541 5489 30544
rect 5523 30572 5535 30575
rect 9982 30572 9988 30584
rect 5523 30544 9988 30572
rect 5523 30541 5535 30544
rect 5477 30535 5535 30541
rect 9982 30532 9988 30544
rect 10040 30532 10046 30584
rect 17529 30575 17587 30581
rect 17529 30541 17541 30575
rect 17575 30572 17587 30575
rect 17575 30544 18400 30572
rect 17575 30541 17587 30544
rect 17529 30535 17587 30541
rect 5014 30504 5020 30516
rect 4975 30476 5020 30504
rect 5014 30464 5020 30476
rect 5072 30504 5078 30516
rect 5293 30507 5351 30513
rect 5293 30504 5305 30507
rect 5072 30476 5305 30504
rect 5072 30464 5078 30476
rect 5293 30473 5305 30476
rect 5339 30504 5351 30507
rect 5382 30504 5388 30516
rect 5339 30476 5388 30504
rect 5339 30473 5351 30476
rect 5293 30467 5351 30473
rect 5382 30464 5388 30476
rect 5440 30464 5446 30516
rect 9430 30464 9436 30516
rect 9488 30504 9494 30516
rect 9890 30504 9896 30516
rect 9488 30476 9896 30504
rect 9488 30464 9494 30476
rect 9890 30464 9896 30476
rect 9948 30464 9954 30516
rect 16882 30464 16888 30516
rect 16940 30504 16946 30516
rect 17805 30507 17863 30513
rect 17805 30504 17817 30507
rect 16940 30476 17817 30504
rect 16940 30464 16946 30476
rect 17805 30473 17817 30476
rect 17851 30504 17863 30507
rect 18081 30507 18139 30513
rect 18081 30504 18093 30507
rect 17851 30476 18093 30504
rect 17851 30473 17863 30476
rect 17805 30467 17863 30473
rect 18081 30473 18093 30476
rect 18127 30473 18139 30507
rect 18081 30467 18139 30473
rect 18372 30448 18400 30544
rect 26910 30532 26916 30584
rect 26968 30572 26974 30584
rect 28569 30575 28627 30581
rect 28569 30572 28581 30575
rect 26968 30544 28581 30572
rect 26968 30532 26974 30544
rect 28569 30541 28581 30544
rect 28615 30572 28627 30575
rect 29121 30575 29179 30581
rect 29121 30572 29133 30575
rect 28615 30544 29133 30572
rect 28615 30541 28627 30544
rect 28569 30535 28627 30541
rect 29121 30541 29133 30544
rect 29167 30541 29179 30575
rect 29121 30535 29179 30541
rect 28842 30504 28848 30516
rect 28755 30476 28848 30504
rect 28842 30464 28848 30476
rect 28900 30504 28906 30516
rect 29305 30507 29363 30513
rect 29305 30504 29317 30507
rect 28900 30476 29317 30504
rect 28900 30464 28906 30476
rect 29305 30473 29317 30476
rect 29351 30473 29363 30507
rect 29305 30467 29363 30473
rect 3910 30396 3916 30448
rect 3968 30436 3974 30448
rect 10166 30436 10172 30448
rect 3968 30408 10172 30436
rect 3968 30396 3974 30408
rect 10166 30396 10172 30408
rect 10224 30396 10230 30448
rect 18354 30436 18360 30448
rect 18315 30408 18360 30436
rect 18354 30396 18360 30408
rect 18412 30396 18418 30448
rect 400 30346 31680 30368
rect 400 30294 18870 30346
rect 18922 30294 18934 30346
rect 18986 30294 18998 30346
rect 19050 30294 19062 30346
rect 19114 30294 19126 30346
rect 19178 30294 31680 30346
rect 400 30272 31680 30294
rect 414 30192 420 30244
rect 472 30232 478 30244
rect 6486 30232 6492 30244
rect 472 30204 6492 30232
rect 472 30192 478 30204
rect 6486 30192 6492 30204
rect 6544 30192 6550 30244
rect 6670 30192 6676 30244
rect 6728 30232 6734 30244
rect 7501 30235 7559 30241
rect 7501 30232 7513 30235
rect 6728 30204 7513 30232
rect 6728 30192 6734 30204
rect 7501 30201 7513 30204
rect 7547 30232 7559 30235
rect 7682 30232 7688 30244
rect 7547 30204 7688 30232
rect 7547 30201 7559 30204
rect 7501 30195 7559 30201
rect 7682 30192 7688 30204
rect 7740 30192 7746 30244
rect 13662 30192 13668 30244
rect 13720 30232 13726 30244
rect 14858 30232 14864 30244
rect 13720 30204 14864 30232
rect 13720 30192 13726 30204
rect 14858 30192 14864 30204
rect 14916 30192 14922 30244
rect 14950 30192 14956 30244
rect 15008 30232 15014 30244
rect 18538 30232 18544 30244
rect 15008 30204 18544 30232
rect 15008 30192 15014 30204
rect 18538 30192 18544 30204
rect 18596 30192 18602 30244
rect 28842 30232 28848 30244
rect 28803 30204 28848 30232
rect 28842 30192 28848 30204
rect 28900 30192 28906 30244
rect 4002 30164 4008 30176
rect 3963 30136 4008 30164
rect 4002 30124 4008 30136
rect 4060 30124 4066 30176
rect 4462 30124 4468 30176
rect 4520 30164 4526 30176
rect 4925 30167 4983 30173
rect 4925 30164 4937 30167
rect 4520 30136 4937 30164
rect 4520 30124 4526 30136
rect 4925 30133 4937 30136
rect 4971 30133 4983 30167
rect 4925 30127 4983 30133
rect 5382 30124 5388 30176
rect 5440 30124 5446 30176
rect 9154 30124 9160 30176
rect 9212 30164 9218 30176
rect 9249 30167 9307 30173
rect 9249 30164 9261 30167
rect 9212 30136 9261 30164
rect 9212 30124 9218 30136
rect 9249 30133 9261 30136
rect 9295 30133 9307 30167
rect 9249 30127 9307 30133
rect 10258 30124 10264 30176
rect 10316 30124 10322 30176
rect 16882 30124 16888 30176
rect 16940 30124 16946 30176
rect 3361 30099 3419 30105
rect 3361 30065 3373 30099
rect 3407 30096 3419 30099
rect 4020 30096 4048 30124
rect 3407 30068 4048 30096
rect 3407 30065 3419 30068
rect 3361 30059 3419 30065
rect 6302 30056 6308 30108
rect 6360 30096 6366 30108
rect 8970 30096 8976 30108
rect 6360 30068 8976 30096
rect 6360 30056 6366 30068
rect 8970 30056 8976 30068
rect 9028 30056 9034 30108
rect 12558 30096 12564 30108
rect 12519 30068 12564 30096
rect 12558 30056 12564 30068
rect 12616 30056 12622 30108
rect 17710 30056 17716 30108
rect 17768 30096 17774 30108
rect 18998 30096 19004 30108
rect 17768 30068 19004 30096
rect 17768 30056 17774 30068
rect 18998 30056 19004 30068
rect 19056 30096 19062 30108
rect 19185 30099 19243 30105
rect 19185 30096 19197 30099
rect 19056 30068 19197 30096
rect 19056 30056 19062 30068
rect 19185 30065 19197 30068
rect 19231 30065 19243 30099
rect 20470 30096 20476 30108
rect 20431 30068 20476 30096
rect 19185 30059 19243 30065
rect 20470 30056 20476 30068
rect 20528 30056 20534 30108
rect 23046 30096 23052 30108
rect 23007 30068 23052 30096
rect 23046 30056 23052 30068
rect 23104 30056 23110 30108
rect 24337 30099 24395 30105
rect 24337 30065 24349 30099
rect 24383 30096 24395 30099
rect 24518 30096 24524 30108
rect 24383 30068 24524 30096
rect 24383 30065 24395 30068
rect 24337 30059 24395 30065
rect 24518 30056 24524 30068
rect 24576 30056 24582 30108
rect 24610 30056 24616 30108
rect 24668 30096 24674 30108
rect 25809 30099 25867 30105
rect 25809 30096 25821 30099
rect 24668 30068 25821 30096
rect 24668 30056 24674 30068
rect 25809 30065 25821 30068
rect 25855 30096 25867 30099
rect 27830 30096 27836 30108
rect 25855 30068 27836 30096
rect 25855 30065 25867 30068
rect 25809 30059 25867 30065
rect 27830 30056 27836 30068
rect 27888 30096 27894 30108
rect 28017 30099 28075 30105
rect 28017 30096 28029 30099
rect 27888 30068 28029 30096
rect 27888 30056 27894 30068
rect 28017 30065 28029 30068
rect 28063 30096 28075 30099
rect 29305 30099 29363 30105
rect 29305 30096 29317 30099
rect 28063 30068 29317 30096
rect 28063 30065 28075 30068
rect 28017 30059 28075 30065
rect 29305 30065 29317 30068
rect 29351 30096 29363 30099
rect 29854 30096 29860 30108
rect 29351 30068 29860 30096
rect 29351 30065 29363 30068
rect 29305 30059 29363 30065
rect 29854 30056 29860 30068
rect 29912 30056 29918 30108
rect 3174 29988 3180 30040
rect 3232 30028 3238 30040
rect 3545 30031 3603 30037
rect 3545 30028 3557 30031
rect 3232 30000 3557 30028
rect 3232 29988 3238 30000
rect 3545 29997 3557 30000
rect 3591 29997 3603 30031
rect 4646 30028 4652 30040
rect 4607 30000 4652 30028
rect 3545 29991 3603 29997
rect 4646 29988 4652 30000
rect 4704 29988 4710 30040
rect 5382 29988 5388 30040
rect 5440 30028 5446 30040
rect 6673 30031 6731 30037
rect 6673 30028 6685 30031
rect 5440 30000 6685 30028
rect 5440 29988 5446 30000
rect 6673 29997 6685 30000
rect 6719 30028 6731 30031
rect 6854 30028 6860 30040
rect 6719 30000 6860 30028
rect 6719 29997 6731 30000
rect 6673 29991 6731 29997
rect 6854 29988 6860 30000
rect 6912 29988 6918 30040
rect 10994 30028 11000 30040
rect 10955 30000 11000 30028
rect 10994 29988 11000 30000
rect 11052 29988 11058 30040
rect 12282 29988 12288 30040
rect 12340 30028 12346 30040
rect 12745 30031 12803 30037
rect 12745 30028 12757 30031
rect 12340 30000 12757 30028
rect 12340 29988 12346 30000
rect 12745 29997 12757 30000
rect 12791 29997 12803 30031
rect 16146 30028 16152 30040
rect 16107 30000 16152 30028
rect 12745 29991 12803 29997
rect 16146 29988 16152 30000
rect 16204 29988 16210 30040
rect 16422 30028 16428 30040
rect 16383 30000 16428 30028
rect 16422 29988 16428 30000
rect 16480 29988 16486 30040
rect 18173 30031 18231 30037
rect 18173 29997 18185 30031
rect 18219 30028 18231 30031
rect 18262 30028 18268 30040
rect 18219 30000 18268 30028
rect 18219 29997 18231 30000
rect 18173 29991 18231 29997
rect 18262 29988 18268 30000
rect 18320 29988 18326 30040
rect 23325 30031 23383 30037
rect 23325 29997 23337 30031
rect 23371 30028 23383 30031
rect 23598 30028 23604 30040
rect 23371 30000 23604 30028
rect 23371 29997 23383 30000
rect 23325 29991 23383 29997
rect 23598 29988 23604 30000
rect 23656 29988 23662 30040
rect 25990 30028 25996 30040
rect 25951 30000 25996 30028
rect 25990 29988 25996 30000
rect 26048 29988 26054 30040
rect 27646 29988 27652 30040
rect 27704 30028 27710 30040
rect 28201 30031 28259 30037
rect 28201 30028 28213 30031
rect 27704 30000 28213 30028
rect 27704 29988 27710 30000
rect 28201 29997 28213 30000
rect 28247 29997 28259 30031
rect 28201 29991 28259 29997
rect 28661 30031 28719 30037
rect 28661 29997 28673 30031
rect 28707 30028 28719 30031
rect 29394 30028 29400 30040
rect 28707 30000 29400 30028
rect 28707 29997 28719 30000
rect 28661 29991 28719 29997
rect 29394 29988 29400 30000
rect 29452 30028 29458 30040
rect 29489 30031 29547 30037
rect 29489 30028 29501 30031
rect 29452 30000 29501 30028
rect 29452 29988 29458 30000
rect 29489 29997 29501 30000
rect 29535 29997 29547 30031
rect 29489 29991 29547 29997
rect 1061 29963 1119 29969
rect 1061 29929 1073 29963
rect 1107 29960 1119 29963
rect 1150 29960 1156 29972
rect 1107 29932 1156 29960
rect 1107 29929 1119 29932
rect 1061 29923 1119 29929
rect 1150 29920 1156 29932
rect 1208 29920 1214 29972
rect 13018 29920 13024 29972
rect 13076 29960 13082 29972
rect 13297 29963 13355 29969
rect 13297 29960 13309 29963
rect 13076 29932 13309 29960
rect 13076 29920 13082 29932
rect 13297 29929 13309 29932
rect 13343 29929 13355 29963
rect 23414 29960 23420 29972
rect 13297 29923 13355 29929
rect 18372 29932 23420 29960
rect 1242 29892 1248 29904
rect 1155 29864 1248 29892
rect 1242 29852 1248 29864
rect 1300 29892 1306 29904
rect 4646 29892 4652 29904
rect 1300 29864 4652 29892
rect 1300 29852 1306 29864
rect 4646 29852 4652 29864
rect 4704 29852 4710 29904
rect 13202 29892 13208 29904
rect 13163 29864 13208 29892
rect 13202 29852 13208 29864
rect 13260 29852 13266 29904
rect 16238 29852 16244 29904
rect 16296 29892 16302 29904
rect 18372 29892 18400 29932
rect 23414 29920 23420 29932
rect 23472 29960 23478 29972
rect 24521 29963 24579 29969
rect 24521 29960 24533 29963
rect 23472 29932 24533 29960
rect 23472 29920 23478 29932
rect 24521 29929 24533 29932
rect 24567 29929 24579 29963
rect 24521 29923 24579 29929
rect 20654 29892 20660 29904
rect 16296 29864 18400 29892
rect 20615 29864 20660 29892
rect 16296 29852 16302 29864
rect 20654 29852 20660 29864
rect 20712 29852 20718 29904
rect 23782 29852 23788 29904
rect 23840 29892 23846 29904
rect 24153 29895 24211 29901
rect 24153 29892 24165 29895
rect 23840 29864 24165 29892
rect 23840 29852 23846 29864
rect 24153 29861 24165 29864
rect 24199 29861 24211 29895
rect 24153 29855 24211 29861
rect 400 29802 31680 29824
rect 400 29750 3510 29802
rect 3562 29750 3574 29802
rect 3626 29750 3638 29802
rect 3690 29750 3702 29802
rect 3754 29750 3766 29802
rect 3818 29750 31680 29802
rect 400 29728 31680 29750
rect 2346 29648 2352 29700
rect 2404 29688 2410 29700
rect 3174 29688 3180 29700
rect 2404 29660 3180 29688
rect 2404 29648 2410 29660
rect 3174 29648 3180 29660
rect 3232 29648 3238 29700
rect 3358 29688 3364 29700
rect 3271 29660 3364 29688
rect 3358 29648 3364 29660
rect 3416 29688 3422 29700
rect 4281 29691 4339 29697
rect 4281 29688 4293 29691
rect 3416 29660 4293 29688
rect 3416 29648 3422 29660
rect 4281 29657 4293 29660
rect 4327 29657 4339 29691
rect 5014 29688 5020 29700
rect 4975 29660 5020 29688
rect 4281 29651 4339 29657
rect 5014 29648 5020 29660
rect 5072 29648 5078 29700
rect 7682 29688 7688 29700
rect 7643 29660 7688 29688
rect 7682 29648 7688 29660
rect 7740 29648 7746 29700
rect 8970 29648 8976 29700
rect 9028 29688 9034 29700
rect 9525 29691 9583 29697
rect 9525 29688 9537 29691
rect 9028 29660 9537 29688
rect 9028 29648 9034 29660
rect 9525 29657 9537 29660
rect 9571 29688 9583 29691
rect 10350 29688 10356 29700
rect 9571 29660 10356 29688
rect 9571 29657 9583 29660
rect 9525 29651 9583 29657
rect 10350 29648 10356 29660
rect 10408 29648 10414 29700
rect 16238 29688 16244 29700
rect 10460 29660 16244 29688
rect 4741 29623 4799 29629
rect 4741 29589 4753 29623
rect 4787 29620 4799 29623
rect 5382 29620 5388 29632
rect 4787 29592 5388 29620
rect 4787 29589 4799 29592
rect 4741 29583 4799 29589
rect 5382 29580 5388 29592
rect 5440 29580 5446 29632
rect 5474 29580 5480 29632
rect 5532 29620 5538 29632
rect 10460 29620 10488 29660
rect 16238 29648 16244 29660
rect 16296 29648 16302 29700
rect 16422 29648 16428 29700
rect 16480 29688 16486 29700
rect 16517 29691 16575 29697
rect 16517 29688 16529 29691
rect 16480 29660 16529 29688
rect 16480 29648 16486 29660
rect 16517 29657 16529 29660
rect 16563 29688 16575 29691
rect 16885 29691 16943 29697
rect 16885 29688 16897 29691
rect 16563 29660 16897 29688
rect 16563 29657 16575 29660
rect 16517 29651 16575 29657
rect 16885 29657 16897 29660
rect 16931 29657 16943 29691
rect 18998 29688 19004 29700
rect 18959 29660 19004 29688
rect 16885 29651 16943 29657
rect 5532 29592 10488 29620
rect 5532 29580 5538 29592
rect 969 29555 1027 29561
rect 969 29521 981 29555
rect 1015 29552 1027 29555
rect 1242 29552 1248 29564
rect 1015 29524 1248 29552
rect 1015 29521 1027 29524
rect 969 29515 1027 29521
rect 1242 29512 1248 29524
rect 1300 29512 1306 29564
rect 3821 29555 3879 29561
rect 3821 29521 3833 29555
rect 3867 29552 3879 29555
rect 4554 29552 4560 29564
rect 3867 29524 4560 29552
rect 3867 29521 3879 29524
rect 3821 29515 3879 29521
rect 4554 29512 4560 29524
rect 4612 29512 4618 29564
rect 9433 29555 9491 29561
rect 9433 29521 9445 29555
rect 9479 29552 9491 29555
rect 10258 29552 10264 29564
rect 9479 29524 10264 29552
rect 9479 29521 9491 29524
rect 9433 29515 9491 29521
rect 10258 29512 10264 29524
rect 10316 29552 10322 29564
rect 10537 29555 10595 29561
rect 10537 29552 10549 29555
rect 10316 29524 10549 29552
rect 10316 29512 10322 29524
rect 10537 29521 10549 29524
rect 10583 29521 10595 29555
rect 10537 29515 10595 29521
rect 10902 29512 10908 29564
rect 10960 29552 10966 29564
rect 11733 29555 11791 29561
rect 11733 29552 11745 29555
rect 10960 29524 11745 29552
rect 10960 29512 10966 29524
rect 11733 29521 11745 29524
rect 11779 29552 11791 29555
rect 12009 29555 12067 29561
rect 12009 29552 12021 29555
rect 11779 29524 12021 29552
rect 11779 29521 11791 29524
rect 11733 29515 11791 29521
rect 12009 29521 12021 29524
rect 12055 29521 12067 29555
rect 12558 29552 12564 29564
rect 12471 29524 12564 29552
rect 12009 29515 12067 29521
rect 12558 29512 12564 29524
rect 12616 29552 12622 29564
rect 13662 29552 13668 29564
rect 12616 29524 13668 29552
rect 12616 29512 12622 29524
rect 13662 29512 13668 29524
rect 13720 29512 13726 29564
rect 15502 29512 15508 29564
rect 15560 29552 15566 29564
rect 16425 29555 16483 29561
rect 16425 29552 16437 29555
rect 15560 29524 16437 29552
rect 15560 29512 15566 29524
rect 16425 29521 16437 29524
rect 16471 29552 16483 29555
rect 16900 29552 16928 29651
rect 18998 29648 19004 29660
rect 19056 29648 19062 29700
rect 20470 29688 20476 29700
rect 20431 29660 20476 29688
rect 20470 29648 20476 29660
rect 20528 29648 20534 29700
rect 23046 29688 23052 29700
rect 23007 29660 23052 29688
rect 23046 29648 23052 29660
rect 23104 29648 23110 29700
rect 23230 29648 23236 29700
rect 23288 29688 23294 29700
rect 23325 29691 23383 29697
rect 23325 29688 23337 29691
rect 23288 29660 23337 29688
rect 23288 29648 23294 29660
rect 23325 29657 23337 29660
rect 23371 29688 23383 29691
rect 23417 29691 23475 29697
rect 23417 29688 23429 29691
rect 23371 29660 23429 29688
rect 23371 29657 23383 29660
rect 23325 29651 23383 29657
rect 23417 29657 23429 29660
rect 23463 29657 23475 29691
rect 23598 29688 23604 29700
rect 23559 29660 23604 29688
rect 23417 29651 23475 29657
rect 23598 29648 23604 29660
rect 23656 29688 23662 29700
rect 24150 29688 24156 29700
rect 23656 29660 24156 29688
rect 23656 29648 23662 29660
rect 24150 29648 24156 29660
rect 24208 29648 24214 29700
rect 26910 29688 26916 29700
rect 26871 29660 26916 29688
rect 26910 29648 26916 29660
rect 26968 29648 26974 29700
rect 27830 29688 27836 29700
rect 27791 29660 27836 29688
rect 27830 29648 27836 29660
rect 27888 29648 27894 29700
rect 17161 29623 17219 29629
rect 17161 29589 17173 29623
rect 17207 29620 17219 29623
rect 18262 29620 18268 29632
rect 17207 29592 18268 29620
rect 17207 29589 17219 29592
rect 17161 29583 17219 29589
rect 17345 29555 17403 29561
rect 17345 29552 17357 29555
rect 16471 29524 16836 29552
rect 16900 29524 17357 29552
rect 16471 29521 16483 29524
rect 16425 29515 16483 29521
rect 16808 29496 16836 29524
rect 17345 29521 17357 29524
rect 17391 29521 17403 29555
rect 17345 29515 17403 29521
rect 2346 29444 2352 29496
rect 2404 29444 2410 29496
rect 4094 29484 4100 29496
rect 4055 29456 4100 29484
rect 4094 29444 4100 29456
rect 4152 29444 4158 29496
rect 6210 29444 6216 29496
rect 6268 29484 6274 29496
rect 7225 29487 7283 29493
rect 7225 29484 7237 29487
rect 6268 29456 7237 29484
rect 6268 29444 6274 29456
rect 7225 29453 7237 29456
rect 7271 29453 7283 29487
rect 7225 29447 7283 29453
rect 1150 29376 1156 29428
rect 1208 29416 1214 29428
rect 1245 29419 1303 29425
rect 1245 29416 1257 29419
rect 1208 29388 1257 29416
rect 1208 29376 1214 29388
rect 1245 29385 1257 29388
rect 1291 29385 1303 29419
rect 2993 29419 3051 29425
rect 2993 29406 3005 29419
rect 3039 29406 3051 29419
rect 4005 29419 4063 29425
rect 4005 29416 4017 29419
rect 2990 29394 2996 29406
rect 1245 29379 1303 29385
rect 2916 29366 2996 29394
rect 877 29351 935 29357
rect 877 29317 889 29351
rect 923 29348 935 29351
rect 2916 29348 2944 29366
rect 2990 29354 2996 29366
rect 3048 29354 3054 29406
rect 3468 29388 4017 29416
rect 923 29320 2944 29348
rect 923 29317 935 29320
rect 877 29311 935 29317
rect 3266 29308 3272 29360
rect 3324 29348 3330 29360
rect 3468 29357 3496 29388
rect 4005 29385 4017 29388
rect 4051 29385 4063 29419
rect 4005 29379 4063 29385
rect 4925 29419 4983 29425
rect 4925 29385 4937 29419
rect 4971 29416 4983 29419
rect 5290 29416 5296 29428
rect 4971 29388 5296 29416
rect 4971 29385 4983 29388
rect 4925 29379 4983 29385
rect 5290 29376 5296 29388
rect 5348 29376 5354 29428
rect 7240 29416 7268 29447
rect 7314 29444 7320 29496
rect 7372 29484 7378 29496
rect 7593 29487 7651 29493
rect 7593 29484 7605 29487
rect 7372 29456 7605 29484
rect 7372 29444 7378 29456
rect 7593 29453 7605 29456
rect 7639 29484 7651 29487
rect 8145 29487 8203 29493
rect 8145 29484 8157 29487
rect 7639 29456 8157 29484
rect 7639 29453 7651 29456
rect 7593 29447 7651 29453
rect 8145 29453 8157 29456
rect 8191 29484 8203 29487
rect 8970 29484 8976 29496
rect 8191 29456 8976 29484
rect 8191 29453 8203 29456
rect 8145 29447 8203 29453
rect 8970 29444 8976 29456
rect 9028 29444 9034 29496
rect 9982 29484 9988 29496
rect 9943 29456 9988 29484
rect 9982 29444 9988 29456
rect 10040 29484 10046 29496
rect 10721 29487 10779 29493
rect 10721 29484 10733 29487
rect 10040 29456 10733 29484
rect 10040 29444 10046 29456
rect 10721 29453 10733 29456
rect 10767 29484 10779 29487
rect 11822 29484 11828 29496
rect 10767 29456 11828 29484
rect 10767 29453 10779 29456
rect 10721 29447 10779 29453
rect 11822 29444 11828 29456
rect 11880 29484 11886 29496
rect 12282 29484 12288 29496
rect 11880 29456 12288 29484
rect 11880 29444 11886 29456
rect 12282 29444 12288 29456
rect 12340 29444 12346 29496
rect 13018 29484 13024 29496
rect 12576 29456 13024 29484
rect 7869 29419 7927 29425
rect 7869 29416 7881 29419
rect 7240 29388 7881 29416
rect 7869 29385 7881 29388
rect 7915 29416 7927 29419
rect 8786 29416 8792 29428
rect 7915 29388 8792 29416
rect 7915 29385 7927 29388
rect 7869 29379 7927 29385
rect 8786 29376 8792 29388
rect 8844 29376 8850 29428
rect 9062 29416 9068 29428
rect 9023 29388 9068 29416
rect 9062 29376 9068 29388
rect 9120 29376 9126 29428
rect 10350 29376 10356 29428
rect 10408 29416 10414 29428
rect 12576 29416 12604 29456
rect 13018 29444 13024 29456
rect 13076 29444 13082 29496
rect 15962 29484 15968 29496
rect 15923 29456 15968 29484
rect 15962 29444 15968 29456
rect 16020 29484 16026 29496
rect 16701 29487 16759 29493
rect 16701 29484 16713 29487
rect 16020 29456 16713 29484
rect 16020 29444 16026 29456
rect 16701 29453 16713 29456
rect 16747 29453 16759 29487
rect 16701 29447 16759 29453
rect 16790 29444 16796 29496
rect 16848 29484 16854 29496
rect 17452 29484 17480 29592
rect 18262 29580 18268 29592
rect 18320 29580 18326 29632
rect 17618 29512 17624 29564
rect 17676 29552 17682 29564
rect 18449 29555 18507 29561
rect 18449 29552 18461 29555
rect 17676 29524 18461 29552
rect 17676 29512 17682 29524
rect 17894 29484 17900 29496
rect 16848 29456 17480 29484
rect 17855 29456 17900 29484
rect 16848 29444 16854 29456
rect 17894 29444 17900 29456
rect 17952 29444 17958 29496
rect 18188 29493 18216 29524
rect 18449 29521 18461 29524
rect 18495 29521 18507 29555
rect 18449 29515 18507 29521
rect 24061 29555 24119 29561
rect 24061 29521 24073 29555
rect 24107 29552 24119 29555
rect 24518 29552 24524 29564
rect 24107 29524 24524 29552
rect 24107 29521 24119 29524
rect 24061 29515 24119 29521
rect 24518 29512 24524 29524
rect 24576 29552 24582 29564
rect 26450 29552 26456 29564
rect 24576 29524 26456 29552
rect 24576 29512 24582 29524
rect 26450 29512 26456 29524
rect 26508 29512 26514 29564
rect 18173 29487 18231 29493
rect 18173 29453 18185 29487
rect 18219 29453 18231 29487
rect 18173 29447 18231 29453
rect 18262 29444 18268 29496
rect 18320 29484 18326 29496
rect 18357 29487 18415 29493
rect 18357 29484 18369 29487
rect 18320 29456 18369 29484
rect 18320 29444 18326 29456
rect 18357 29453 18369 29456
rect 18403 29453 18415 29487
rect 19550 29484 19556 29496
rect 19511 29456 19556 29484
rect 18357 29447 18415 29453
rect 19550 29444 19556 29456
rect 19608 29484 19614 29496
rect 20105 29487 20163 29493
rect 20105 29484 20117 29487
rect 19608 29456 20117 29484
rect 19608 29444 19614 29456
rect 20105 29453 20117 29456
rect 20151 29484 20163 29487
rect 20565 29487 20623 29493
rect 20565 29484 20577 29487
rect 20151 29456 20577 29484
rect 20151 29453 20163 29456
rect 20105 29447 20163 29453
rect 20565 29453 20577 29456
rect 20611 29484 20623 29487
rect 20654 29484 20660 29496
rect 20611 29456 20660 29484
rect 20611 29453 20623 29456
rect 20565 29447 20623 29453
rect 20654 29444 20660 29456
rect 20712 29484 20718 29496
rect 20841 29487 20899 29493
rect 20841 29484 20853 29487
rect 20712 29456 20853 29484
rect 20712 29444 20718 29456
rect 20841 29453 20853 29456
rect 20887 29484 20899 29487
rect 21393 29487 21451 29493
rect 21393 29484 21405 29487
rect 20887 29456 21405 29484
rect 20887 29453 20899 29456
rect 20841 29447 20899 29453
rect 21393 29453 21405 29456
rect 21439 29453 21451 29487
rect 24150 29484 24156 29496
rect 24111 29456 24156 29484
rect 21393 29447 21451 29453
rect 24150 29444 24156 29456
rect 24208 29444 24214 29496
rect 26928 29484 26956 29648
rect 28569 29555 28627 29561
rect 28569 29521 28581 29555
rect 28615 29552 28627 29555
rect 28842 29552 28848 29564
rect 28615 29524 28848 29552
rect 28615 29521 28627 29524
rect 28569 29515 28627 29521
rect 28842 29512 28848 29524
rect 28900 29512 28906 29564
rect 27005 29487 27063 29493
rect 27005 29484 27017 29487
rect 26928 29456 27017 29484
rect 27005 29453 27017 29456
rect 27051 29484 27063 29487
rect 27830 29484 27836 29496
rect 27051 29456 27836 29484
rect 27051 29453 27063 29456
rect 27005 29447 27063 29453
rect 27830 29444 27836 29456
rect 27888 29444 27894 29496
rect 10408 29388 12604 29416
rect 12745 29419 12803 29425
rect 10408 29376 10414 29388
rect 12745 29385 12757 29419
rect 12791 29416 12803 29419
rect 13294 29416 13300 29428
rect 12791 29388 13300 29416
rect 12791 29385 12803 29388
rect 12745 29379 12803 29385
rect 13294 29376 13300 29388
rect 13352 29376 13358 29428
rect 15042 29416 15048 29428
rect 3453 29351 3511 29357
rect 3453 29348 3465 29351
rect 3324 29320 3465 29348
rect 3324 29308 3330 29320
rect 3453 29317 3465 29320
rect 3499 29317 3511 29351
rect 3453 29311 3511 29317
rect 3729 29351 3787 29357
rect 3729 29317 3741 29351
rect 3775 29348 3787 29351
rect 4186 29348 4192 29360
rect 3775 29320 4192 29348
rect 3775 29317 3787 29320
rect 3729 29311 3787 29317
rect 4186 29308 4192 29320
rect 4244 29348 4250 29360
rect 4554 29348 4560 29360
rect 4244 29320 4560 29348
rect 4244 29308 4250 29320
rect 4554 29308 4560 29320
rect 4612 29308 4618 29360
rect 4646 29308 4652 29360
rect 4704 29348 4710 29360
rect 5201 29351 5259 29357
rect 5201 29348 5213 29351
rect 4704 29320 5213 29348
rect 4704 29308 4710 29320
rect 5201 29317 5213 29320
rect 5247 29348 5259 29351
rect 6302 29348 6308 29360
rect 5247 29320 6308 29348
rect 5247 29317 5259 29320
rect 5201 29311 5259 29317
rect 6302 29308 6308 29320
rect 6360 29308 6366 29360
rect 9154 29348 9160 29360
rect 9115 29320 9160 29348
rect 9154 29308 9160 29320
rect 9212 29308 9218 29360
rect 12929 29351 12987 29357
rect 12929 29317 12941 29351
rect 12975 29348 12987 29351
rect 13110 29348 13116 29360
rect 12975 29320 13116 29348
rect 12975 29317 12987 29320
rect 12929 29311 12987 29317
rect 13110 29308 13116 29320
rect 13168 29308 13174 29360
rect 13202 29308 13208 29360
rect 13260 29348 13266 29360
rect 14324 29348 14352 29416
rect 15003 29388 15048 29416
rect 15042 29376 15048 29388
rect 15100 29376 15106 29428
rect 15410 29376 15416 29428
rect 15468 29416 15474 29428
rect 15781 29419 15839 29425
rect 15781 29416 15793 29419
rect 15468 29388 15793 29416
rect 15468 29376 15474 29388
rect 15781 29385 15793 29388
rect 15827 29416 15839 29419
rect 16241 29419 16299 29425
rect 16241 29416 16253 29419
rect 15827 29388 16253 29416
rect 15827 29385 15839 29388
rect 15781 29379 15839 29385
rect 16241 29385 16253 29388
rect 16287 29416 16299 29419
rect 17618 29416 17624 29428
rect 16287 29388 17624 29416
rect 16287 29385 16299 29388
rect 16241 29379 16299 29385
rect 17618 29376 17624 29388
rect 17676 29376 17682 29428
rect 19829 29419 19887 29425
rect 19829 29385 19841 29419
rect 19875 29385 19887 29419
rect 21114 29416 21120 29428
rect 21075 29388 21120 29416
rect 19829 29379 19887 29385
rect 13260 29320 14352 29348
rect 15597 29351 15655 29357
rect 13260 29308 13266 29320
rect 15597 29317 15609 29351
rect 15643 29348 15655 29351
rect 16146 29348 16152 29360
rect 15643 29320 16152 29348
rect 15643 29317 15655 29320
rect 15597 29311 15655 29317
rect 16146 29308 16152 29320
rect 16204 29348 16210 29360
rect 17342 29348 17348 29360
rect 16204 29320 17348 29348
rect 16204 29308 16210 29320
rect 17342 29308 17348 29320
rect 17400 29308 17406 29360
rect 18354 29308 18360 29360
rect 18412 29348 18418 29360
rect 19461 29351 19519 29357
rect 19461 29348 19473 29351
rect 18412 29320 19473 29348
rect 18412 29308 18418 29320
rect 19461 29317 19473 29320
rect 19507 29348 19519 29351
rect 19844 29348 19872 29379
rect 21114 29376 21120 29388
rect 21172 29416 21178 29428
rect 21577 29419 21635 29425
rect 21577 29416 21589 29419
rect 21172 29388 21589 29416
rect 21172 29376 21178 29388
rect 21577 29385 21589 29388
rect 21623 29385 21635 29419
rect 21577 29379 21635 29385
rect 23874 29376 23880 29428
rect 23932 29416 23938 29428
rect 24429 29419 24487 29425
rect 24429 29416 24441 29419
rect 23932 29388 24441 29416
rect 23932 29376 23938 29388
rect 24429 29385 24441 29388
rect 24475 29416 24487 29419
rect 24518 29416 24524 29428
rect 24475 29388 24524 29416
rect 24475 29385 24487 29388
rect 24429 29379 24487 29385
rect 24518 29376 24524 29388
rect 24576 29376 24582 29428
rect 24886 29376 24892 29428
rect 24944 29376 24950 29428
rect 26082 29376 26088 29428
rect 26140 29416 26146 29428
rect 26177 29419 26235 29425
rect 26177 29416 26189 29419
rect 26140 29388 26189 29416
rect 26140 29376 26146 29388
rect 26177 29385 26189 29388
rect 26223 29385 26235 29419
rect 26177 29379 26235 29385
rect 26910 29376 26916 29428
rect 26968 29416 26974 29428
rect 27281 29419 27339 29425
rect 27281 29416 27293 29419
rect 26968 29388 27293 29416
rect 26968 29376 26974 29388
rect 27281 29385 27293 29388
rect 27327 29416 27339 29419
rect 27557 29419 27615 29425
rect 27557 29416 27569 29419
rect 27327 29388 27569 29416
rect 27327 29385 27339 29388
rect 27281 29379 27339 29385
rect 27557 29385 27569 29388
rect 27603 29385 27615 29419
rect 27557 29379 27615 29385
rect 27646 29376 27652 29428
rect 27704 29416 27710 29428
rect 27925 29419 27983 29425
rect 27925 29416 27937 29419
rect 27704 29388 27937 29416
rect 27704 29376 27710 29388
rect 27925 29385 27937 29388
rect 27971 29385 27983 29419
rect 28198 29416 28204 29428
rect 28111 29388 28204 29416
rect 27925 29379 27983 29385
rect 28198 29376 28204 29388
rect 28256 29416 28262 29428
rect 28845 29419 28903 29425
rect 28845 29416 28857 29419
rect 28256 29388 28857 29416
rect 28256 29376 28262 29388
rect 28845 29385 28857 29388
rect 28891 29385 28903 29419
rect 28845 29379 28903 29385
rect 29394 29376 29400 29428
rect 29452 29376 29458 29428
rect 30593 29419 30651 29425
rect 30593 29385 30605 29419
rect 30639 29385 30651 29419
rect 30593 29379 30651 29385
rect 20102 29348 20108 29360
rect 19507 29320 20108 29348
rect 19507 29317 19519 29320
rect 19461 29311 19519 29317
rect 20102 29308 20108 29320
rect 20160 29308 20166 29360
rect 23690 29308 23696 29360
rect 23748 29348 23754 29360
rect 23785 29351 23843 29357
rect 23785 29348 23797 29351
rect 23748 29320 23797 29348
rect 23748 29308 23754 29320
rect 23785 29317 23797 29320
rect 23831 29317 23843 29351
rect 24904 29348 24932 29376
rect 25990 29348 25996 29360
rect 24904 29320 25996 29348
rect 23785 29311 23843 29317
rect 25990 29308 25996 29320
rect 26048 29348 26054 29360
rect 26269 29351 26327 29357
rect 26269 29348 26281 29351
rect 26048 29320 26281 29348
rect 26048 29308 26054 29320
rect 26269 29317 26281 29320
rect 26315 29317 26327 29351
rect 26269 29311 26327 29317
rect 26545 29351 26603 29357
rect 26545 29317 26557 29351
rect 26591 29348 26603 29351
rect 27738 29348 27744 29360
rect 26591 29320 27744 29348
rect 26591 29317 26603 29320
rect 26545 29311 26603 29317
rect 27738 29308 27744 29320
rect 27796 29308 27802 29360
rect 28385 29351 28443 29357
rect 28385 29317 28397 29351
rect 28431 29348 28443 29351
rect 28474 29348 28480 29360
rect 28431 29320 28480 29348
rect 28431 29317 28443 29320
rect 28385 29311 28443 29317
rect 28474 29308 28480 29320
rect 28532 29348 28538 29360
rect 30608 29348 30636 29379
rect 28532 29320 30636 29348
rect 28532 29308 28538 29320
rect 400 29258 31680 29280
rect 400 29206 18870 29258
rect 18922 29206 18934 29258
rect 18986 29206 18998 29258
rect 19050 29206 19062 29258
rect 19114 29206 19126 29258
rect 19178 29206 31680 29258
rect 400 29184 31680 29206
rect 1061 29147 1119 29153
rect 1061 29113 1073 29147
rect 1107 29144 1119 29147
rect 2346 29144 2352 29156
rect 1107 29116 2352 29144
rect 1107 29113 1119 29116
rect 1061 29107 1119 29113
rect 2346 29104 2352 29116
rect 2404 29104 2410 29156
rect 3913 29147 3971 29153
rect 3913 29113 3925 29147
rect 3959 29144 3971 29147
rect 4094 29144 4100 29156
rect 3959 29116 4100 29144
rect 3959 29113 3971 29116
rect 3913 29107 3971 29113
rect 4094 29104 4100 29116
rect 4152 29104 4158 29156
rect 4462 29104 4468 29156
rect 4520 29144 4526 29156
rect 5290 29144 5296 29156
rect 4520 29116 5296 29144
rect 4520 29104 4526 29116
rect 5290 29104 5296 29116
rect 5348 29104 5354 29156
rect 16241 29147 16299 29153
rect 16241 29113 16253 29147
rect 16287 29144 16299 29147
rect 16882 29144 16888 29156
rect 16287 29116 16888 29144
rect 16287 29113 16299 29116
rect 16241 29107 16299 29113
rect 16882 29104 16888 29116
rect 16940 29104 16946 29156
rect 17894 29144 17900 29156
rect 16992 29116 17900 29144
rect 4557 29079 4615 29085
rect 4557 29045 4569 29079
rect 4603 29076 4615 29079
rect 4603 29048 5704 29076
rect 4603 29045 4615 29048
rect 4557 29039 4615 29045
rect 5676 29020 5704 29048
rect 13294 29036 13300 29088
rect 13352 29076 13358 29088
rect 15226 29076 15232 29088
rect 13352 29048 14214 29076
rect 13352 29036 13358 29048
rect 2990 28968 2996 29020
rect 3048 29008 3054 29020
rect 3637 29011 3695 29017
rect 3637 29008 3649 29011
rect 3048 28980 3649 29008
rect 3048 28968 3054 28980
rect 3637 28977 3649 28980
rect 3683 29008 3695 29011
rect 4002 29008 4008 29020
rect 3683 28980 4008 29008
rect 3683 28977 3695 28980
rect 3637 28971 3695 28977
rect 4002 28968 4008 28980
rect 4060 28968 4066 29020
rect 4278 28968 4284 29020
rect 4336 29008 4342 29020
rect 5017 29011 5075 29017
rect 5017 29008 5029 29011
rect 4336 28980 5029 29008
rect 4336 28968 4342 28980
rect 5017 28977 5029 28980
rect 5063 28977 5075 29011
rect 5658 29008 5664 29020
rect 5571 28980 5664 29008
rect 5017 28971 5075 28977
rect 5658 28968 5664 28980
rect 5716 28968 5722 29020
rect 6854 29008 6860 29020
rect 6815 28980 6860 29008
rect 6854 28968 6860 28980
rect 6912 28968 6918 29020
rect 8970 29008 8976 29020
rect 8931 28980 8976 29008
rect 8970 28968 8976 28980
rect 9028 28968 9034 29020
rect 9062 28968 9068 29020
rect 9120 29008 9126 29020
rect 9157 29011 9215 29017
rect 9157 29008 9169 29011
rect 9120 28980 9169 29008
rect 9120 28968 9126 28980
rect 9157 28977 9169 28980
rect 9203 29008 9215 29011
rect 10629 29011 10687 29017
rect 10629 29008 10641 29011
rect 9203 28980 10641 29008
rect 9203 28977 9215 28980
rect 9157 28971 9215 28977
rect 10629 28977 10641 28980
rect 10675 29008 10687 29011
rect 10994 29008 11000 29020
rect 10675 28980 11000 29008
rect 10675 28977 10687 28980
rect 10629 28971 10687 28977
rect 10994 28968 11000 28980
rect 11052 28968 11058 29020
rect 11822 29008 11828 29020
rect 11783 28980 11828 29008
rect 11822 28968 11828 28980
rect 11880 28968 11886 29020
rect 13113 29011 13171 29017
rect 13113 28977 13125 29011
rect 13159 29008 13171 29011
rect 13662 29008 13668 29020
rect 13159 28980 13668 29008
rect 13159 28977 13171 28980
rect 13113 28971 13171 28977
rect 13662 28968 13668 28980
rect 13720 28968 13726 29020
rect 4922 28940 4928 28952
rect 4883 28912 4928 28940
rect 4922 28900 4928 28912
rect 4980 28900 4986 28952
rect 5566 28940 5572 28952
rect 5527 28912 5572 28940
rect 5566 28900 5572 28912
rect 5624 28900 5630 28952
rect 11914 28900 11920 28952
rect 11972 28940 11978 28952
rect 12009 28943 12067 28949
rect 12009 28940 12021 28943
rect 11972 28912 12021 28940
rect 11972 28900 11978 28912
rect 12009 28909 12021 28912
rect 12055 28909 12067 28943
rect 13294 28940 13300 28952
rect 13255 28912 13300 28940
rect 12009 28903 12067 28909
rect 13294 28900 13300 28912
rect 13352 28900 13358 28952
rect 14186 28940 14214 29048
rect 15060 29048 15232 29076
rect 15060 29017 15088 29048
rect 15226 29036 15232 29048
rect 15284 29036 15290 29088
rect 15045 29011 15103 29017
rect 15045 28977 15057 29011
rect 15091 28977 15103 29011
rect 15318 29008 15324 29020
rect 15279 28980 15324 29008
rect 15045 28971 15103 28977
rect 15318 28968 15324 28980
rect 15376 28968 15382 29020
rect 15413 29011 15471 29017
rect 15413 28977 15425 29011
rect 15459 29008 15471 29011
rect 15502 29008 15508 29020
rect 15459 28980 15508 29008
rect 15459 28977 15471 28980
rect 15413 28971 15471 28977
rect 14582 28940 14588 28952
rect 14186 28912 14588 28940
rect 14582 28900 14588 28912
rect 14640 28900 14646 28952
rect 14674 28900 14680 28952
rect 14732 28940 14738 28952
rect 15428 28940 15456 28971
rect 15502 28968 15508 28980
rect 15560 28968 15566 29020
rect 16057 29011 16115 29017
rect 16057 28977 16069 29011
rect 16103 29008 16115 29011
rect 16146 29008 16152 29020
rect 16103 28980 16152 29008
rect 16103 28977 16115 28980
rect 16057 28971 16115 28977
rect 16146 28968 16152 28980
rect 16204 29008 16210 29020
rect 16992 29008 17020 29116
rect 17894 29104 17900 29116
rect 17952 29144 17958 29156
rect 18081 29147 18139 29153
rect 18081 29144 18093 29147
rect 17952 29116 18093 29144
rect 17952 29104 17958 29116
rect 18081 29113 18093 29116
rect 18127 29113 18139 29147
rect 24150 29144 24156 29156
rect 24111 29116 24156 29144
rect 18081 29107 18139 29113
rect 24150 29104 24156 29116
rect 24208 29104 24214 29156
rect 24613 29147 24671 29153
rect 24613 29113 24625 29147
rect 24659 29144 24671 29147
rect 24886 29144 24892 29156
rect 24659 29116 24892 29144
rect 24659 29113 24671 29116
rect 24613 29107 24671 29113
rect 24886 29104 24892 29116
rect 24944 29104 24950 29156
rect 29394 29144 29400 29156
rect 29355 29116 29400 29144
rect 29394 29104 29400 29116
rect 29452 29104 29458 29156
rect 29946 29144 29952 29156
rect 29907 29116 29952 29144
rect 29946 29104 29952 29116
rect 30004 29104 30010 29156
rect 17618 29076 17624 29088
rect 17084 29048 17624 29076
rect 17084 29017 17112 29048
rect 17618 29036 17624 29048
rect 17676 29036 17682 29088
rect 23414 29036 23420 29088
rect 23472 29076 23478 29088
rect 24337 29079 24395 29085
rect 24337 29076 24349 29079
rect 23472 29048 24349 29076
rect 23472 29036 23478 29048
rect 24337 29045 24349 29048
rect 24383 29045 24395 29079
rect 24337 29039 24395 29045
rect 27646 29036 27652 29088
rect 27704 29036 27710 29088
rect 16204 28980 17020 29008
rect 17069 29011 17127 29017
rect 16204 28968 16210 28980
rect 17069 28977 17081 29011
rect 17115 28977 17127 29011
rect 17069 28971 17127 28977
rect 17437 29011 17495 29017
rect 17437 28977 17449 29011
rect 17483 28977 17495 29011
rect 17437 28971 17495 28977
rect 14732 28912 15456 28940
rect 15689 28943 15747 28949
rect 14732 28900 14738 28912
rect 15689 28909 15701 28943
rect 15735 28909 15747 28943
rect 15689 28903 15747 28909
rect 5290 28872 5296 28884
rect 5251 28844 5296 28872
rect 5290 28832 5296 28844
rect 5348 28832 5354 28884
rect 7314 28872 7320 28884
rect 5768 28844 7320 28872
rect 1886 28804 1892 28816
rect 1847 28776 1892 28804
rect 1886 28764 1892 28776
rect 1944 28764 1950 28816
rect 2070 28804 2076 28816
rect 2031 28776 2076 28804
rect 2070 28764 2076 28776
rect 2128 28764 2134 28816
rect 3174 28764 3180 28816
rect 3232 28804 3238 28816
rect 3453 28807 3511 28813
rect 3453 28804 3465 28807
rect 3232 28776 3465 28804
rect 3232 28764 3238 28776
rect 3453 28773 3465 28776
rect 3499 28804 3511 28807
rect 4005 28807 4063 28813
rect 4005 28804 4017 28807
rect 3499 28776 4017 28804
rect 3499 28773 3511 28776
rect 3453 28767 3511 28773
rect 4005 28773 4017 28776
rect 4051 28773 4063 28807
rect 4005 28767 4063 28773
rect 4281 28807 4339 28813
rect 4281 28773 4293 28807
rect 4327 28804 4339 28807
rect 5014 28804 5020 28816
rect 4327 28776 5020 28804
rect 4327 28773 4339 28776
rect 4281 28767 4339 28773
rect 5014 28764 5020 28776
rect 5072 28804 5078 28816
rect 5768 28804 5796 28844
rect 7314 28832 7320 28844
rect 7372 28832 7378 28884
rect 8145 28875 8203 28881
rect 8145 28841 8157 28875
rect 8191 28872 8203 28875
rect 9522 28872 9528 28884
rect 8191 28844 9528 28872
rect 8191 28841 8203 28844
rect 8145 28835 8203 28841
rect 9522 28832 9528 28844
rect 9580 28832 9586 28884
rect 15042 28832 15048 28884
rect 15100 28872 15106 28884
rect 15704 28872 15732 28903
rect 16974 28872 16980 28884
rect 15100 28844 15732 28872
rect 16935 28844 16980 28872
rect 15100 28832 15106 28844
rect 16974 28832 16980 28844
rect 17032 28832 17038 28884
rect 17158 28832 17164 28884
rect 17216 28872 17222 28884
rect 17452 28872 17480 28971
rect 18722 28968 18728 29020
rect 18780 29008 18786 29020
rect 18909 29011 18967 29017
rect 18909 29008 18921 29011
rect 18780 28980 18921 29008
rect 18780 28968 18786 28980
rect 18909 28977 18921 28980
rect 18955 28977 18967 29011
rect 18909 28971 18967 28977
rect 20102 28968 20108 29020
rect 20160 29008 20166 29020
rect 20197 29011 20255 29017
rect 20197 29008 20209 29011
rect 20160 28980 20209 29008
rect 20160 28968 20166 28980
rect 20197 28977 20209 28980
rect 20243 28977 20255 29011
rect 20197 28971 20255 28977
rect 21114 28968 21120 29020
rect 21172 29008 21178 29020
rect 23506 29008 23512 29020
rect 21172 28980 23512 29008
rect 21172 28968 21178 28980
rect 23506 28968 23512 28980
rect 23564 28968 23570 29020
rect 26910 29008 26916 29020
rect 26871 28980 26916 29008
rect 26910 28968 26916 28980
rect 26968 28968 26974 29020
rect 29762 29008 29768 29020
rect 29723 28980 29768 29008
rect 29762 28968 29768 28980
rect 29820 28968 29826 29020
rect 17526 28900 17532 28952
rect 17584 28940 17590 28952
rect 17713 28943 17771 28949
rect 17713 28940 17725 28943
rect 17584 28912 17725 28940
rect 17584 28900 17590 28912
rect 17713 28909 17725 28912
rect 17759 28909 17771 28943
rect 17713 28903 17771 28909
rect 20286 28900 20292 28952
rect 20344 28940 20350 28952
rect 20381 28943 20439 28949
rect 20381 28940 20393 28943
rect 20344 28912 20393 28940
rect 20344 28900 20350 28912
rect 20381 28909 20393 28912
rect 20427 28909 20439 28943
rect 20381 28903 20439 28909
rect 23785 28943 23843 28949
rect 23785 28909 23797 28943
rect 23831 28940 23843 28943
rect 24610 28940 24616 28952
rect 23831 28912 24616 28940
rect 23831 28909 23843 28912
rect 23785 28903 23843 28909
rect 24610 28900 24616 28912
rect 24668 28900 24674 28952
rect 27186 28940 27192 28952
rect 27147 28912 27192 28940
rect 27186 28900 27192 28912
rect 27244 28900 27250 28952
rect 27278 28900 27284 28952
rect 27336 28940 27342 28952
rect 28937 28943 28995 28949
rect 28937 28940 28949 28943
rect 27336 28912 28949 28940
rect 27336 28900 27342 28912
rect 28937 28909 28949 28912
rect 28983 28909 28995 28943
rect 28937 28903 28995 28909
rect 17216 28844 19228 28872
rect 17216 28832 17222 28844
rect 6210 28804 6216 28816
rect 5072 28776 5796 28804
rect 6171 28776 6216 28804
rect 5072 28764 5078 28776
rect 6210 28764 6216 28776
rect 6268 28764 6274 28816
rect 6946 28804 6952 28816
rect 6907 28776 6952 28804
rect 6946 28764 6952 28776
rect 7004 28764 7010 28816
rect 8878 28764 8884 28816
rect 8936 28804 8942 28816
rect 9249 28807 9307 28813
rect 9249 28804 9261 28807
rect 8936 28776 9261 28804
rect 8936 28764 8942 28776
rect 9249 28773 9261 28776
rect 9295 28804 9307 28807
rect 9617 28807 9675 28813
rect 9617 28804 9629 28807
rect 9295 28776 9629 28804
rect 9295 28773 9307 28776
rect 9249 28767 9307 28773
rect 9617 28773 9629 28776
rect 9663 28773 9675 28807
rect 10442 28804 10448 28816
rect 10403 28776 10448 28804
rect 9617 28767 9675 28773
rect 10442 28764 10448 28776
rect 10500 28764 10506 28816
rect 18078 28764 18084 28816
rect 18136 28804 18142 28816
rect 19200 28813 19228 28844
rect 18265 28807 18323 28813
rect 18265 28804 18277 28807
rect 18136 28776 18277 28804
rect 18136 28764 18142 28776
rect 18265 28773 18277 28776
rect 18311 28773 18323 28807
rect 18265 28767 18323 28773
rect 19185 28807 19243 28813
rect 19185 28773 19197 28807
rect 19231 28804 19243 28807
rect 19274 28804 19280 28816
rect 19231 28776 19280 28804
rect 19231 28773 19243 28776
rect 19185 28767 19243 28773
rect 19274 28764 19280 28776
rect 19332 28764 19338 28816
rect 24981 28807 25039 28813
rect 24981 28773 24993 28807
rect 25027 28804 25039 28807
rect 26174 28804 26180 28816
rect 25027 28776 26180 28804
rect 25027 28773 25039 28776
rect 24981 28767 25039 28773
rect 26174 28764 26180 28776
rect 26232 28764 26238 28816
rect 29581 28807 29639 28813
rect 29581 28773 29593 28807
rect 29627 28804 29639 28807
rect 29854 28804 29860 28816
rect 29627 28776 29860 28804
rect 29627 28773 29639 28776
rect 29581 28767 29639 28773
rect 29854 28764 29860 28776
rect 29912 28764 29918 28816
rect 400 28714 31680 28736
rect 400 28662 3510 28714
rect 3562 28662 3574 28714
rect 3626 28662 3638 28714
rect 3690 28662 3702 28714
rect 3754 28662 3766 28714
rect 3818 28662 31680 28714
rect 400 28640 31680 28662
rect 1150 28560 1156 28612
rect 1208 28600 1214 28612
rect 1613 28603 1671 28609
rect 1613 28600 1625 28603
rect 1208 28572 1625 28600
rect 1208 28560 1214 28572
rect 1613 28569 1625 28572
rect 1659 28600 1671 28603
rect 4278 28600 4284 28612
rect 1659 28572 2208 28600
rect 4239 28572 4284 28600
rect 1659 28569 1671 28572
rect 1613 28563 1671 28569
rect 2180 28541 2208 28572
rect 4278 28560 4284 28572
rect 4336 28560 4342 28612
rect 5290 28600 5296 28612
rect 5251 28572 5296 28600
rect 5290 28560 5296 28572
rect 5348 28560 5354 28612
rect 5658 28600 5664 28612
rect 5619 28572 5664 28600
rect 5658 28560 5664 28572
rect 5716 28560 5722 28612
rect 6210 28560 6216 28612
rect 6268 28600 6274 28612
rect 6397 28603 6455 28609
rect 6397 28600 6409 28603
rect 6268 28572 6409 28600
rect 6268 28560 6274 28572
rect 6397 28569 6409 28572
rect 6443 28569 6455 28603
rect 6854 28600 6860 28612
rect 6815 28572 6860 28600
rect 6397 28563 6455 28569
rect 6854 28560 6860 28572
rect 6912 28560 6918 28612
rect 8970 28560 8976 28612
rect 9028 28600 9034 28612
rect 9709 28603 9767 28609
rect 9709 28600 9721 28603
rect 9028 28572 9721 28600
rect 9028 28560 9034 28572
rect 9709 28569 9721 28572
rect 9755 28569 9767 28603
rect 9709 28563 9767 28569
rect 10074 28560 10080 28612
rect 10132 28600 10138 28612
rect 12837 28603 12895 28609
rect 12837 28600 12849 28603
rect 10132 28572 12849 28600
rect 10132 28560 10138 28572
rect 12837 28569 12849 28572
rect 12883 28600 12895 28603
rect 13294 28600 13300 28612
rect 12883 28572 13300 28600
rect 12883 28569 12895 28572
rect 12837 28563 12895 28569
rect 2165 28535 2223 28541
rect 2165 28501 2177 28535
rect 2211 28501 2223 28535
rect 5477 28535 5535 28541
rect 5477 28532 5489 28535
rect 2165 28495 2223 28501
rect 4756 28504 5489 28532
rect 4756 28476 4784 28504
rect 5477 28501 5489 28504
rect 5523 28532 5535 28535
rect 5566 28532 5572 28544
rect 5523 28504 5572 28532
rect 5523 28501 5535 28504
rect 5477 28495 5535 28501
rect 5566 28492 5572 28504
rect 5624 28492 5630 28544
rect 7961 28535 8019 28541
rect 7961 28501 7973 28535
rect 8007 28532 8019 28535
rect 8421 28535 8479 28541
rect 8421 28532 8433 28535
rect 8007 28504 8433 28532
rect 8007 28501 8019 28504
rect 7961 28495 8019 28501
rect 8421 28501 8433 28504
rect 8467 28532 8479 28535
rect 9154 28532 9160 28544
rect 8467 28504 9160 28532
rect 8467 28501 8479 28504
rect 8421 28495 8479 28501
rect 9154 28492 9160 28504
rect 9212 28492 9218 28544
rect 9617 28535 9675 28541
rect 9617 28501 9629 28535
rect 9663 28532 9675 28535
rect 10994 28532 11000 28544
rect 9663 28504 11000 28532
rect 9663 28501 9675 28504
rect 9617 28495 9675 28501
rect 10994 28492 11000 28504
rect 11052 28492 11058 28544
rect 11822 28492 11828 28544
rect 11880 28532 11886 28544
rect 12009 28535 12067 28541
rect 12009 28532 12021 28535
rect 11880 28504 12021 28532
rect 11880 28492 11886 28504
rect 12009 28501 12021 28504
rect 12055 28501 12067 28535
rect 12009 28495 12067 28501
rect 1521 28467 1579 28473
rect 1521 28433 1533 28467
rect 1567 28464 1579 28467
rect 3085 28467 3143 28473
rect 3085 28464 3097 28467
rect 1567 28436 3097 28464
rect 1567 28433 1579 28436
rect 1521 28427 1579 28433
rect 3085 28433 3097 28436
rect 3131 28464 3143 28467
rect 4738 28464 4744 28476
rect 3131 28436 4744 28464
rect 3131 28433 3143 28436
rect 3085 28427 3143 28433
rect 4738 28424 4744 28436
rect 4796 28424 4802 28476
rect 4830 28424 4836 28476
rect 4888 28464 4894 28476
rect 4925 28467 4983 28473
rect 4925 28464 4937 28467
rect 4888 28436 4937 28464
rect 4888 28424 4894 28436
rect 4925 28433 4937 28436
rect 4971 28433 4983 28467
rect 4925 28427 4983 28433
rect 7682 28424 7688 28476
rect 7740 28464 7746 28476
rect 8237 28467 8295 28473
rect 8237 28464 8249 28467
rect 7740 28436 8249 28464
rect 7740 28424 7746 28436
rect 8237 28433 8249 28436
rect 8283 28433 8295 28467
rect 8237 28427 8295 28433
rect 9341 28467 9399 28473
rect 9341 28433 9353 28467
rect 9387 28464 9399 28467
rect 9522 28464 9528 28476
rect 9387 28436 9528 28464
rect 9387 28433 9399 28436
rect 9341 28427 9399 28433
rect 9522 28424 9528 28436
rect 9580 28424 9586 28476
rect 1886 28396 1892 28408
rect 1847 28368 1892 28396
rect 1886 28356 1892 28368
rect 1944 28356 1950 28408
rect 2070 28356 2076 28408
rect 2128 28396 2134 28408
rect 2165 28399 2223 28405
rect 2165 28396 2177 28399
rect 2128 28368 2177 28396
rect 2128 28356 2134 28368
rect 2165 28365 2177 28368
rect 2211 28365 2223 28399
rect 2165 28359 2223 28365
rect 2254 28356 2260 28408
rect 2312 28396 2318 28408
rect 2809 28399 2867 28405
rect 2809 28396 2821 28399
rect 2312 28368 2821 28396
rect 2312 28356 2318 28368
rect 2809 28365 2821 28368
rect 2855 28396 2867 28399
rect 3174 28396 3180 28408
rect 2855 28368 3180 28396
rect 2855 28365 2867 28368
rect 2809 28359 2867 28365
rect 3174 28356 3180 28368
rect 3232 28396 3238 28408
rect 3545 28399 3603 28405
rect 3545 28396 3557 28399
rect 3232 28368 3557 28396
rect 3232 28356 3238 28368
rect 3545 28365 3557 28368
rect 3591 28365 3603 28399
rect 3545 28359 3603 28365
rect 3560 28328 3588 28359
rect 4186 28356 4192 28408
rect 4244 28396 4250 28408
rect 4465 28399 4523 28405
rect 4465 28396 4477 28399
rect 4244 28368 4477 28396
rect 4244 28356 4250 28368
rect 4465 28365 4477 28368
rect 4511 28365 4523 28399
rect 4465 28359 4523 28365
rect 4649 28399 4707 28405
rect 4649 28365 4661 28399
rect 4695 28365 4707 28399
rect 5014 28396 5020 28408
rect 4975 28368 5020 28396
rect 4649 28359 4707 28365
rect 4664 28328 4692 28359
rect 5014 28356 5020 28368
rect 5072 28356 5078 28408
rect 5658 28356 5664 28408
rect 5716 28396 5722 28408
rect 6305 28399 6363 28405
rect 6305 28396 6317 28399
rect 5716 28368 6317 28396
rect 5716 28356 5722 28368
rect 6305 28365 6317 28368
rect 6351 28396 6363 28399
rect 6946 28396 6952 28408
rect 6351 28368 6952 28396
rect 6351 28365 6363 28368
rect 6305 28359 6363 28365
rect 6946 28356 6952 28368
rect 7004 28396 7010 28408
rect 7041 28399 7099 28405
rect 7041 28396 7053 28399
rect 7004 28368 7053 28396
rect 7004 28356 7010 28368
rect 7041 28365 7053 28368
rect 7087 28365 7099 28399
rect 7590 28396 7596 28408
rect 7503 28368 7596 28396
rect 7041 28359 7099 28365
rect 7590 28356 7596 28368
rect 7648 28396 7654 28408
rect 8421 28399 8479 28405
rect 8421 28396 8433 28399
rect 7648 28368 8433 28396
rect 7648 28356 7654 28368
rect 8421 28365 8433 28368
rect 8467 28365 8479 28399
rect 9062 28396 9068 28408
rect 9023 28368 9068 28396
rect 8421 28359 8479 28365
rect 9062 28356 9068 28368
rect 9120 28396 9126 28408
rect 9893 28399 9951 28405
rect 9893 28396 9905 28399
rect 9120 28368 9905 28396
rect 9120 28356 9126 28368
rect 9893 28365 9905 28368
rect 9939 28396 9951 28399
rect 10077 28399 10135 28405
rect 10077 28396 10089 28399
rect 9939 28368 10089 28396
rect 9939 28365 9951 28368
rect 9893 28359 9951 28365
rect 10077 28365 10089 28368
rect 10123 28396 10135 28399
rect 10442 28396 10448 28408
rect 10123 28368 10448 28396
rect 10123 28365 10135 28368
rect 10077 28359 10135 28365
rect 10442 28356 10448 28368
rect 10500 28356 10506 28408
rect 12852 28396 12880 28563
rect 13294 28560 13300 28572
rect 13352 28560 13358 28612
rect 13662 28600 13668 28612
rect 13623 28572 13668 28600
rect 13662 28560 13668 28572
rect 13720 28560 13726 28612
rect 14582 28560 14588 28612
rect 14640 28600 14646 28612
rect 14953 28603 15011 28609
rect 14953 28600 14965 28603
rect 14640 28572 14965 28600
rect 14640 28560 14646 28572
rect 14953 28569 14965 28572
rect 14999 28569 15011 28603
rect 15410 28600 15416 28612
rect 15371 28572 15416 28600
rect 14953 28563 15011 28569
rect 15410 28560 15416 28572
rect 15468 28560 15474 28612
rect 16974 28600 16980 28612
rect 16935 28572 16980 28600
rect 16974 28560 16980 28572
rect 17032 28600 17038 28612
rect 17713 28603 17771 28609
rect 17713 28600 17725 28603
rect 17032 28572 17725 28600
rect 17032 28560 17038 28572
rect 17713 28569 17725 28572
rect 17759 28569 17771 28603
rect 17713 28563 17771 28569
rect 13312 28532 13340 28560
rect 13941 28535 13999 28541
rect 13941 28532 13953 28535
rect 13312 28504 13953 28532
rect 13941 28501 13953 28504
rect 13987 28501 13999 28535
rect 17158 28532 17164 28544
rect 17119 28504 17164 28532
rect 13941 28495 13999 28501
rect 17158 28492 17164 28504
rect 17216 28492 17222 28544
rect 17618 28532 17624 28544
rect 17579 28504 17624 28532
rect 17618 28492 17624 28504
rect 17676 28492 17682 28544
rect 13202 28464 13208 28476
rect 13163 28436 13208 28464
rect 13202 28424 13208 28436
rect 13260 28464 13266 28476
rect 13757 28467 13815 28473
rect 13757 28464 13769 28467
rect 13260 28436 13769 28464
rect 13260 28424 13266 28436
rect 13757 28433 13769 28436
rect 13803 28433 13815 28467
rect 13757 28427 13815 28433
rect 14493 28467 14551 28473
rect 14493 28433 14505 28467
rect 14539 28464 14551 28467
rect 16146 28464 16152 28476
rect 14539 28436 16152 28464
rect 14539 28433 14551 28436
rect 14493 28427 14551 28433
rect 16146 28424 16152 28436
rect 16204 28424 16210 28476
rect 17437 28467 17495 28473
rect 17437 28433 17449 28467
rect 17483 28464 17495 28467
rect 17526 28464 17532 28476
rect 17483 28436 17532 28464
rect 17483 28433 17495 28436
rect 17437 28427 17495 28433
rect 17526 28424 17532 28436
rect 17584 28424 17590 28476
rect 17728 28464 17756 28563
rect 23506 28560 23512 28612
rect 23564 28600 23570 28612
rect 23693 28603 23751 28609
rect 23693 28600 23705 28603
rect 23564 28572 23705 28600
rect 23564 28560 23570 28572
rect 23693 28569 23705 28572
rect 23739 28569 23751 28603
rect 24518 28600 24524 28612
rect 24479 28572 24524 28600
rect 23693 28563 23751 28569
rect 24518 28560 24524 28572
rect 24576 28600 24582 28612
rect 27186 28600 27192 28612
rect 24576 28572 25116 28600
rect 27147 28572 27192 28600
rect 24576 28560 24582 28572
rect 23969 28535 24027 28541
rect 23969 28501 23981 28535
rect 24015 28532 24027 28535
rect 24610 28532 24616 28544
rect 24015 28504 24616 28532
rect 24015 28501 24027 28504
rect 23969 28495 24027 28501
rect 24610 28492 24616 28504
rect 24668 28492 24674 28544
rect 18357 28467 18415 28473
rect 18357 28464 18369 28467
rect 17728 28436 18369 28464
rect 18357 28433 18369 28436
rect 18403 28433 18415 28467
rect 18357 28427 18415 28433
rect 18722 28424 18728 28476
rect 18780 28464 18786 28476
rect 20105 28467 20163 28473
rect 20105 28464 20117 28467
rect 18780 28436 20117 28464
rect 18780 28424 18786 28436
rect 20105 28433 20117 28436
rect 20151 28433 20163 28467
rect 21850 28464 21856 28476
rect 21763 28436 21856 28464
rect 20105 28427 20163 28433
rect 21850 28424 21856 28436
rect 21908 28464 21914 28476
rect 23046 28464 23052 28476
rect 21908 28436 22448 28464
rect 21908 28424 21914 28436
rect 13021 28399 13079 28405
rect 13021 28396 13033 28399
rect 12852 28368 13033 28396
rect 13021 28365 13033 28368
rect 13067 28365 13079 28399
rect 13021 28359 13079 28365
rect 13110 28356 13116 28408
rect 13168 28396 13174 28408
rect 14769 28399 14827 28405
rect 14769 28396 14781 28399
rect 13168 28368 14781 28396
rect 13168 28356 13174 28368
rect 14769 28365 14781 28368
rect 14815 28396 14827 28399
rect 15042 28396 15048 28408
rect 14815 28368 15048 28396
rect 14815 28365 14827 28368
rect 14769 28359 14827 28365
rect 15042 28356 15048 28368
rect 15100 28356 15106 28408
rect 15781 28399 15839 28405
rect 15781 28365 15793 28399
rect 15827 28396 15839 28399
rect 15827 28368 16560 28396
rect 15827 28365 15839 28368
rect 15781 28359 15839 28365
rect 6121 28331 6179 28337
rect 6121 28328 6133 28331
rect 3560 28300 4692 28328
rect 5860 28300 6133 28328
rect 1334 28260 1340 28272
rect 1295 28232 1340 28260
rect 1334 28220 1340 28232
rect 1392 28220 1398 28272
rect 3450 28260 3456 28272
rect 3411 28232 3456 28260
rect 3450 28220 3456 28232
rect 3508 28220 3514 28272
rect 3913 28263 3971 28269
rect 3913 28229 3925 28263
rect 3959 28260 3971 28263
rect 4186 28260 4192 28272
rect 3959 28232 4192 28260
rect 3959 28229 3971 28232
rect 3913 28223 3971 28229
rect 4186 28220 4192 28232
rect 4244 28220 4250 28272
rect 5750 28220 5756 28272
rect 5808 28260 5814 28272
rect 5860 28269 5888 28300
rect 6121 28297 6133 28300
rect 6167 28297 6179 28331
rect 6121 28291 6179 28297
rect 9430 28288 9436 28340
rect 9488 28328 9494 28340
rect 10261 28331 10319 28337
rect 10261 28328 10273 28331
rect 9488 28300 10273 28328
rect 9488 28288 9494 28300
rect 10261 28297 10273 28300
rect 10307 28328 10319 28331
rect 11089 28331 11147 28337
rect 11089 28328 11101 28331
rect 10307 28300 11101 28328
rect 10307 28297 10319 28300
rect 10261 28291 10319 28297
rect 11089 28297 11101 28300
rect 11135 28297 11147 28331
rect 11089 28291 11147 28297
rect 15410 28288 15416 28340
rect 15468 28328 15474 28340
rect 15597 28331 15655 28337
rect 15597 28328 15609 28331
rect 15468 28300 15609 28328
rect 15468 28288 15474 28300
rect 15597 28297 15609 28300
rect 15643 28328 15655 28331
rect 15962 28328 15968 28340
rect 15643 28300 15968 28328
rect 15643 28297 15655 28300
rect 15597 28291 15655 28297
rect 15962 28288 15968 28300
rect 16020 28328 16026 28340
rect 16425 28331 16483 28337
rect 16425 28328 16437 28331
rect 16020 28300 16437 28328
rect 16020 28288 16026 28300
rect 16425 28297 16437 28300
rect 16471 28297 16483 28331
rect 16425 28291 16483 28297
rect 5845 28263 5903 28269
rect 5845 28260 5857 28263
rect 5808 28232 5857 28260
rect 5808 28220 5814 28232
rect 5845 28229 5857 28232
rect 5891 28229 5903 28263
rect 7682 28260 7688 28272
rect 7643 28232 7688 28260
rect 5845 28223 5903 28229
rect 7682 28220 7688 28232
rect 7740 28220 7746 28272
rect 10534 28260 10540 28272
rect 10495 28232 10540 28260
rect 10534 28220 10540 28232
rect 10592 28220 10598 28272
rect 10994 28260 11000 28272
rect 10955 28232 11000 28260
rect 10994 28220 11000 28232
rect 11052 28220 11058 28272
rect 11270 28220 11276 28272
rect 11328 28260 11334 28272
rect 11825 28263 11883 28269
rect 11825 28260 11837 28263
rect 11328 28232 11837 28260
rect 11328 28220 11334 28232
rect 11825 28229 11837 28232
rect 11871 28260 11883 28263
rect 11914 28260 11920 28272
rect 11871 28232 11920 28260
rect 11871 28229 11883 28232
rect 11825 28223 11883 28229
rect 11914 28220 11920 28232
rect 11972 28220 11978 28272
rect 14674 28260 14680 28272
rect 14635 28232 14680 28260
rect 14674 28220 14680 28232
rect 14732 28220 14738 28272
rect 15226 28260 15232 28272
rect 15187 28232 15232 28260
rect 15226 28220 15232 28232
rect 15284 28220 15290 28272
rect 16333 28263 16391 28269
rect 16333 28229 16345 28263
rect 16379 28260 16391 28263
rect 16532 28260 16560 28368
rect 17342 28356 17348 28408
rect 17400 28396 17406 28408
rect 18078 28396 18084 28408
rect 17400 28368 18084 28396
rect 17400 28356 17406 28368
rect 18078 28356 18084 28368
rect 18136 28356 18142 28408
rect 22420 28405 22448 28436
rect 22972 28436 23052 28464
rect 22972 28405 23000 28436
rect 23046 28424 23052 28436
rect 23104 28424 23110 28476
rect 25088 28473 25116 28572
rect 27186 28560 27192 28572
rect 27244 28560 27250 28612
rect 27557 28603 27615 28609
rect 27557 28569 27569 28603
rect 27603 28600 27615 28603
rect 27646 28600 27652 28612
rect 27603 28572 27652 28600
rect 27603 28569 27615 28572
rect 27557 28563 27615 28569
rect 27646 28560 27652 28572
rect 27704 28560 27710 28612
rect 28198 28600 28204 28612
rect 28159 28572 28204 28600
rect 28198 28560 28204 28572
rect 28256 28600 28262 28612
rect 29946 28600 29952 28612
rect 28256 28572 28796 28600
rect 29907 28572 29952 28600
rect 28256 28560 28262 28572
rect 26910 28492 26916 28544
rect 26968 28532 26974 28544
rect 27281 28535 27339 28541
rect 27281 28532 27293 28535
rect 26968 28504 27293 28532
rect 26968 28492 26974 28504
rect 27281 28501 27293 28504
rect 27327 28501 27339 28535
rect 27281 28495 27339 28501
rect 25073 28467 25131 28473
rect 25073 28433 25085 28467
rect 25119 28433 25131 28467
rect 25073 28427 25131 28433
rect 25901 28467 25959 28473
rect 25901 28433 25913 28467
rect 25947 28464 25959 28467
rect 26174 28464 26180 28476
rect 25947 28436 26180 28464
rect 25947 28433 25959 28436
rect 25901 28427 25959 28433
rect 26174 28424 26180 28436
rect 26232 28464 26238 28476
rect 28106 28464 28112 28476
rect 26232 28436 28112 28464
rect 26232 28424 26238 28436
rect 28106 28424 28112 28436
rect 28164 28424 28170 28476
rect 28768 28473 28796 28572
rect 29946 28560 29952 28572
rect 30004 28560 30010 28612
rect 28753 28467 28811 28473
rect 28753 28433 28765 28467
rect 28799 28433 28811 28467
rect 28753 28427 28811 28433
rect 21577 28399 21635 28405
rect 21577 28365 21589 28399
rect 21623 28396 21635 28399
rect 22405 28399 22463 28405
rect 21623 28368 22264 28396
rect 21623 28365 21635 28368
rect 21577 28359 21635 28365
rect 19366 28288 19372 28340
rect 19424 28288 19430 28340
rect 20102 28288 20108 28340
rect 20160 28328 20166 28340
rect 22236 28337 22264 28368
rect 22405 28365 22417 28399
rect 22451 28396 22463 28399
rect 22773 28399 22831 28405
rect 22773 28396 22785 28399
rect 22451 28368 22785 28396
rect 22451 28365 22463 28368
rect 22405 28359 22463 28365
rect 22773 28365 22785 28368
rect 22819 28396 22831 28399
rect 22957 28399 23015 28405
rect 22957 28396 22969 28399
rect 22819 28368 22969 28396
rect 22819 28365 22831 28368
rect 22773 28359 22831 28365
rect 22957 28365 22969 28368
rect 23003 28365 23015 28399
rect 22957 28359 23015 28365
rect 23690 28356 23696 28408
rect 23748 28396 23754 28408
rect 24978 28396 24984 28408
rect 23748 28368 24840 28396
rect 24939 28368 24984 28396
rect 23748 28356 23754 28368
rect 20381 28331 20439 28337
rect 20381 28328 20393 28331
rect 20160 28300 20393 28328
rect 20160 28288 20166 28300
rect 20381 28297 20393 28300
rect 20427 28297 20439 28331
rect 20381 28291 20439 28297
rect 22221 28331 22279 28337
rect 22221 28297 22233 28331
rect 22267 28328 22279 28331
rect 22494 28328 22500 28340
rect 22267 28300 22500 28328
rect 22267 28297 22279 28300
rect 22221 28291 22279 28297
rect 22494 28288 22500 28300
rect 22552 28288 22558 28340
rect 23046 28288 23052 28340
rect 23104 28328 23110 28340
rect 24812 28337 24840 28368
rect 24978 28356 24984 28368
rect 25036 28356 25042 28408
rect 25809 28399 25867 28405
rect 25809 28365 25821 28399
rect 25855 28365 25867 28399
rect 28014 28396 28020 28408
rect 27927 28368 28020 28396
rect 25809 28359 25867 28365
rect 23233 28331 23291 28337
rect 23233 28328 23245 28331
rect 23104 28300 23245 28328
rect 23104 28288 23110 28300
rect 23233 28297 23245 28300
rect 23279 28328 23291 28331
rect 23509 28331 23567 28337
rect 23509 28328 23521 28331
rect 23279 28300 23521 28328
rect 23279 28297 23291 28300
rect 23233 28291 23291 28297
rect 23509 28297 23521 28300
rect 23555 28297 23567 28331
rect 23509 28291 23567 28297
rect 24797 28331 24855 28337
rect 24797 28297 24809 28331
rect 24843 28328 24855 28331
rect 25824 28328 25852 28359
rect 28014 28356 28020 28368
rect 28072 28396 28078 28408
rect 28661 28399 28719 28405
rect 28661 28396 28673 28399
rect 28072 28368 28673 28396
rect 28072 28356 28078 28368
rect 28661 28365 28673 28368
rect 28707 28365 28719 28399
rect 28661 28359 28719 28365
rect 29489 28399 29547 28405
rect 29489 28365 29501 28399
rect 29535 28365 29547 28399
rect 29489 28359 29547 28365
rect 26082 28328 26088 28340
rect 24843 28300 26088 28328
rect 24843 28297 24855 28300
rect 24797 28291 24855 28297
rect 26082 28288 26088 28300
rect 26140 28288 26146 28340
rect 29504 28328 29532 28359
rect 29578 28356 29584 28408
rect 29636 28396 29642 28408
rect 29636 28368 29681 28396
rect 29636 28356 29642 28368
rect 28492 28300 29532 28328
rect 16606 28260 16612 28272
rect 16379 28232 16612 28260
rect 16379 28229 16391 28232
rect 16333 28223 16391 28229
rect 16606 28220 16612 28232
rect 16664 28220 16670 28272
rect 17986 28260 17992 28272
rect 17947 28232 17992 28260
rect 17986 28220 17992 28232
rect 18044 28220 18050 28272
rect 19384 28260 19412 28288
rect 28492 28272 28520 28300
rect 20197 28263 20255 28269
rect 20197 28260 20209 28263
rect 19384 28232 20209 28260
rect 20197 28229 20209 28232
rect 20243 28260 20255 28263
rect 20286 28260 20292 28272
rect 20243 28232 20292 28260
rect 20243 28229 20255 28232
rect 20197 28223 20255 28229
rect 20286 28220 20292 28232
rect 20344 28220 20350 28272
rect 27005 28263 27063 28269
rect 27005 28229 27017 28263
rect 27051 28260 27063 28263
rect 27278 28260 27284 28272
rect 27051 28232 27284 28260
rect 27051 28229 27063 28232
rect 27005 28223 27063 28229
rect 27278 28220 27284 28232
rect 27336 28220 27342 28272
rect 28385 28263 28443 28269
rect 28385 28229 28397 28263
rect 28431 28260 28443 28263
rect 28474 28260 28480 28272
rect 28431 28232 28480 28260
rect 28431 28229 28443 28232
rect 28385 28223 28443 28229
rect 28474 28220 28480 28232
rect 28532 28220 28538 28272
rect 29026 28220 29032 28272
rect 29084 28260 29090 28272
rect 29762 28260 29768 28272
rect 29084 28232 29768 28260
rect 29084 28220 29090 28232
rect 29762 28220 29768 28232
rect 29820 28220 29826 28272
rect 400 28170 31680 28192
rect 400 28118 18870 28170
rect 18922 28118 18934 28170
rect 18986 28118 18998 28170
rect 19050 28118 19062 28170
rect 19114 28118 19126 28170
rect 19178 28118 31680 28170
rect 400 28096 31680 28118
rect 2717 28059 2775 28065
rect 2717 28025 2729 28059
rect 2763 28056 2775 28059
rect 3082 28056 3088 28068
rect 2763 28028 3088 28056
rect 2763 28025 2775 28028
rect 2717 28019 2775 28025
rect 3082 28016 3088 28028
rect 3140 28056 3146 28068
rect 3358 28056 3364 28068
rect 3140 28028 3364 28056
rect 3140 28016 3146 28028
rect 3358 28016 3364 28028
rect 3416 28016 3422 28068
rect 4278 28056 4284 28068
rect 4239 28028 4284 28056
rect 4278 28016 4284 28028
rect 4336 28056 4342 28068
rect 4465 28059 4523 28065
rect 4465 28056 4477 28059
rect 4336 28028 4477 28056
rect 4336 28016 4342 28028
rect 4465 28025 4477 28028
rect 4511 28025 4523 28059
rect 4465 28019 4523 28025
rect 4741 28059 4799 28065
rect 4741 28025 4753 28059
rect 4787 28056 4799 28059
rect 4922 28056 4928 28068
rect 4787 28028 4928 28056
rect 4787 28025 4799 28028
rect 4741 28019 4799 28025
rect 4922 28016 4928 28028
rect 4980 28056 4986 28068
rect 7682 28056 7688 28068
rect 4980 28028 7688 28056
rect 4980 28016 4986 28028
rect 7682 28016 7688 28028
rect 7740 28016 7746 28068
rect 8145 28059 8203 28065
rect 8145 28025 8157 28059
rect 8191 28056 8203 28059
rect 9062 28056 9068 28068
rect 8191 28028 9068 28056
rect 8191 28025 8203 28028
rect 8145 28019 8203 28025
rect 9062 28016 9068 28028
rect 9120 28016 9126 28068
rect 9246 28056 9252 28068
rect 9207 28028 9252 28056
rect 9246 28016 9252 28028
rect 9304 28016 9310 28068
rect 10353 28059 10411 28065
rect 10353 28025 10365 28059
rect 10399 28056 10411 28059
rect 10534 28056 10540 28068
rect 10399 28028 10540 28056
rect 10399 28025 10411 28028
rect 10353 28019 10411 28025
rect 10534 28016 10540 28028
rect 10592 28016 10598 28068
rect 15873 28059 15931 28065
rect 15873 28025 15885 28059
rect 15919 28056 15931 28059
rect 16146 28056 16152 28068
rect 15919 28028 16152 28056
rect 15919 28025 15931 28028
rect 15873 28019 15931 28025
rect 16146 28016 16152 28028
rect 16204 28016 16210 28068
rect 17986 28016 17992 28068
rect 18044 28056 18050 28068
rect 18722 28056 18728 28068
rect 18044 28028 18728 28056
rect 18044 28016 18050 28028
rect 18722 28016 18728 28028
rect 18780 28056 18786 28068
rect 18909 28059 18967 28065
rect 18909 28056 18921 28059
rect 18780 28028 18921 28056
rect 18780 28016 18786 28028
rect 18909 28025 18921 28028
rect 18955 28025 18967 28059
rect 18909 28019 18967 28025
rect 19185 28059 19243 28065
rect 19185 28025 19197 28059
rect 19231 28056 19243 28059
rect 19274 28056 19280 28068
rect 19231 28028 19280 28056
rect 19231 28025 19243 28028
rect 19185 28019 19243 28025
rect 19274 28016 19280 28028
rect 19332 28016 19338 28068
rect 23046 28056 23052 28068
rect 23007 28028 23052 28056
rect 23046 28016 23052 28028
rect 23104 28016 23110 28068
rect 24978 28056 24984 28068
rect 24939 28028 24984 28056
rect 24978 28016 24984 28028
rect 25036 28016 25042 28068
rect 27830 28056 27836 28068
rect 26376 28028 27836 28056
rect 1334 27948 1340 28000
rect 1392 27988 1398 28000
rect 3913 27991 3971 27997
rect 1392 27960 2116 27988
rect 1392 27948 1398 27960
rect 1889 27923 1947 27929
rect 1889 27889 1901 27923
rect 1935 27920 1947 27923
rect 1978 27920 1984 27932
rect 1935 27892 1984 27920
rect 1935 27889 1947 27892
rect 1889 27883 1947 27889
rect 1978 27880 1984 27892
rect 2036 27880 2042 27932
rect 2088 27929 2116 27960
rect 3913 27957 3925 27991
rect 3959 27988 3971 27991
rect 4094 27988 4100 28000
rect 3959 27960 4100 27988
rect 3959 27957 3971 27960
rect 3913 27951 3971 27957
rect 4094 27948 4100 27960
rect 4152 27948 4158 28000
rect 8786 27948 8792 28000
rect 8844 27988 8850 28000
rect 8844 27960 9476 27988
rect 8844 27948 8850 27960
rect 9448 27932 9476 27960
rect 11270 27948 11276 28000
rect 11328 27948 11334 28000
rect 14950 27948 14956 28000
rect 15008 27988 15014 28000
rect 15137 27991 15195 27997
rect 15137 27988 15149 27991
rect 15008 27960 15149 27988
rect 15008 27948 15014 27960
rect 15137 27957 15149 27960
rect 15183 27988 15195 27991
rect 17526 27988 17532 28000
rect 15183 27960 17532 27988
rect 15183 27957 15195 27960
rect 15137 27951 15195 27957
rect 17526 27948 17532 27960
rect 17584 27948 17590 28000
rect 18173 27991 18231 27997
rect 18173 27957 18185 27991
rect 18219 27988 18231 27991
rect 19366 27988 19372 28000
rect 18219 27960 19372 27988
rect 18219 27957 18231 27960
rect 18173 27951 18231 27957
rect 19366 27948 19372 27960
rect 19424 27948 19430 28000
rect 20565 27991 20623 27997
rect 20565 27957 20577 27991
rect 20611 27988 20623 27991
rect 20930 27988 20936 28000
rect 20611 27960 20936 27988
rect 20611 27957 20623 27960
rect 20565 27951 20623 27957
rect 20930 27948 20936 27960
rect 20988 27988 20994 28000
rect 24610 27988 24616 28000
rect 20988 27960 22540 27988
rect 24523 27960 24616 27988
rect 20988 27948 20994 27960
rect 22512 27932 22540 27960
rect 24610 27948 24616 27960
rect 24668 27988 24674 28000
rect 26376 27988 26404 28028
rect 27830 28016 27836 28028
rect 27888 28016 27894 28068
rect 28661 28059 28719 28065
rect 28661 28025 28673 28059
rect 28707 28056 28719 28059
rect 29578 28056 29584 28068
rect 28707 28028 29584 28056
rect 28707 28025 28719 28028
rect 28661 28019 28719 28025
rect 27186 27988 27192 28000
rect 24668 27960 26404 27988
rect 27147 27960 27192 27988
rect 24668 27948 24674 27960
rect 27186 27948 27192 27960
rect 27244 27948 27250 28000
rect 2073 27923 2131 27929
rect 2073 27889 2085 27923
rect 2119 27920 2131 27923
rect 2162 27920 2168 27932
rect 2119 27892 2168 27920
rect 2119 27889 2131 27892
rect 2073 27883 2131 27889
rect 2162 27880 2168 27892
rect 2220 27880 2226 27932
rect 3358 27920 3364 27932
rect 3319 27892 3364 27920
rect 3358 27880 3364 27892
rect 3416 27880 3422 27932
rect 3450 27880 3456 27932
rect 3508 27920 3514 27932
rect 3545 27923 3603 27929
rect 3545 27920 3557 27923
rect 3508 27892 3557 27920
rect 3508 27880 3514 27892
rect 3545 27889 3557 27892
rect 3591 27920 3603 27923
rect 4002 27920 4008 27932
rect 3591 27892 4008 27920
rect 3591 27889 3603 27892
rect 3545 27883 3603 27889
rect 4002 27880 4008 27892
rect 4060 27880 4066 27932
rect 5658 27920 5664 27932
rect 5619 27892 5664 27920
rect 5658 27880 5664 27892
rect 5716 27880 5722 27932
rect 9249 27923 9307 27929
rect 9249 27889 9261 27923
rect 9295 27920 9307 27923
rect 9338 27920 9344 27932
rect 9295 27892 9344 27920
rect 9295 27889 9307 27892
rect 9249 27883 9307 27889
rect 9338 27880 9344 27892
rect 9396 27880 9402 27932
rect 9430 27880 9436 27932
rect 9488 27920 9494 27932
rect 9488 27892 9581 27920
rect 9488 27880 9494 27892
rect 10350 27880 10356 27932
rect 10408 27920 10414 27932
rect 10537 27923 10595 27929
rect 10537 27920 10549 27923
rect 10408 27892 10549 27920
rect 10408 27880 10414 27892
rect 10537 27889 10549 27892
rect 10583 27889 10595 27923
rect 10537 27883 10595 27889
rect 15321 27923 15379 27929
rect 15321 27889 15333 27923
rect 15367 27920 15379 27923
rect 15962 27920 15968 27932
rect 15367 27892 15968 27920
rect 15367 27889 15379 27892
rect 15321 27883 15379 27889
rect 15962 27880 15968 27892
rect 16020 27880 16026 27932
rect 16790 27920 16796 27932
rect 16751 27892 16796 27920
rect 16790 27880 16796 27892
rect 16848 27880 16854 27932
rect 20194 27920 20200 27932
rect 20155 27892 20200 27920
rect 20194 27880 20200 27892
rect 20252 27880 20258 27932
rect 22402 27920 22408 27932
rect 22363 27892 22408 27920
rect 22402 27880 22408 27892
rect 22460 27880 22466 27932
rect 22494 27880 22500 27932
rect 22552 27920 22558 27932
rect 24334 27920 24340 27932
rect 22552 27892 24340 27920
rect 22552 27880 22558 27892
rect 24334 27880 24340 27892
rect 24392 27880 24398 27932
rect 27278 27880 27284 27932
rect 27336 27920 27342 27932
rect 27925 27923 27983 27929
rect 27925 27920 27937 27923
rect 27336 27892 27937 27920
rect 27336 27880 27342 27892
rect 27925 27889 27937 27892
rect 27971 27889 27983 27923
rect 27925 27883 27983 27889
rect 28017 27923 28075 27929
rect 28017 27889 28029 27923
rect 28063 27920 28075 27923
rect 28106 27920 28112 27932
rect 28063 27892 28112 27920
rect 28063 27889 28075 27892
rect 28017 27883 28075 27889
rect 28106 27880 28112 27892
rect 28164 27920 28170 27932
rect 28676 27920 28704 28019
rect 29578 28016 29584 28028
rect 29636 28016 29642 28068
rect 29670 27920 29676 27932
rect 28164 27892 28704 27920
rect 29631 27892 29676 27920
rect 28164 27880 28170 27892
rect 29670 27880 29676 27892
rect 29728 27880 29734 27932
rect 2438 27852 2444 27864
rect 2399 27824 2444 27852
rect 2438 27812 2444 27824
rect 2496 27812 2502 27864
rect 4097 27855 4155 27861
rect 4097 27821 4109 27855
rect 4143 27852 4155 27855
rect 4830 27852 4836 27864
rect 4143 27824 4836 27852
rect 4143 27821 4155 27824
rect 4097 27815 4155 27821
rect 4830 27812 4836 27824
rect 4888 27812 4894 27864
rect 5014 27812 5020 27864
rect 5072 27852 5078 27864
rect 5385 27855 5443 27861
rect 5385 27852 5397 27855
rect 5072 27824 5397 27852
rect 5072 27812 5078 27824
rect 5385 27821 5397 27824
rect 5431 27852 5443 27855
rect 5750 27852 5756 27864
rect 5431 27824 5756 27852
rect 5431 27821 5443 27824
rect 5385 27815 5443 27821
rect 5750 27812 5756 27824
rect 5808 27812 5814 27864
rect 5842 27812 5848 27864
rect 5900 27852 5906 27864
rect 10810 27852 10816 27864
rect 5900 27824 5945 27852
rect 10771 27824 10816 27852
rect 5900 27812 5906 27824
rect 10810 27812 10816 27824
rect 10868 27812 10874 27864
rect 12561 27855 12619 27861
rect 12561 27821 12573 27855
rect 12607 27852 12619 27855
rect 12650 27852 12656 27864
rect 12607 27824 12656 27852
rect 12607 27821 12619 27824
rect 12561 27815 12619 27821
rect 12650 27812 12656 27824
rect 12708 27812 12714 27864
rect 22218 27812 22224 27864
rect 22276 27852 22282 27864
rect 22589 27855 22647 27861
rect 22589 27852 22601 27855
rect 22276 27824 22601 27852
rect 22276 27812 22282 27824
rect 22589 27821 22601 27824
rect 22635 27821 22647 27855
rect 22589 27815 22647 27821
rect 27097 27855 27155 27861
rect 27097 27821 27109 27855
rect 27143 27852 27155 27855
rect 27554 27852 27560 27864
rect 27143 27824 27560 27852
rect 27143 27821 27155 27824
rect 27097 27815 27155 27821
rect 27554 27812 27560 27824
rect 27612 27812 27618 27864
rect 30038 27852 30044 27864
rect 29999 27824 30044 27852
rect 30038 27812 30044 27824
rect 30096 27812 30102 27864
rect 7501 27787 7559 27793
rect 7501 27753 7513 27787
rect 7547 27784 7559 27787
rect 8878 27784 8884 27796
rect 7547 27756 8884 27784
rect 7547 27753 7559 27756
rect 7501 27747 7559 27753
rect 8878 27744 8884 27756
rect 8936 27744 8942 27796
rect 14858 27744 14864 27796
rect 14916 27784 14922 27796
rect 23506 27784 23512 27796
rect 14916 27756 23512 27784
rect 14916 27744 14922 27756
rect 23506 27744 23512 27756
rect 23564 27744 23570 27796
rect 7317 27719 7375 27725
rect 7317 27685 7329 27719
rect 7363 27716 7375 27719
rect 7866 27716 7872 27728
rect 7363 27688 7872 27716
rect 7363 27685 7375 27688
rect 7317 27679 7375 27685
rect 7866 27676 7872 27688
rect 7924 27676 7930 27728
rect 15410 27716 15416 27728
rect 15371 27688 15416 27716
rect 15410 27676 15416 27688
rect 15468 27676 15474 27728
rect 16606 27716 16612 27728
rect 16567 27688 16612 27716
rect 16606 27676 16612 27688
rect 16664 27676 16670 27728
rect 400 27626 31680 27648
rect 400 27574 3510 27626
rect 3562 27574 3574 27626
rect 3626 27574 3638 27626
rect 3690 27574 3702 27626
rect 3754 27574 3766 27626
rect 3818 27574 31680 27626
rect 400 27552 31680 27574
rect 2162 27512 2168 27524
rect 2123 27484 2168 27512
rect 2162 27472 2168 27484
rect 2220 27472 2226 27524
rect 3913 27515 3971 27521
rect 3913 27481 3925 27515
rect 3959 27512 3971 27515
rect 4094 27512 4100 27524
rect 3959 27484 4100 27512
rect 3959 27481 3971 27484
rect 3913 27475 3971 27481
rect 4094 27472 4100 27484
rect 4152 27472 4158 27524
rect 4830 27472 4836 27524
rect 4888 27512 4894 27524
rect 5385 27515 5443 27521
rect 5385 27512 5397 27515
rect 4888 27484 5397 27512
rect 4888 27472 4894 27484
rect 5385 27481 5397 27484
rect 5431 27481 5443 27515
rect 5385 27475 5443 27481
rect 6026 27472 6032 27524
rect 6084 27512 6090 27524
rect 6949 27515 7007 27521
rect 6949 27512 6961 27515
rect 6084 27484 6961 27512
rect 6084 27472 6090 27484
rect 6949 27481 6961 27484
rect 6995 27512 7007 27515
rect 9430 27512 9436 27524
rect 6995 27484 8004 27512
rect 9391 27484 9436 27512
rect 6995 27481 7007 27484
rect 6949 27475 7007 27481
rect 2349 27447 2407 27453
rect 2349 27413 2361 27447
rect 2395 27444 2407 27447
rect 2438 27444 2444 27456
rect 2395 27416 2444 27444
rect 2395 27413 2407 27416
rect 2349 27407 2407 27413
rect 2438 27404 2444 27416
rect 2496 27444 2502 27456
rect 3266 27444 3272 27456
rect 2496 27416 3272 27444
rect 2496 27404 2502 27416
rect 3266 27404 3272 27416
rect 3324 27444 3330 27456
rect 5014 27444 5020 27456
rect 3324 27416 5020 27444
rect 3324 27404 3330 27416
rect 5014 27404 5020 27416
rect 5072 27404 5078 27456
rect 5293 27447 5351 27453
rect 5293 27413 5305 27447
rect 5339 27444 5351 27447
rect 5658 27444 5664 27456
rect 5339 27416 5664 27444
rect 5339 27413 5351 27416
rect 5293 27407 5351 27413
rect 5658 27404 5664 27416
rect 5716 27404 5722 27456
rect 6854 27404 6860 27456
rect 6912 27444 6918 27456
rect 7041 27447 7099 27453
rect 7041 27444 7053 27447
rect 6912 27416 7053 27444
rect 6912 27404 6918 27416
rect 7041 27413 7053 27416
rect 7087 27444 7099 27447
rect 7225 27447 7283 27453
rect 7225 27444 7237 27447
rect 7087 27416 7237 27444
rect 7087 27413 7099 27416
rect 7041 27407 7099 27413
rect 7225 27413 7237 27416
rect 7271 27413 7283 27447
rect 7590 27444 7596 27456
rect 7551 27416 7596 27444
rect 7225 27407 7283 27413
rect 7590 27404 7596 27416
rect 7648 27404 7654 27456
rect 1337 27379 1395 27385
rect 1337 27345 1349 27379
rect 1383 27376 1395 27379
rect 1426 27376 1432 27388
rect 1383 27348 1432 27376
rect 1383 27345 1395 27348
rect 1337 27339 1395 27345
rect 1426 27336 1432 27348
rect 1484 27336 1490 27388
rect 2070 27336 2076 27388
rect 2128 27376 2134 27388
rect 2714 27376 2720 27388
rect 2128 27348 2720 27376
rect 2128 27336 2134 27348
rect 2714 27336 2720 27348
rect 2772 27376 2778 27388
rect 3177 27379 3235 27385
rect 3177 27376 3189 27379
rect 2772 27348 3189 27376
rect 2772 27336 2778 27348
rect 3177 27345 3189 27348
rect 3223 27345 3235 27379
rect 3177 27339 3235 27345
rect 4925 27379 4983 27385
rect 4925 27345 4937 27379
rect 4971 27376 4983 27379
rect 5842 27376 5848 27388
rect 4971 27348 5848 27376
rect 4971 27345 4983 27348
rect 4925 27339 4983 27345
rect 5842 27336 5848 27348
rect 5900 27336 5906 27388
rect 1153 27311 1211 27317
rect 1153 27277 1165 27311
rect 1199 27277 1211 27311
rect 1153 27271 1211 27277
rect 2533 27311 2591 27317
rect 2533 27277 2545 27311
rect 2579 27308 2591 27311
rect 2898 27308 2904 27320
rect 2579 27280 2904 27308
rect 2579 27277 2591 27280
rect 2533 27271 2591 27277
rect 1168 27184 1196 27271
rect 2898 27268 2904 27280
rect 2956 27268 2962 27320
rect 3082 27308 3088 27320
rect 3043 27280 3088 27308
rect 3082 27268 3088 27280
rect 3140 27268 3146 27320
rect 7866 27308 7872 27320
rect 7827 27280 7872 27308
rect 7866 27268 7872 27280
rect 7924 27268 7930 27320
rect 7976 27317 8004 27484
rect 9430 27472 9436 27484
rect 9488 27472 9494 27524
rect 10350 27512 10356 27524
rect 10311 27484 10356 27512
rect 10350 27472 10356 27484
rect 10408 27472 10414 27524
rect 10810 27512 10816 27524
rect 10771 27484 10816 27512
rect 10810 27472 10816 27484
rect 10868 27472 10874 27524
rect 10997 27515 11055 27521
rect 10997 27481 11009 27515
rect 11043 27512 11055 27515
rect 11270 27512 11276 27524
rect 11043 27484 11276 27512
rect 11043 27481 11055 27484
rect 10997 27475 11055 27481
rect 11270 27472 11276 27484
rect 11328 27472 11334 27524
rect 14769 27515 14827 27521
rect 14769 27481 14781 27515
rect 14815 27512 14827 27515
rect 15410 27512 15416 27524
rect 14815 27484 15416 27512
rect 14815 27481 14827 27484
rect 14769 27475 14827 27481
rect 15410 27472 15416 27484
rect 15468 27472 15474 27524
rect 15962 27512 15968 27524
rect 15875 27484 15968 27512
rect 15962 27472 15968 27484
rect 16020 27512 16026 27524
rect 16422 27512 16428 27524
rect 16020 27484 16428 27512
rect 16020 27472 16026 27484
rect 16422 27472 16428 27484
rect 16480 27512 16486 27524
rect 17158 27512 17164 27524
rect 16480 27484 17164 27512
rect 16480 27472 16486 27484
rect 17158 27472 17164 27484
rect 17216 27472 17222 27524
rect 20930 27512 20936 27524
rect 20891 27484 20936 27512
rect 20930 27472 20936 27484
rect 20988 27472 20994 27524
rect 24334 27472 24340 27524
rect 24392 27512 24398 27524
rect 25073 27515 25131 27521
rect 25073 27512 25085 27515
rect 24392 27484 25085 27512
rect 24392 27472 24398 27484
rect 25073 27481 25085 27484
rect 25119 27481 25131 27515
rect 27186 27512 27192 27524
rect 27147 27484 27192 27512
rect 25073 27475 25131 27481
rect 27186 27472 27192 27484
rect 27244 27472 27250 27524
rect 27554 27512 27560 27524
rect 27515 27484 27560 27512
rect 27554 27472 27560 27484
rect 27612 27472 27618 27524
rect 29949 27515 30007 27521
rect 29949 27481 29961 27515
rect 29995 27512 30007 27515
rect 30038 27512 30044 27524
rect 29995 27484 30044 27512
rect 29995 27481 30007 27484
rect 29949 27475 30007 27481
rect 30038 27472 30044 27484
rect 30096 27472 30102 27524
rect 14950 27444 14956 27456
rect 14911 27416 14956 27444
rect 14950 27404 14956 27416
rect 15008 27404 15014 27456
rect 15042 27404 15048 27456
rect 15100 27444 15106 27456
rect 15505 27447 15563 27453
rect 15505 27444 15517 27447
rect 15100 27416 15517 27444
rect 15100 27404 15106 27416
rect 9338 27376 9344 27388
rect 9251 27348 9344 27376
rect 9338 27336 9344 27348
rect 9396 27376 9402 27388
rect 10626 27376 10632 27388
rect 9396 27348 10632 27376
rect 9396 27336 9402 27348
rect 10626 27336 10632 27348
rect 10684 27376 10690 27388
rect 11365 27379 11423 27385
rect 11365 27376 11377 27379
rect 10684 27348 11377 27376
rect 10684 27336 10690 27348
rect 11365 27345 11377 27348
rect 11411 27376 11423 27379
rect 12650 27376 12656 27388
rect 11411 27348 12656 27376
rect 11411 27345 11423 27348
rect 11365 27339 11423 27345
rect 12650 27336 12656 27348
rect 12708 27336 12714 27388
rect 7961 27311 8019 27317
rect 7961 27277 7973 27311
rect 8007 27277 8019 27311
rect 8694 27308 8700 27320
rect 8655 27280 8700 27308
rect 7961 27271 8019 27277
rect 8694 27268 8700 27280
rect 8752 27268 8758 27320
rect 8878 27308 8884 27320
rect 8839 27280 8884 27308
rect 8878 27268 8884 27280
rect 8936 27268 8942 27320
rect 9246 27268 9252 27320
rect 9304 27308 9310 27320
rect 9617 27311 9675 27317
rect 9617 27308 9629 27311
rect 9304 27280 9629 27308
rect 9304 27268 9310 27280
rect 9617 27277 9629 27280
rect 9663 27277 9675 27311
rect 9617 27271 9675 27277
rect 10994 27268 11000 27320
rect 11052 27308 11058 27320
rect 11549 27311 11607 27317
rect 11549 27308 11561 27311
rect 11052 27280 11561 27308
rect 11052 27268 11058 27280
rect 11549 27277 11561 27280
rect 11595 27308 11607 27311
rect 12193 27311 12251 27317
rect 12193 27308 12205 27311
rect 11595 27280 12205 27308
rect 11595 27277 11607 27280
rect 11549 27271 11607 27277
rect 12193 27277 12205 27280
rect 12239 27277 12251 27311
rect 12558 27308 12564 27320
rect 12519 27280 12564 27308
rect 12193 27271 12251 27277
rect 12558 27268 12564 27280
rect 12616 27268 12622 27320
rect 15152 27317 15180 27416
rect 15505 27413 15517 27416
rect 15551 27413 15563 27447
rect 15505 27407 15563 27413
rect 16609 27447 16667 27453
rect 16609 27413 16621 27447
rect 16655 27444 16667 27447
rect 16790 27444 16796 27456
rect 16655 27416 16796 27444
rect 16655 27413 16667 27416
rect 16609 27407 16667 27413
rect 16790 27404 16796 27416
rect 16848 27404 16854 27456
rect 27465 27447 27523 27453
rect 27465 27413 27477 27447
rect 27511 27444 27523 27447
rect 28106 27444 28112 27456
rect 27511 27416 28112 27444
rect 27511 27413 27523 27416
rect 27465 27407 27523 27413
rect 28106 27404 28112 27416
rect 28164 27404 28170 27456
rect 16882 27336 16888 27388
rect 16940 27376 16946 27388
rect 20194 27376 20200 27388
rect 16940 27348 20200 27376
rect 16940 27336 16946 27348
rect 20194 27336 20200 27348
rect 20252 27376 20258 27388
rect 20473 27379 20531 27385
rect 20473 27376 20485 27379
rect 20252 27348 20485 27376
rect 20252 27336 20258 27348
rect 20473 27345 20485 27348
rect 20519 27345 20531 27379
rect 22954 27376 22960 27388
rect 22915 27348 22960 27376
rect 20473 27339 20531 27345
rect 22954 27336 22960 27348
rect 23012 27336 23018 27388
rect 15137 27311 15195 27317
rect 15137 27277 15149 27311
rect 15183 27277 15195 27311
rect 15137 27271 15195 27277
rect 19921 27311 19979 27317
rect 19921 27277 19933 27311
rect 19967 27308 19979 27311
rect 21114 27308 21120 27320
rect 19967 27280 21120 27308
rect 19967 27277 19979 27280
rect 19921 27271 19979 27277
rect 1978 27240 1984 27252
rect 1891 27212 1984 27240
rect 1978 27200 1984 27212
rect 2036 27240 2042 27252
rect 3266 27240 3272 27252
rect 2036 27212 3272 27240
rect 2036 27200 2042 27212
rect 3266 27200 3272 27212
rect 3324 27200 3330 27252
rect 3358 27200 3364 27252
rect 3416 27240 3422 27252
rect 3637 27243 3695 27249
rect 3637 27240 3649 27243
rect 3416 27212 3649 27240
rect 3416 27200 3422 27212
rect 3637 27209 3649 27212
rect 3683 27209 3695 27243
rect 3637 27203 3695 27209
rect 6765 27243 6823 27249
rect 6765 27209 6777 27243
rect 6811 27240 6823 27243
rect 8712 27240 8740 27268
rect 6811 27212 8740 27240
rect 6811 27209 6823 27212
rect 6765 27203 6823 27209
rect 9982 27200 9988 27252
rect 10040 27240 10046 27252
rect 11181 27243 11239 27249
rect 11181 27240 11193 27243
rect 10040 27212 11193 27240
rect 10040 27200 10046 27212
rect 11181 27209 11193 27212
rect 11227 27240 11239 27243
rect 11733 27243 11791 27249
rect 11733 27240 11745 27243
rect 11227 27212 11745 27240
rect 11227 27209 11239 27212
rect 11181 27203 11239 27209
rect 11733 27209 11745 27212
rect 11779 27209 11791 27243
rect 11733 27203 11791 27209
rect 15962 27200 15968 27252
rect 16020 27240 16026 27252
rect 19737 27243 19795 27249
rect 19737 27240 19749 27243
rect 16020 27212 19749 27240
rect 16020 27200 16026 27212
rect 19737 27209 19749 27212
rect 19783 27240 19795 27243
rect 19936 27240 19964 27271
rect 21114 27268 21120 27280
rect 21172 27268 21178 27320
rect 19783 27212 19964 27240
rect 20197 27243 20255 27249
rect 19783 27209 19795 27212
rect 19737 27203 19795 27209
rect 20197 27209 20209 27243
rect 20243 27209 20255 27243
rect 22313 27243 22371 27249
rect 22313 27240 22325 27243
rect 20197 27203 20255 27209
rect 20672 27212 22325 27240
rect 1061 27175 1119 27181
rect 1061 27141 1073 27175
rect 1107 27172 1119 27175
rect 1150 27172 1156 27184
rect 1107 27144 1156 27172
rect 1107 27141 1119 27144
rect 1061 27135 1119 27141
rect 1150 27132 1156 27144
rect 1208 27132 1214 27184
rect 1518 27132 1524 27184
rect 1576 27172 1582 27184
rect 1705 27175 1763 27181
rect 1705 27172 1717 27175
rect 1576 27144 1717 27172
rect 1576 27132 1582 27144
rect 1705 27141 1717 27144
rect 1751 27141 1763 27175
rect 1705 27135 1763 27141
rect 3545 27175 3603 27181
rect 3545 27141 3557 27175
rect 3591 27172 3603 27175
rect 4002 27172 4008 27184
rect 3591 27144 4008 27172
rect 3591 27141 3603 27144
rect 3545 27135 3603 27141
rect 4002 27132 4008 27144
rect 4060 27172 4066 27184
rect 6946 27172 6952 27184
rect 4060 27144 6952 27172
rect 4060 27132 4066 27144
rect 6946 27132 6952 27144
rect 7004 27132 7010 27184
rect 12282 27132 12288 27184
rect 12340 27172 12346 27184
rect 14950 27172 14956 27184
rect 12340 27144 14956 27172
rect 12340 27132 12346 27144
rect 14950 27132 14956 27144
rect 15008 27132 15014 27184
rect 15226 27132 15232 27184
rect 15284 27172 15290 27184
rect 15321 27175 15379 27181
rect 15321 27172 15333 27175
rect 15284 27144 15333 27172
rect 15284 27132 15290 27144
rect 15321 27141 15333 27144
rect 15367 27172 15379 27175
rect 15689 27175 15747 27181
rect 15689 27172 15701 27175
rect 15367 27144 15701 27172
rect 15367 27141 15379 27144
rect 15321 27135 15379 27141
rect 15689 27141 15701 27144
rect 15735 27141 15747 27175
rect 15689 27135 15747 27141
rect 16606 27132 16612 27184
rect 16664 27172 16670 27184
rect 16701 27175 16759 27181
rect 16701 27172 16713 27175
rect 16664 27144 16713 27172
rect 16664 27132 16670 27144
rect 16701 27141 16713 27144
rect 16747 27141 16759 27175
rect 20212 27172 20240 27203
rect 20672 27184 20700 27212
rect 22313 27209 22325 27212
rect 22359 27240 22371 27243
rect 22402 27240 22408 27252
rect 22359 27212 22408 27240
rect 22359 27209 22371 27212
rect 22313 27203 22371 27209
rect 22402 27200 22408 27212
rect 22460 27200 22466 27252
rect 22589 27243 22647 27249
rect 22589 27209 22601 27243
rect 22635 27240 22647 27243
rect 23233 27243 23291 27249
rect 23233 27240 23245 27243
rect 22635 27212 23245 27240
rect 22635 27209 22647 27212
rect 22589 27203 22647 27209
rect 23233 27209 23245 27212
rect 23279 27240 23291 27243
rect 23322 27240 23328 27252
rect 23279 27212 23328 27240
rect 23279 27209 23291 27212
rect 23233 27203 23291 27209
rect 23322 27200 23328 27212
rect 23380 27200 23386 27252
rect 23690 27200 23696 27252
rect 23748 27200 23754 27252
rect 24981 27243 25039 27249
rect 24981 27240 24993 27243
rect 24720 27212 24993 27240
rect 20654 27172 20660 27184
rect 20212 27144 20660 27172
rect 16701 27135 16759 27141
rect 20654 27132 20660 27144
rect 20712 27132 20718 27184
rect 22218 27172 22224 27184
rect 22179 27144 22224 27172
rect 22218 27132 22224 27144
rect 22276 27132 22282 27184
rect 22773 27175 22831 27181
rect 22773 27141 22785 27175
rect 22819 27172 22831 27175
rect 24518 27172 24524 27184
rect 22819 27144 24524 27172
rect 22819 27141 22831 27144
rect 22773 27135 22831 27141
rect 24518 27132 24524 27144
rect 24576 27172 24582 27184
rect 24720 27172 24748 27212
rect 24981 27209 24993 27212
rect 25027 27209 25039 27243
rect 24981 27203 25039 27209
rect 24576 27144 24748 27172
rect 27097 27175 27155 27181
rect 24576 27132 24582 27144
rect 27097 27141 27109 27175
rect 27143 27172 27155 27175
rect 27278 27172 27284 27184
rect 27143 27144 27284 27172
rect 27143 27141 27155 27144
rect 27097 27135 27155 27141
rect 27278 27132 27284 27144
rect 27336 27132 27342 27184
rect 28290 27132 28296 27184
rect 28348 27172 28354 27184
rect 29670 27172 29676 27184
rect 28348 27144 29676 27172
rect 28348 27132 28354 27144
rect 29670 27132 29676 27144
rect 29728 27132 29734 27184
rect 400 27082 31680 27104
rect 400 27030 18870 27082
rect 18922 27030 18934 27082
rect 18986 27030 18998 27082
rect 19050 27030 19062 27082
rect 19114 27030 19126 27082
rect 19178 27030 31680 27082
rect 400 27008 31680 27030
rect 2714 26968 2720 26980
rect 2675 26940 2720 26968
rect 2714 26928 2720 26940
rect 2772 26928 2778 26980
rect 7501 26971 7559 26977
rect 7501 26937 7513 26971
rect 7547 26968 7559 26971
rect 7590 26968 7596 26980
rect 7547 26940 7596 26968
rect 7547 26937 7559 26940
rect 7501 26931 7559 26937
rect 7590 26928 7596 26940
rect 7648 26928 7654 26980
rect 8694 26968 8700 26980
rect 8607 26940 8700 26968
rect 8694 26928 8700 26940
rect 8752 26968 8758 26980
rect 10534 26968 10540 26980
rect 8752 26940 10540 26968
rect 8752 26928 8758 26940
rect 10534 26928 10540 26940
rect 10592 26928 10598 26980
rect 11825 26971 11883 26977
rect 11825 26937 11837 26971
rect 11871 26968 11883 26971
rect 12558 26968 12564 26980
rect 11871 26940 12564 26968
rect 11871 26937 11883 26940
rect 11825 26931 11883 26937
rect 12558 26928 12564 26940
rect 12616 26928 12622 26980
rect 22218 26928 22224 26980
rect 22276 26968 22282 26980
rect 23049 26971 23107 26977
rect 23049 26968 23061 26971
rect 22276 26940 23061 26968
rect 22276 26928 22282 26940
rect 23049 26937 23061 26940
rect 23095 26968 23107 26971
rect 23690 26968 23696 26980
rect 23095 26940 23696 26968
rect 23095 26937 23107 26940
rect 23049 26931 23107 26937
rect 23690 26928 23696 26940
rect 23748 26928 23754 26980
rect 24429 26971 24487 26977
rect 24429 26937 24441 26971
rect 24475 26968 24487 26971
rect 24610 26968 24616 26980
rect 24475 26940 24616 26968
rect 24475 26937 24487 26940
rect 24429 26931 24487 26937
rect 24610 26928 24616 26940
rect 24668 26928 24674 26980
rect 9249 26903 9307 26909
rect 9249 26869 9261 26903
rect 9295 26900 9307 26903
rect 10810 26900 10816 26912
rect 9295 26872 10816 26900
rect 9295 26869 9307 26872
rect 9249 26863 9307 26869
rect 10810 26860 10816 26872
rect 10868 26860 10874 26912
rect 26085 26903 26143 26909
rect 14876 26872 16560 26900
rect 14876 26844 14904 26872
rect 3266 26792 3272 26844
rect 3324 26832 3330 26844
rect 3361 26835 3419 26841
rect 3361 26832 3373 26835
rect 3324 26804 3373 26832
rect 3324 26792 3330 26804
rect 3361 26801 3373 26804
rect 3407 26801 3419 26835
rect 6578 26832 6584 26844
rect 6539 26804 6584 26832
rect 3361 26795 3419 26801
rect 6578 26792 6584 26804
rect 6636 26792 6642 26844
rect 9798 26832 9804 26844
rect 9759 26804 9804 26832
rect 9798 26792 9804 26804
rect 9856 26792 9862 26844
rect 9982 26832 9988 26844
rect 9943 26804 9988 26832
rect 9982 26792 9988 26804
rect 10040 26792 10046 26844
rect 10077 26835 10135 26841
rect 10077 26801 10089 26835
rect 10123 26801 10135 26835
rect 10626 26832 10632 26844
rect 10587 26804 10632 26832
rect 10077 26795 10135 26801
rect 6946 26764 6952 26776
rect 6907 26736 6952 26764
rect 6946 26724 6952 26736
rect 7004 26724 7010 26776
rect 9614 26724 9620 26776
rect 9672 26764 9678 26776
rect 10092 26764 10120 26795
rect 10626 26792 10632 26804
rect 10684 26792 10690 26844
rect 14858 26832 14864 26844
rect 14819 26804 14864 26832
rect 14858 26792 14864 26804
rect 14916 26792 14922 26844
rect 15137 26835 15195 26841
rect 15137 26801 15149 26835
rect 15183 26832 15195 26835
rect 15226 26832 15232 26844
rect 15183 26804 15232 26832
rect 15183 26801 15195 26804
rect 15137 26795 15195 26801
rect 15226 26792 15232 26804
rect 15284 26792 15290 26844
rect 16422 26832 16428 26844
rect 16383 26804 16428 26832
rect 16422 26792 16428 26804
rect 16480 26792 16486 26844
rect 16532 26841 16560 26872
rect 26085 26869 26097 26903
rect 26131 26900 26143 26903
rect 26174 26900 26180 26912
rect 26131 26872 26180 26900
rect 26131 26869 26143 26872
rect 26085 26863 26143 26869
rect 26174 26860 26180 26872
rect 26232 26860 26238 26912
rect 16517 26835 16575 26841
rect 16517 26801 16529 26835
rect 16563 26832 16575 26835
rect 16606 26832 16612 26844
rect 16563 26804 16612 26832
rect 16563 26801 16575 26804
rect 16517 26795 16575 26801
rect 16606 26792 16612 26804
rect 16664 26792 16670 26844
rect 21209 26835 21267 26841
rect 21209 26801 21221 26835
rect 21255 26832 21267 26835
rect 21850 26832 21856 26844
rect 21255 26804 21856 26832
rect 21255 26801 21267 26804
rect 21209 26795 21267 26801
rect 21850 26792 21856 26804
rect 21908 26792 21914 26844
rect 25809 26835 25867 26841
rect 25809 26801 25821 26835
rect 25855 26832 25867 26835
rect 25898 26832 25904 26844
rect 25855 26804 25904 26832
rect 25855 26801 25867 26804
rect 25809 26795 25867 26801
rect 25898 26792 25904 26804
rect 25956 26792 25962 26844
rect 28566 26832 28572 26844
rect 28527 26804 28572 26832
rect 28566 26792 28572 26804
rect 28624 26792 28630 26844
rect 10350 26764 10356 26776
rect 9672 26736 10120 26764
rect 10311 26736 10356 26764
rect 9672 26724 9678 26736
rect 10350 26724 10356 26736
rect 10408 26724 10414 26776
rect 15318 26764 15324 26776
rect 15279 26736 15324 26764
rect 15318 26724 15324 26736
rect 15376 26724 15382 26776
rect 785 26699 843 26705
rect 785 26665 797 26699
rect 831 26696 843 26699
rect 2714 26696 2720 26708
rect 831 26668 2720 26696
rect 831 26665 843 26668
rect 785 26659 843 26665
rect 2714 26656 2720 26668
rect 2772 26656 2778 26708
rect 6854 26696 6860 26708
rect 6815 26668 6860 26696
rect 6854 26656 6860 26668
rect 6912 26656 6918 26708
rect 14953 26699 15011 26705
rect 14953 26665 14965 26699
rect 14999 26696 15011 26699
rect 15134 26696 15140 26708
rect 14999 26668 15140 26696
rect 14999 26665 15011 26668
rect 14953 26659 15011 26665
rect 15134 26656 15140 26668
rect 15192 26696 15198 26708
rect 16440 26696 16468 26792
rect 21390 26764 21396 26776
rect 21351 26736 21396 26764
rect 21390 26724 21396 26736
rect 21448 26724 21454 26776
rect 15192 26668 16468 26696
rect 15192 26656 15198 26668
rect 969 26631 1027 26637
rect 969 26597 981 26631
rect 1015 26628 1027 26631
rect 1426 26628 1432 26640
rect 1015 26600 1432 26628
rect 1015 26597 1027 26600
rect 969 26591 1027 26597
rect 1426 26588 1432 26600
rect 1484 26588 1490 26640
rect 3358 26588 3364 26640
rect 3416 26628 3422 26640
rect 6762 26637 6768 26640
rect 3453 26631 3511 26637
rect 3453 26628 3465 26631
rect 3416 26600 3465 26628
rect 3416 26588 3422 26600
rect 3453 26597 3465 26600
rect 3499 26597 3511 26631
rect 3453 26591 3511 26597
rect 6746 26631 6768 26637
rect 6746 26597 6758 26631
rect 6746 26591 6768 26597
rect 6762 26588 6768 26591
rect 6820 26588 6826 26640
rect 7222 26628 7228 26640
rect 7183 26600 7228 26628
rect 7222 26588 7228 26600
rect 7280 26588 7286 26640
rect 14677 26631 14735 26637
rect 14677 26597 14689 26631
rect 14723 26628 14735 26631
rect 15042 26628 15048 26640
rect 14723 26600 15048 26628
rect 14723 26597 14735 26600
rect 14677 26591 14735 26597
rect 15042 26588 15048 26600
rect 15100 26628 15106 26640
rect 16701 26631 16759 26637
rect 16701 26628 16713 26631
rect 15100 26600 16713 26628
rect 15100 26588 15106 26600
rect 16701 26597 16713 26600
rect 16747 26628 16759 26631
rect 16790 26628 16796 26640
rect 16747 26600 16796 26628
rect 16747 26597 16759 26600
rect 16701 26591 16759 26597
rect 16790 26588 16796 26600
rect 16848 26588 16854 26640
rect 28750 26628 28756 26640
rect 28711 26600 28756 26628
rect 28750 26588 28756 26600
rect 28808 26588 28814 26640
rect 400 26538 31680 26560
rect 400 26486 3510 26538
rect 3562 26486 3574 26538
rect 3626 26486 3638 26538
rect 3690 26486 3702 26538
rect 3754 26486 3766 26538
rect 3818 26486 31680 26538
rect 400 26464 31680 26486
rect 2898 26384 2904 26436
rect 2956 26424 2962 26436
rect 5661 26427 5719 26433
rect 5661 26424 5673 26427
rect 2956 26396 5673 26424
rect 2956 26384 2962 26396
rect 5661 26393 5673 26396
rect 5707 26424 5719 26427
rect 6397 26427 6455 26433
rect 6397 26424 6409 26427
rect 5707 26396 6409 26424
rect 5707 26393 5719 26396
rect 5661 26387 5719 26393
rect 6397 26393 6409 26396
rect 6443 26424 6455 26427
rect 6762 26424 6768 26436
rect 6443 26396 6768 26424
rect 6443 26393 6455 26396
rect 6397 26387 6455 26393
rect 6762 26384 6768 26396
rect 6820 26424 6826 26436
rect 7317 26427 7375 26433
rect 7317 26424 7329 26427
rect 6820 26396 7329 26424
rect 6820 26384 6826 26396
rect 7317 26393 7329 26396
rect 7363 26393 7375 26427
rect 7317 26387 7375 26393
rect 8145 26427 8203 26433
rect 8145 26393 8157 26427
rect 8191 26424 8203 26427
rect 8697 26427 8755 26433
rect 8697 26424 8709 26427
rect 8191 26396 8709 26424
rect 8191 26393 8203 26396
rect 8145 26387 8203 26393
rect 8697 26393 8709 26396
rect 8743 26424 8755 26427
rect 9798 26424 9804 26436
rect 8743 26396 9804 26424
rect 8743 26393 8755 26396
rect 8697 26387 8755 26393
rect 9798 26384 9804 26396
rect 9856 26424 9862 26436
rect 10261 26427 10319 26433
rect 10261 26424 10273 26427
rect 9856 26396 10273 26424
rect 9856 26384 9862 26396
rect 10261 26393 10273 26396
rect 10307 26393 10319 26427
rect 10261 26387 10319 26393
rect 11822 26384 11828 26436
rect 11880 26424 11886 26436
rect 12469 26427 12527 26433
rect 12469 26424 12481 26427
rect 11880 26396 12481 26424
rect 11880 26384 11886 26396
rect 12469 26393 12481 26396
rect 12515 26393 12527 26427
rect 12469 26387 12527 26393
rect 14125 26427 14183 26433
rect 14125 26393 14137 26427
rect 14171 26424 14183 26427
rect 14950 26424 14956 26436
rect 14171 26396 14956 26424
rect 14171 26393 14183 26396
rect 14125 26387 14183 26393
rect 14950 26384 14956 26396
rect 15008 26424 15014 26436
rect 15502 26424 15508 26436
rect 15008 26396 15508 26424
rect 15008 26384 15014 26396
rect 15502 26384 15508 26396
rect 15560 26384 15566 26436
rect 16422 26424 16428 26436
rect 16383 26396 16428 26424
rect 16422 26384 16428 26396
rect 16480 26384 16486 26436
rect 16606 26424 16612 26436
rect 16567 26396 16612 26424
rect 16606 26384 16612 26396
rect 16664 26384 16670 26436
rect 16790 26424 16796 26436
rect 16751 26396 16796 26424
rect 16790 26384 16796 26396
rect 16848 26384 16854 26436
rect 21390 26424 21396 26436
rect 21351 26396 21396 26424
rect 21390 26384 21396 26396
rect 21448 26384 21454 26436
rect 21761 26427 21819 26433
rect 21761 26393 21773 26427
rect 21807 26424 21819 26427
rect 21850 26424 21856 26436
rect 21807 26396 21856 26424
rect 21807 26393 21819 26396
rect 21761 26387 21819 26393
rect 6946 26356 6952 26368
rect 6907 26328 6952 26356
rect 6946 26316 6952 26328
rect 7004 26316 7010 26368
rect 10169 26359 10227 26365
rect 10169 26325 10181 26359
rect 10215 26356 10227 26359
rect 10810 26356 10816 26368
rect 10215 26328 10816 26356
rect 10215 26325 10227 26328
rect 10169 26319 10227 26325
rect 10810 26316 10816 26328
rect 10868 26316 10874 26368
rect 20657 26359 20715 26365
rect 20657 26325 20669 26359
rect 20703 26356 20715 26359
rect 21776 26356 21804 26387
rect 21850 26384 21856 26396
rect 21908 26384 21914 26436
rect 24613 26427 24671 26433
rect 24613 26393 24625 26427
rect 24659 26424 24671 26427
rect 24978 26424 24984 26436
rect 24659 26396 24984 26424
rect 24659 26393 24671 26396
rect 24613 26387 24671 26393
rect 24978 26384 24984 26396
rect 25036 26384 25042 26436
rect 26085 26427 26143 26433
rect 26085 26393 26097 26427
rect 26131 26424 26143 26427
rect 26174 26424 26180 26436
rect 26131 26396 26180 26424
rect 26131 26393 26143 26396
rect 26085 26387 26143 26393
rect 26174 26384 26180 26396
rect 26232 26384 26238 26436
rect 28566 26424 28572 26436
rect 28527 26396 28572 26424
rect 28566 26384 28572 26396
rect 28624 26384 28630 26436
rect 28750 26424 28756 26436
rect 28711 26396 28756 26424
rect 28750 26384 28756 26396
rect 28808 26384 28814 26436
rect 20703 26328 21804 26356
rect 28584 26356 28612 26384
rect 30038 26356 30044 26368
rect 28584 26328 30044 26356
rect 20703 26325 20715 26328
rect 20657 26319 20715 26325
rect 2714 26288 2720 26300
rect 2675 26260 2720 26288
rect 2714 26248 2720 26260
rect 2772 26248 2778 26300
rect 6854 26248 6860 26300
rect 6912 26288 6918 26300
rect 7133 26291 7191 26297
rect 7133 26288 7145 26291
rect 6912 26260 7145 26288
rect 6912 26248 6918 26260
rect 7133 26257 7145 26260
rect 7179 26257 7191 26291
rect 7133 26251 7191 26257
rect 8513 26291 8571 26297
rect 8513 26257 8525 26291
rect 8559 26288 8571 26291
rect 9985 26291 10043 26297
rect 9985 26288 9997 26291
rect 8559 26260 9997 26288
rect 8559 26257 8571 26260
rect 8513 26251 8571 26257
rect 690 26220 696 26232
rect 651 26192 696 26220
rect 690 26180 696 26192
rect 748 26180 754 26232
rect 2732 26220 2760 26248
rect 4281 26223 4339 26229
rect 4281 26220 4293 26223
rect 2732 26192 4293 26220
rect 4281 26189 4293 26192
rect 4327 26220 4339 26223
rect 5937 26223 5995 26229
rect 4327 26192 4554 26220
rect 4327 26189 4339 26192
rect 4281 26183 4339 26189
rect 969 26155 1027 26161
rect 969 26121 981 26155
rect 1015 26121 1027 26155
rect 969 26115 1027 26121
rect 782 26044 788 26096
rect 840 26084 846 26096
rect 984 26084 1012 26115
rect 1426 26112 1432 26164
rect 1484 26112 1490 26164
rect 4526 26152 4554 26192
rect 5937 26189 5949 26223
rect 5983 26220 5995 26223
rect 6118 26220 6124 26232
rect 5983 26192 6124 26220
rect 5983 26189 5995 26192
rect 5937 26183 5995 26189
rect 6118 26180 6124 26192
rect 6176 26180 6182 26232
rect 6213 26223 6271 26229
rect 6213 26189 6225 26223
rect 6259 26220 6271 26223
rect 6765 26223 6823 26229
rect 6765 26220 6777 26223
rect 6259 26192 6777 26220
rect 6259 26189 6271 26192
rect 6213 26183 6271 26189
rect 6765 26189 6777 26192
rect 6811 26189 6823 26223
rect 6765 26183 6823 26189
rect 4833 26155 4891 26161
rect 4833 26152 4845 26155
rect 4526 26124 4845 26152
rect 4833 26121 4845 26124
rect 4879 26152 4891 26155
rect 6228 26152 6256 26183
rect 8694 26180 8700 26232
rect 8752 26220 8758 26232
rect 9246 26220 9252 26232
rect 8752 26192 9252 26220
rect 8752 26180 8758 26192
rect 9246 26180 9252 26192
rect 9304 26180 9310 26232
rect 9632 26229 9660 26260
rect 9985 26257 9997 26260
rect 10031 26288 10043 26291
rect 10626 26288 10632 26300
rect 10031 26260 10632 26288
rect 10031 26257 10043 26260
rect 9985 26251 10043 26257
rect 10626 26248 10632 26260
rect 10684 26248 10690 26300
rect 13941 26291 13999 26297
rect 13941 26257 13953 26291
rect 13987 26288 13999 26291
rect 14309 26291 14367 26297
rect 13987 26260 14214 26288
rect 13987 26257 13999 26260
rect 13941 26251 13999 26257
rect 9341 26223 9399 26229
rect 9341 26189 9353 26223
rect 9387 26189 9399 26223
rect 9341 26183 9399 26189
rect 9617 26223 9675 26229
rect 9617 26189 9629 26223
rect 9663 26189 9675 26223
rect 9617 26183 9675 26189
rect 9801 26223 9859 26229
rect 9801 26189 9813 26223
rect 9847 26220 9859 26223
rect 10534 26220 10540 26232
rect 9847 26192 10540 26220
rect 9847 26189 9859 26192
rect 9801 26183 9859 26189
rect 4879 26124 6256 26152
rect 4879 26121 4891 26124
rect 4833 26115 4891 26121
rect 840 26056 1012 26084
rect 840 26044 846 26056
rect 3266 26044 3272 26096
rect 3324 26084 3330 26096
rect 3361 26087 3419 26093
rect 3361 26084 3373 26087
rect 3324 26056 3373 26084
rect 3324 26044 3330 26056
rect 3361 26053 3373 26056
rect 3407 26053 3419 26087
rect 3361 26047 3419 26053
rect 3450 26044 3456 26096
rect 3508 26084 3514 26096
rect 3545 26087 3603 26093
rect 3545 26084 3557 26087
rect 3508 26056 3557 26084
rect 3508 26044 3514 26056
rect 3545 26053 3557 26056
rect 3591 26053 3603 26087
rect 4554 26084 4560 26096
rect 4515 26056 4560 26084
rect 3545 26047 3603 26053
rect 4554 26044 4560 26056
rect 4612 26084 4618 26096
rect 4925 26087 4983 26093
rect 4925 26084 4937 26087
rect 4612 26056 4937 26084
rect 4612 26044 4618 26056
rect 4925 26053 4937 26056
rect 4971 26053 4983 26087
rect 4925 26047 4983 26053
rect 7866 26044 7872 26096
rect 7924 26084 7930 26096
rect 8234 26084 8240 26096
rect 7924 26056 8240 26084
rect 7924 26044 7930 26056
rect 8234 26044 8240 26056
rect 8292 26084 8298 26096
rect 9356 26084 9384 26183
rect 10534 26180 10540 26192
rect 10592 26180 10598 26232
rect 11733 26223 11791 26229
rect 11733 26189 11745 26223
rect 11779 26220 11791 26223
rect 11822 26220 11828 26232
rect 11779 26192 11828 26220
rect 11779 26189 11791 26192
rect 11733 26183 11791 26189
rect 11822 26180 11828 26192
rect 11880 26180 11886 26232
rect 14186 26220 14214 26260
rect 14309 26257 14321 26291
rect 14355 26288 14367 26291
rect 14674 26288 14680 26300
rect 14355 26260 14680 26288
rect 14355 26257 14367 26260
rect 14309 26251 14367 26257
rect 14674 26248 14680 26260
rect 14732 26288 14738 26300
rect 16422 26288 16428 26300
rect 14732 26260 16428 26288
rect 14732 26248 14738 26260
rect 14861 26223 14919 26229
rect 14861 26220 14873 26223
rect 14186 26192 14873 26220
rect 14861 26189 14873 26192
rect 14907 26189 14919 26223
rect 15042 26220 15048 26232
rect 15003 26192 15048 26220
rect 14861 26183 14919 26189
rect 10718 26112 10724 26164
rect 10776 26152 10782 26164
rect 12009 26155 12067 26161
rect 12009 26152 12021 26155
rect 10776 26124 12021 26152
rect 10776 26112 10782 26124
rect 12009 26121 12021 26124
rect 12055 26152 12067 26155
rect 12285 26155 12343 26161
rect 12285 26152 12297 26155
rect 12055 26124 12297 26152
rect 12055 26121 12067 26124
rect 12009 26115 12067 26121
rect 12285 26121 12297 26124
rect 12331 26121 12343 26155
rect 14876 26152 14904 26183
rect 15042 26180 15048 26192
rect 15100 26180 15106 26232
rect 15428 26229 15456 26260
rect 16422 26248 16428 26260
rect 16480 26248 16486 26300
rect 15413 26223 15471 26229
rect 15413 26189 15425 26223
rect 15459 26189 15471 26223
rect 15413 26183 15471 26189
rect 15502 26180 15508 26232
rect 15560 26220 15566 26232
rect 17713 26223 17771 26229
rect 15560 26192 15605 26220
rect 15560 26180 15566 26192
rect 17713 26189 17725 26223
rect 17759 26220 17771 26223
rect 17802 26220 17808 26232
rect 17759 26192 17808 26220
rect 17759 26189 17771 26192
rect 17713 26183 17771 26189
rect 17802 26180 17808 26192
rect 17860 26220 17866 26232
rect 18449 26223 18507 26229
rect 18449 26220 18461 26223
rect 17860 26192 18461 26220
rect 17860 26180 17866 26192
rect 18449 26189 18461 26192
rect 18495 26220 18507 26223
rect 20102 26220 20108 26232
rect 18495 26192 20108 26220
rect 18495 26189 18507 26192
rect 18449 26183 18507 26189
rect 20102 26180 20108 26192
rect 20160 26180 20166 26232
rect 20194 26180 20200 26232
rect 20252 26220 20258 26232
rect 20764 26229 20792 26328
rect 30038 26316 30044 26328
rect 30096 26316 30102 26368
rect 26913 26291 26971 26297
rect 26913 26257 26925 26291
rect 26959 26288 26971 26291
rect 27557 26291 27615 26297
rect 27557 26288 27569 26291
rect 26959 26260 27569 26288
rect 26959 26257 26971 26260
rect 26913 26251 26971 26257
rect 27557 26257 27569 26260
rect 27603 26288 27615 26291
rect 28014 26288 28020 26300
rect 27603 26260 28020 26288
rect 27603 26257 27615 26260
rect 27557 26251 27615 26257
rect 28014 26248 28020 26260
rect 28072 26248 28078 26300
rect 20749 26223 20807 26229
rect 20749 26220 20761 26223
rect 20252 26192 20761 26220
rect 20252 26180 20258 26192
rect 20749 26189 20761 26192
rect 20795 26189 20807 26223
rect 20749 26183 20807 26189
rect 24889 26223 24947 26229
rect 24889 26189 24901 26223
rect 24935 26220 24947 26223
rect 24935 26192 25668 26220
rect 24935 26189 24947 26192
rect 24889 26183 24947 26189
rect 15226 26152 15232 26164
rect 14876 26124 15232 26152
rect 12285 26115 12343 26121
rect 15226 26112 15232 26124
rect 15284 26152 15290 26164
rect 17989 26155 18047 26161
rect 15284 26124 15824 26152
rect 15284 26112 15290 26124
rect 14674 26084 14680 26096
rect 8292 26056 9384 26084
rect 14635 26056 14680 26084
rect 8292 26044 8298 26056
rect 14674 26044 14680 26056
rect 14732 26044 14738 26096
rect 15796 26093 15824 26124
rect 17989 26121 18001 26155
rect 18035 26121 18047 26155
rect 17989 26115 18047 26121
rect 15781 26087 15839 26093
rect 15781 26053 15793 26087
rect 15827 26084 15839 26087
rect 17710 26084 17716 26096
rect 15827 26056 17716 26084
rect 15827 26053 15839 26056
rect 15781 26047 15839 26053
rect 17710 26044 17716 26056
rect 17768 26044 17774 26096
rect 18004 26084 18032 26115
rect 20930 26112 20936 26164
rect 20988 26152 20994 26164
rect 21025 26155 21083 26161
rect 21025 26152 21037 26155
rect 20988 26124 21037 26152
rect 20988 26112 20994 26124
rect 21025 26121 21037 26124
rect 21071 26152 21083 26155
rect 21485 26155 21543 26161
rect 21485 26152 21497 26155
rect 21071 26124 21497 26152
rect 21071 26121 21083 26124
rect 21025 26115 21083 26121
rect 21485 26121 21497 26124
rect 21531 26121 21543 26155
rect 21485 26115 21543 26121
rect 24242 26112 24248 26164
rect 24300 26152 24306 26164
rect 24705 26155 24763 26161
rect 24705 26152 24717 26155
rect 24300 26124 24717 26152
rect 24300 26112 24306 26124
rect 24705 26121 24717 26124
rect 24751 26152 24763 26155
rect 25533 26155 25591 26161
rect 25533 26152 25545 26155
rect 24751 26124 25545 26152
rect 24751 26121 24763 26124
rect 24705 26115 24763 26121
rect 25533 26121 25545 26124
rect 25579 26121 25591 26155
rect 25533 26115 25591 26121
rect 18262 26084 18268 26096
rect 18004 26056 18268 26084
rect 18262 26044 18268 26056
rect 18320 26044 18326 26096
rect 25441 26087 25499 26093
rect 25441 26053 25453 26087
rect 25487 26084 25499 26087
rect 25640 26084 25668 26192
rect 27094 26180 27100 26232
rect 27152 26220 27158 26232
rect 27189 26223 27247 26229
rect 27189 26220 27201 26223
rect 27152 26192 27201 26220
rect 27152 26180 27158 26192
rect 27189 26189 27201 26192
rect 27235 26220 27247 26223
rect 27649 26223 27707 26229
rect 27649 26220 27661 26223
rect 27235 26192 27661 26220
rect 27235 26189 27247 26192
rect 27189 26183 27247 26189
rect 27649 26189 27661 26192
rect 27695 26189 27707 26223
rect 27649 26183 27707 26189
rect 29397 26223 29455 26229
rect 29397 26189 29409 26223
rect 29443 26220 29455 26223
rect 29854 26220 29860 26232
rect 29443 26192 29860 26220
rect 29443 26189 29455 26192
rect 29397 26183 29455 26189
rect 29854 26180 29860 26192
rect 29912 26180 29918 26232
rect 27005 26155 27063 26161
rect 27005 26121 27017 26155
rect 27051 26152 27063 26155
rect 27833 26155 27891 26161
rect 27833 26152 27845 26155
rect 27051 26124 27845 26152
rect 27051 26121 27063 26124
rect 27005 26115 27063 26121
rect 27833 26121 27845 26124
rect 27879 26121 27891 26155
rect 27833 26115 27891 26121
rect 25898 26084 25904 26096
rect 25487 26056 25904 26084
rect 25487 26053 25499 26056
rect 25441 26047 25499 26053
rect 25898 26044 25904 26056
rect 25956 26044 25962 26096
rect 27020 26084 27048 26115
rect 29302 26112 29308 26164
rect 29360 26152 29366 26164
rect 29673 26155 29731 26161
rect 29673 26152 29685 26155
rect 29360 26124 29685 26152
rect 29360 26112 29366 26124
rect 29673 26121 29685 26124
rect 29719 26152 29731 26155
rect 29949 26155 30007 26161
rect 29949 26152 29961 26155
rect 29719 26124 29961 26152
rect 29719 26121 29731 26124
rect 29673 26115 29731 26121
rect 29949 26121 29961 26124
rect 29995 26121 30007 26155
rect 29949 26115 30007 26121
rect 27186 26084 27192 26096
rect 27020 26056 27192 26084
rect 27186 26044 27192 26056
rect 27244 26044 27250 26096
rect 29854 26044 29860 26096
rect 29912 26084 29918 26096
rect 30133 26087 30191 26093
rect 30133 26084 30145 26087
rect 29912 26056 30145 26084
rect 29912 26044 29918 26056
rect 30133 26053 30145 26056
rect 30179 26053 30191 26087
rect 30133 26047 30191 26053
rect 400 25994 31680 26016
rect 400 25942 18870 25994
rect 18922 25942 18934 25994
rect 18986 25942 18998 25994
rect 19050 25942 19062 25994
rect 19114 25942 19126 25994
rect 19178 25942 31680 25994
rect 400 25920 31680 25942
rect 1797 25883 1855 25889
rect 1797 25849 1809 25883
rect 1843 25880 1855 25883
rect 1886 25880 1892 25892
rect 1843 25852 1892 25880
rect 1843 25849 1855 25852
rect 1797 25843 1855 25849
rect 1886 25840 1892 25852
rect 1944 25880 1950 25892
rect 2622 25880 2628 25892
rect 1944 25852 2628 25880
rect 1944 25840 1950 25852
rect 2622 25840 2628 25852
rect 2680 25840 2686 25892
rect 8694 25880 8700 25892
rect 8655 25852 8700 25880
rect 8694 25840 8700 25852
rect 8752 25840 8758 25892
rect 9525 25883 9583 25889
rect 9525 25849 9537 25883
rect 9571 25880 9583 25883
rect 9982 25880 9988 25892
rect 9571 25852 9988 25880
rect 9571 25849 9583 25852
rect 9525 25843 9583 25849
rect 3082 25772 3088 25824
rect 3140 25812 3146 25824
rect 6026 25812 6032 25824
rect 3140 25784 4416 25812
rect 5987 25784 6032 25812
rect 3140 25772 3146 25784
rect 3358 25704 3364 25756
rect 3416 25744 3422 25756
rect 4388 25753 4416 25784
rect 6026 25772 6032 25784
rect 6084 25772 6090 25824
rect 6578 25772 6584 25824
rect 6636 25812 6642 25824
rect 6673 25815 6731 25821
rect 6673 25812 6685 25815
rect 6636 25784 6685 25812
rect 6636 25772 6642 25784
rect 6673 25781 6685 25784
rect 6719 25812 6731 25815
rect 9540 25812 9568 25843
rect 9982 25840 9988 25852
rect 10040 25840 10046 25892
rect 14674 25880 14680 25892
rect 14635 25852 14680 25880
rect 14674 25840 14680 25852
rect 14732 25840 14738 25892
rect 14858 25840 14864 25892
rect 14916 25880 14922 25892
rect 15137 25883 15195 25889
rect 15137 25880 15149 25883
rect 14916 25852 15149 25880
rect 14916 25840 14922 25852
rect 15137 25849 15149 25852
rect 15183 25849 15195 25883
rect 15318 25880 15324 25892
rect 15279 25852 15324 25880
rect 15137 25843 15195 25849
rect 15318 25840 15324 25852
rect 15376 25840 15382 25892
rect 23785 25883 23843 25889
rect 23785 25849 23797 25883
rect 23831 25880 23843 25883
rect 24886 25880 24892 25892
rect 23831 25852 24892 25880
rect 23831 25849 23843 25852
rect 23785 25843 23843 25849
rect 24886 25840 24892 25852
rect 24944 25840 24950 25892
rect 6719 25784 9568 25812
rect 6719 25781 6731 25784
rect 6673 25775 6731 25781
rect 15042 25772 15048 25824
rect 15100 25812 15106 25824
rect 16149 25815 16207 25821
rect 16149 25812 16161 25815
rect 15100 25784 16161 25812
rect 15100 25772 15106 25784
rect 16149 25781 16161 25784
rect 16195 25781 16207 25815
rect 18357 25815 18415 25821
rect 18357 25812 18369 25815
rect 16149 25775 16207 25781
rect 17820 25784 18369 25812
rect 4005 25747 4063 25753
rect 4005 25744 4017 25747
rect 3416 25716 4017 25744
rect 3416 25704 3422 25716
rect 4005 25713 4017 25716
rect 4051 25713 4063 25747
rect 4005 25707 4063 25713
rect 4373 25747 4431 25753
rect 4373 25713 4385 25747
rect 4419 25713 4431 25747
rect 5750 25744 5756 25756
rect 5711 25716 5756 25744
rect 4373 25707 4431 25713
rect 5750 25704 5756 25716
rect 5808 25704 5814 25756
rect 7682 25704 7688 25756
rect 7740 25744 7746 25756
rect 9249 25747 9307 25753
rect 9249 25744 9261 25747
rect 7740 25716 9261 25744
rect 7740 25704 7746 25716
rect 9249 25713 9261 25716
rect 9295 25744 9307 25747
rect 9798 25744 9804 25756
rect 9295 25716 9804 25744
rect 9295 25713 9307 25716
rect 9249 25707 9307 25713
rect 9798 25704 9804 25716
rect 9856 25744 9862 25756
rect 10350 25744 10356 25756
rect 9856 25716 10356 25744
rect 9856 25704 9862 25716
rect 10350 25704 10356 25716
rect 10408 25704 10414 25756
rect 14953 25747 15011 25753
rect 14953 25713 14965 25747
rect 14999 25744 15011 25747
rect 15134 25744 15140 25756
rect 14999 25716 15140 25744
rect 14999 25713 15011 25716
rect 14953 25707 15011 25713
rect 15134 25704 15140 25716
rect 15192 25704 15198 25756
rect 16790 25704 16796 25756
rect 16848 25744 16854 25756
rect 17820 25753 17848 25784
rect 18357 25781 18369 25784
rect 18403 25781 18415 25815
rect 18357 25775 18415 25781
rect 22494 25772 22500 25824
rect 22552 25772 22558 25824
rect 27281 25815 27339 25821
rect 27281 25781 27293 25815
rect 27327 25812 27339 25815
rect 27554 25812 27560 25824
rect 27327 25784 27560 25812
rect 27327 25781 27339 25784
rect 27281 25775 27339 25781
rect 27554 25772 27560 25784
rect 27612 25772 27618 25824
rect 17805 25747 17863 25753
rect 17805 25744 17817 25747
rect 16848 25716 17817 25744
rect 16848 25704 16854 25716
rect 17805 25713 17817 25716
rect 17851 25713 17863 25747
rect 17805 25707 17863 25713
rect 18265 25747 18323 25753
rect 18265 25713 18277 25747
rect 18311 25744 18323 25747
rect 18446 25744 18452 25756
rect 18311 25716 18452 25744
rect 18311 25713 18323 25716
rect 18265 25707 18323 25713
rect 18446 25704 18452 25716
rect 18504 25704 18510 25756
rect 20194 25744 20200 25756
rect 20155 25716 20200 25744
rect 20194 25704 20200 25716
rect 20252 25704 20258 25756
rect 21390 25704 21396 25756
rect 21448 25744 21454 25756
rect 21577 25747 21635 25753
rect 21577 25744 21589 25747
rect 21448 25716 21589 25744
rect 21448 25704 21454 25716
rect 21577 25713 21589 25716
rect 21623 25713 21635 25747
rect 24518 25744 24524 25756
rect 24479 25716 24524 25744
rect 21577 25707 21635 25713
rect 24518 25704 24524 25716
rect 24576 25704 24582 25756
rect 26726 25744 26732 25756
rect 26687 25716 26732 25744
rect 26726 25704 26732 25716
rect 26784 25704 26790 25756
rect 26913 25747 26971 25753
rect 26913 25713 26925 25747
rect 26959 25744 26971 25747
rect 27094 25744 27100 25756
rect 26959 25716 27100 25744
rect 26959 25713 26971 25716
rect 26913 25707 26971 25713
rect 27094 25704 27100 25716
rect 27152 25704 27158 25756
rect 27830 25704 27836 25756
rect 27888 25744 27894 25756
rect 28109 25747 28167 25753
rect 28109 25744 28121 25747
rect 27888 25716 28121 25744
rect 27888 25704 27894 25716
rect 28109 25713 28121 25716
rect 28155 25713 28167 25747
rect 28109 25707 28167 25713
rect 690 25636 696 25688
rect 748 25676 754 25688
rect 877 25679 935 25685
rect 877 25676 889 25679
rect 748 25648 889 25676
rect 748 25636 754 25648
rect 877 25645 889 25648
rect 923 25645 935 25679
rect 877 25639 935 25645
rect 2714 25636 2720 25688
rect 2772 25676 2778 25688
rect 3453 25679 3511 25685
rect 3453 25676 3465 25679
rect 2772 25648 3465 25676
rect 2772 25636 2778 25648
rect 3453 25645 3465 25648
rect 3499 25645 3511 25679
rect 3910 25676 3916 25688
rect 3871 25648 3916 25676
rect 3453 25639 3511 25645
rect 782 25540 788 25552
rect 743 25512 788 25540
rect 782 25500 788 25512
rect 840 25500 846 25552
rect 3468 25540 3496 25639
rect 3910 25636 3916 25648
rect 3968 25636 3974 25688
rect 4278 25676 4284 25688
rect 4239 25648 4284 25676
rect 4278 25636 4284 25648
rect 4336 25636 4342 25688
rect 6857 25679 6915 25685
rect 6857 25645 6869 25679
rect 6903 25676 6915 25679
rect 7222 25676 7228 25688
rect 6903 25648 7228 25676
rect 6903 25645 6915 25648
rect 6857 25639 6915 25645
rect 7222 25636 7228 25648
rect 7280 25676 7286 25688
rect 12742 25676 12748 25688
rect 7280 25648 12748 25676
rect 7280 25636 7286 25648
rect 12742 25636 12748 25648
rect 12800 25636 12806 25688
rect 15502 25636 15508 25688
rect 15560 25676 15566 25688
rect 16330 25676 16336 25688
rect 15560 25648 16336 25676
rect 15560 25636 15566 25648
rect 16330 25636 16336 25648
rect 16388 25676 16394 25688
rect 16517 25679 16575 25685
rect 16517 25676 16529 25679
rect 16388 25648 16529 25676
rect 16388 25636 16394 25648
rect 16517 25645 16529 25648
rect 16563 25645 16575 25679
rect 17710 25676 17716 25688
rect 17623 25648 17716 25676
rect 16517 25639 16575 25645
rect 17710 25636 17716 25648
rect 17768 25676 17774 25688
rect 18170 25676 18176 25688
rect 17768 25648 18176 25676
rect 17768 25636 17774 25648
rect 18170 25636 18176 25648
rect 18228 25636 18234 25688
rect 20378 25676 20384 25688
rect 20339 25648 20384 25676
rect 20378 25636 20384 25648
rect 20436 25636 20442 25688
rect 21850 25676 21856 25688
rect 21811 25648 21856 25676
rect 21850 25636 21856 25648
rect 21908 25636 21914 25688
rect 22218 25636 22224 25688
rect 22276 25676 22282 25688
rect 23230 25676 23236 25688
rect 22276 25648 23236 25676
rect 22276 25636 22282 25648
rect 23230 25636 23236 25648
rect 23288 25676 23294 25688
rect 23601 25679 23659 25685
rect 23601 25676 23613 25679
rect 23288 25648 23613 25676
rect 23288 25636 23294 25648
rect 23601 25645 23613 25648
rect 23647 25645 23659 25679
rect 23601 25639 23659 25645
rect 28385 25679 28443 25685
rect 28385 25645 28397 25679
rect 28431 25676 28443 25679
rect 28566 25676 28572 25688
rect 28431 25648 28572 25676
rect 28431 25645 28443 25648
rect 28385 25639 28443 25645
rect 28566 25636 28572 25648
rect 28624 25676 28630 25688
rect 28661 25679 28719 25685
rect 28661 25676 28673 25679
rect 28624 25648 28673 25676
rect 28624 25636 28630 25648
rect 28661 25645 28673 25648
rect 28707 25645 28719 25679
rect 28661 25639 28719 25645
rect 6486 25568 6492 25620
rect 6544 25608 6550 25620
rect 10626 25608 10632 25620
rect 6544 25580 10632 25608
rect 6544 25568 6550 25580
rect 10626 25568 10632 25580
rect 10684 25568 10690 25620
rect 15594 25568 15600 25620
rect 15652 25608 15658 25620
rect 16609 25611 16667 25617
rect 16609 25608 16621 25611
rect 15652 25580 16621 25608
rect 15652 25568 15658 25580
rect 16609 25577 16621 25580
rect 16655 25577 16667 25611
rect 16609 25571 16667 25577
rect 17437 25611 17495 25617
rect 17437 25577 17449 25611
rect 17483 25608 17495 25611
rect 18262 25608 18268 25620
rect 17483 25580 18268 25608
rect 17483 25577 17495 25580
rect 17437 25571 17495 25577
rect 18262 25568 18268 25580
rect 18320 25568 18326 25620
rect 4922 25540 4928 25552
rect 3468 25512 4928 25540
rect 4922 25500 4928 25512
rect 4980 25500 4986 25552
rect 9614 25540 9620 25552
rect 9575 25512 9620 25540
rect 9614 25500 9620 25512
rect 9672 25500 9678 25552
rect 13018 25500 13024 25552
rect 13076 25540 13082 25552
rect 14674 25540 14680 25552
rect 13076 25512 14680 25540
rect 13076 25500 13082 25512
rect 14674 25500 14680 25512
rect 14732 25500 14738 25552
rect 16238 25500 16244 25552
rect 16296 25549 16302 25552
rect 16296 25543 16345 25549
rect 16296 25509 16299 25543
rect 16333 25509 16345 25543
rect 16422 25540 16428 25552
rect 16383 25512 16428 25540
rect 16296 25503 16345 25509
rect 16296 25500 16302 25503
rect 16422 25500 16428 25512
rect 16480 25500 16486 25552
rect 17342 25500 17348 25552
rect 17400 25540 17406 25552
rect 17529 25543 17587 25549
rect 17529 25540 17541 25543
rect 17400 25512 17541 25540
rect 17400 25500 17406 25512
rect 17529 25509 17541 25512
rect 17575 25509 17587 25543
rect 17529 25503 17587 25509
rect 24426 25500 24432 25552
rect 24484 25540 24490 25552
rect 24613 25543 24671 25549
rect 24613 25540 24625 25543
rect 24484 25512 24625 25540
rect 24484 25500 24490 25512
rect 24613 25509 24625 25512
rect 24659 25509 24671 25543
rect 24613 25503 24671 25509
rect 400 25450 31680 25472
rect 400 25398 3510 25450
rect 3562 25398 3574 25450
rect 3626 25398 3638 25450
rect 3690 25398 3702 25450
rect 3754 25398 3766 25450
rect 3818 25398 31680 25450
rect 400 25376 31680 25398
rect 3453 25339 3511 25345
rect 3453 25305 3465 25339
rect 3499 25336 3511 25339
rect 4278 25336 4284 25348
rect 3499 25308 4284 25336
rect 3499 25305 3511 25308
rect 3453 25299 3511 25305
rect 4278 25296 4284 25308
rect 4336 25336 4342 25348
rect 4922 25336 4928 25348
rect 4336 25308 4784 25336
rect 4883 25308 4928 25336
rect 4336 25296 4342 25308
rect 782 25228 788 25280
rect 840 25268 846 25280
rect 1613 25271 1671 25277
rect 1613 25268 1625 25271
rect 840 25240 1625 25268
rect 840 25228 846 25240
rect 1613 25237 1625 25240
rect 1659 25268 1671 25271
rect 2073 25271 2131 25277
rect 2073 25268 2085 25271
rect 1659 25240 2085 25268
rect 1659 25237 1671 25240
rect 1613 25231 1671 25237
rect 2073 25237 2085 25240
rect 2119 25237 2131 25271
rect 3266 25268 3272 25280
rect 3179 25240 3272 25268
rect 2073 25231 2131 25237
rect 3266 25228 3272 25240
rect 3324 25268 3330 25280
rect 4756 25268 4784 25308
rect 4922 25296 4928 25308
rect 4980 25296 4986 25348
rect 5661 25339 5719 25345
rect 5661 25305 5673 25339
rect 5707 25336 5719 25339
rect 6026 25336 6032 25348
rect 5707 25308 6032 25336
rect 5707 25305 5719 25308
rect 5661 25299 5719 25305
rect 6026 25296 6032 25308
rect 6084 25296 6090 25348
rect 12469 25339 12527 25345
rect 12469 25305 12481 25339
rect 12515 25336 12527 25339
rect 12558 25336 12564 25348
rect 12515 25308 12564 25336
rect 12515 25305 12527 25308
rect 12469 25299 12527 25305
rect 12558 25296 12564 25308
rect 12616 25336 12622 25348
rect 12837 25339 12895 25345
rect 12837 25336 12849 25339
rect 12616 25308 12849 25336
rect 12616 25296 12622 25308
rect 12837 25305 12849 25308
rect 12883 25305 12895 25339
rect 12837 25299 12895 25305
rect 16241 25339 16299 25345
rect 16241 25305 16253 25339
rect 16287 25336 16299 25339
rect 16422 25336 16428 25348
rect 16287 25308 16428 25336
rect 16287 25305 16299 25308
rect 16241 25299 16299 25305
rect 16422 25296 16428 25308
rect 16480 25296 16486 25348
rect 20194 25336 20200 25348
rect 20155 25308 20200 25336
rect 20194 25296 20200 25308
rect 20252 25296 20258 25348
rect 21301 25339 21359 25345
rect 21301 25305 21313 25339
rect 21347 25336 21359 25339
rect 21390 25336 21396 25348
rect 21347 25308 21396 25336
rect 21347 25305 21359 25308
rect 21301 25299 21359 25305
rect 21390 25296 21396 25308
rect 21448 25296 21454 25348
rect 22218 25336 22224 25348
rect 22179 25308 22224 25336
rect 22218 25296 22224 25308
rect 22276 25296 22282 25348
rect 22494 25336 22500 25348
rect 22455 25308 22500 25336
rect 22494 25296 22500 25308
rect 22552 25336 22558 25348
rect 22681 25339 22739 25345
rect 22681 25336 22693 25339
rect 22552 25308 22693 25336
rect 22552 25296 22558 25308
rect 22681 25305 22693 25308
rect 22727 25305 22739 25339
rect 23322 25336 23328 25348
rect 23283 25308 23328 25336
rect 22681 25299 22739 25305
rect 23322 25296 23328 25308
rect 23380 25336 23386 25348
rect 23969 25339 24027 25345
rect 23969 25336 23981 25339
rect 23380 25308 23981 25336
rect 23380 25296 23386 25308
rect 23969 25305 23981 25308
rect 24015 25305 24027 25339
rect 23969 25299 24027 25305
rect 24518 25296 24524 25348
rect 24576 25336 24582 25348
rect 24981 25339 25039 25345
rect 24981 25336 24993 25339
rect 24576 25308 24993 25336
rect 24576 25296 24582 25308
rect 24981 25305 24993 25308
rect 25027 25305 25039 25339
rect 24981 25299 25039 25305
rect 26453 25339 26511 25345
rect 26453 25305 26465 25339
rect 26499 25336 26511 25339
rect 26821 25339 26879 25345
rect 26821 25336 26833 25339
rect 26499 25308 26833 25336
rect 26499 25305 26511 25308
rect 26453 25299 26511 25305
rect 26821 25305 26833 25308
rect 26867 25336 26879 25339
rect 27094 25336 27100 25348
rect 26867 25308 27100 25336
rect 26867 25305 26879 25308
rect 26821 25299 26879 25305
rect 5750 25268 5756 25280
rect 3324 25240 4416 25268
rect 4756 25240 5756 25268
rect 3324 25228 3330 25240
rect 4388 25209 4416 25240
rect 5750 25228 5756 25240
rect 5808 25268 5814 25280
rect 13205 25271 13263 25277
rect 5808 25240 5888 25268
rect 5808 25228 5814 25240
rect 4373 25203 4431 25209
rect 2180 25172 4140 25200
rect 2180 25141 2208 25172
rect 1429 25135 1487 25141
rect 1429 25101 1441 25135
rect 1475 25132 1487 25135
rect 2165 25135 2223 25141
rect 2165 25132 2177 25135
rect 1475 25104 2177 25132
rect 1475 25101 1487 25104
rect 1429 25095 1487 25101
rect 2165 25101 2177 25104
rect 2211 25101 2223 25135
rect 2346 25132 2352 25144
rect 2307 25104 2352 25132
rect 2165 25095 2223 25101
rect 2346 25092 2352 25104
rect 2404 25092 2410 25144
rect 2622 25132 2628 25144
rect 2583 25104 2628 25132
rect 2622 25092 2628 25104
rect 2680 25092 2686 25144
rect 2714 25092 2720 25144
rect 2772 25132 2778 25144
rect 4112 25141 4140 25172
rect 4373 25169 4385 25203
rect 4419 25169 4431 25203
rect 4373 25163 4431 25169
rect 4097 25135 4155 25141
rect 2772 25104 2865 25132
rect 2772 25092 2778 25104
rect 4097 25101 4109 25135
rect 4143 25132 4155 25135
rect 4554 25132 4560 25144
rect 4143 25104 4560 25132
rect 4143 25101 4155 25104
rect 4097 25095 4155 25101
rect 4554 25092 4560 25104
rect 4612 25092 4618 25144
rect 1245 25067 1303 25073
rect 1245 25033 1257 25067
rect 1291 25064 1303 25067
rect 2732 25064 2760 25092
rect 1291 25036 2760 25064
rect 3913 25067 3971 25073
rect 1291 25033 1303 25036
rect 1245 25027 1303 25033
rect 3913 25033 3925 25067
rect 3959 25064 3971 25067
rect 4278 25064 4284 25076
rect 3959 25036 4284 25064
rect 3959 25033 3971 25036
rect 3913 25027 3971 25033
rect 4278 25024 4284 25036
rect 4336 25064 4342 25076
rect 4741 25067 4799 25073
rect 4741 25064 4753 25067
rect 4336 25036 4753 25064
rect 4336 25024 4342 25036
rect 4741 25033 4753 25036
rect 4787 25033 4799 25067
rect 4741 25027 4799 25033
rect 3082 24956 3088 25008
rect 3140 24996 3146 25008
rect 3545 24999 3603 25005
rect 3545 24996 3557 24999
rect 3140 24968 3557 24996
rect 3140 24956 3146 24968
rect 3545 24965 3557 24968
rect 3591 24965 3603 24999
rect 3818 24996 3824 25008
rect 3779 24968 3824 24996
rect 3545 24959 3603 24965
rect 3818 24956 3824 24968
rect 3876 24956 3882 25008
rect 4554 24996 4560 25008
rect 4515 24968 4560 24996
rect 4554 24956 4560 24968
rect 4612 24956 4618 25008
rect 5860 25005 5888 25240
rect 13205 25237 13217 25271
rect 13251 25268 13263 25271
rect 14950 25268 14956 25280
rect 13251 25240 14956 25268
rect 13251 25237 13263 25240
rect 13205 25231 13263 25237
rect 14950 25228 14956 25240
rect 15008 25228 15014 25280
rect 16330 25268 16336 25280
rect 16291 25240 16336 25268
rect 16330 25228 16336 25240
rect 16388 25228 16394 25280
rect 16790 25268 16796 25280
rect 16751 25240 16796 25268
rect 16790 25228 16796 25240
rect 16848 25228 16854 25280
rect 18630 25228 18636 25280
rect 18688 25268 18694 25280
rect 20378 25268 20384 25280
rect 18688 25240 20384 25268
rect 18688 25228 18694 25240
rect 20378 25228 20384 25240
rect 20436 25268 20442 25280
rect 21025 25271 21083 25277
rect 21025 25268 21037 25271
rect 20436 25240 21037 25268
rect 20436 25228 20442 25240
rect 21025 25237 21037 25240
rect 21071 25237 21083 25271
rect 21025 25231 21083 25237
rect 10442 25200 10448 25212
rect 10355 25172 10448 25200
rect 5934 25092 5940 25144
rect 5992 25132 5998 25144
rect 10368 25141 10396 25172
rect 10442 25160 10448 25172
rect 10500 25200 10506 25212
rect 10997 25203 11055 25209
rect 10997 25200 11009 25203
rect 10500 25172 11009 25200
rect 10500 25160 10506 25172
rect 10997 25169 11009 25172
rect 11043 25200 11055 25203
rect 16238 25200 16244 25212
rect 11043 25172 16244 25200
rect 11043 25169 11055 25172
rect 10997 25163 11055 25169
rect 16238 25160 16244 25172
rect 16296 25200 16302 25212
rect 16609 25203 16667 25209
rect 16609 25200 16621 25203
rect 16296 25172 16621 25200
rect 16296 25160 16302 25172
rect 16609 25169 16621 25172
rect 16655 25200 16667 25203
rect 18354 25200 18360 25212
rect 16655 25172 18360 25200
rect 16655 25169 16667 25172
rect 16609 25163 16667 25169
rect 18354 25160 18360 25172
rect 18412 25160 18418 25212
rect 20013 25203 20071 25209
rect 20013 25169 20025 25203
rect 20059 25200 20071 25203
rect 20473 25203 20531 25209
rect 20473 25200 20485 25203
rect 20059 25172 20485 25200
rect 20059 25169 20071 25172
rect 20013 25163 20071 25169
rect 20473 25169 20485 25172
rect 20519 25200 20531 25203
rect 21666 25200 21672 25212
rect 20519 25172 21672 25200
rect 20519 25169 20531 25172
rect 20473 25163 20531 25169
rect 21666 25160 21672 25172
rect 21724 25160 21730 25212
rect 21853 25203 21911 25209
rect 21853 25169 21865 25203
rect 21899 25200 21911 25203
rect 22512 25200 22540 25296
rect 23601 25271 23659 25277
rect 23601 25237 23613 25271
rect 23647 25268 23659 25271
rect 24536 25268 24564 25296
rect 24886 25268 24892 25280
rect 23647 25240 24564 25268
rect 24799 25240 24892 25268
rect 23647 25237 23659 25240
rect 23601 25231 23659 25237
rect 24444 25209 24472 25240
rect 24886 25228 24892 25240
rect 24944 25268 24950 25280
rect 26174 25268 26180 25280
rect 24944 25240 26180 25268
rect 24944 25228 24950 25240
rect 26174 25228 26180 25240
rect 26232 25228 26238 25280
rect 24429 25203 24487 25209
rect 21899 25172 22540 25200
rect 23846 25172 24380 25200
rect 21899 25169 21911 25172
rect 21853 25163 21911 25169
rect 6121 25135 6179 25141
rect 6121 25132 6133 25135
rect 5992 25104 6133 25132
rect 5992 25092 5998 25104
rect 6121 25101 6133 25104
rect 6167 25132 6179 25135
rect 6673 25135 6731 25141
rect 6673 25132 6685 25135
rect 6167 25104 6685 25132
rect 6167 25101 6179 25104
rect 6121 25095 6179 25101
rect 6673 25101 6685 25104
rect 6719 25101 6731 25135
rect 6673 25095 6731 25101
rect 10353 25135 10411 25141
rect 10353 25101 10365 25135
rect 10399 25101 10411 25135
rect 10353 25095 10411 25101
rect 12469 25135 12527 25141
rect 12469 25101 12481 25135
rect 12515 25132 12527 25135
rect 17342 25132 17348 25144
rect 12515 25104 12696 25132
rect 17303 25104 17348 25132
rect 12515 25101 12527 25104
rect 12469 25095 12527 25101
rect 6394 25064 6400 25076
rect 6355 25036 6400 25064
rect 6394 25024 6400 25036
rect 6452 25064 6458 25076
rect 6857 25067 6915 25073
rect 6857 25064 6869 25067
rect 6452 25036 6869 25064
rect 6452 25024 6458 25036
rect 6857 25033 6869 25036
rect 6903 25064 6915 25067
rect 8234 25064 8240 25076
rect 6903 25036 8240 25064
rect 6903 25033 6915 25036
rect 6857 25027 6915 25033
rect 8234 25024 8240 25036
rect 8292 25024 8298 25076
rect 10629 25067 10687 25073
rect 10629 25033 10641 25067
rect 10675 25064 10687 25067
rect 10675 25036 11224 25064
rect 10675 25033 10687 25036
rect 10629 25027 10687 25033
rect 5845 24999 5903 25005
rect 5845 24965 5857 24999
rect 5891 24996 5903 24999
rect 7038 24996 7044 25008
rect 5891 24968 7044 24996
rect 5891 24965 5903 24968
rect 5845 24959 5903 24965
rect 7038 24956 7044 24968
rect 7096 24956 7102 25008
rect 11196 25005 11224 25036
rect 12668 25008 12696 25104
rect 17342 25092 17348 25104
rect 17400 25092 17406 25144
rect 20286 25132 20292 25144
rect 20247 25104 20292 25132
rect 20286 25092 20292 25104
rect 20344 25132 20350 25144
rect 20654 25132 20660 25144
rect 20344 25104 20660 25132
rect 20344 25092 20350 25104
rect 20654 25092 20660 25104
rect 20712 25132 20718 25144
rect 20841 25135 20899 25141
rect 20841 25132 20853 25135
rect 20712 25104 20853 25132
rect 20712 25092 20718 25104
rect 20841 25101 20853 25104
rect 20887 25132 20899 25135
rect 21393 25135 21451 25141
rect 21393 25132 21405 25135
rect 20887 25104 21405 25132
rect 20887 25101 20899 25104
rect 20841 25095 20899 25101
rect 21393 25101 21405 25104
rect 21439 25132 21451 25135
rect 21577 25135 21635 25141
rect 21577 25132 21589 25135
rect 21439 25104 21589 25132
rect 21439 25101 21451 25104
rect 21393 25095 21451 25101
rect 21577 25101 21589 25104
rect 21623 25101 21635 25135
rect 23846 25132 23874 25172
rect 24352 25141 24380 25172
rect 24429 25169 24441 25203
rect 24475 25169 24487 25203
rect 24429 25163 24487 25169
rect 21577 25095 21635 25101
rect 23156 25104 23874 25132
rect 24337 25135 24395 25141
rect 13481 25067 13539 25073
rect 13481 25033 13493 25067
rect 13527 25064 13539 25067
rect 16882 25064 16888 25076
rect 13527 25036 16888 25064
rect 13527 25033 13539 25036
rect 13481 25027 13539 25033
rect 11181 24999 11239 25005
rect 11181 24965 11193 24999
rect 11227 24996 11239 24999
rect 11454 24996 11460 25008
rect 11227 24968 11460 24996
rect 11227 24965 11239 24968
rect 11181 24959 11239 24965
rect 11454 24956 11460 24968
rect 11512 24956 11518 25008
rect 12650 24996 12656 25008
rect 12611 24968 12656 24996
rect 12650 24956 12656 24968
rect 12708 24956 12714 25008
rect 13294 24996 13300 25008
rect 13255 24968 13300 24996
rect 13294 24956 13300 24968
rect 13352 24996 13358 25008
rect 13496 24996 13524 25027
rect 16882 25024 16888 25036
rect 16940 25024 16946 25076
rect 17621 25067 17679 25073
rect 17621 25064 17633 25067
rect 16992 25036 17633 25064
rect 16992 25008 17020 25036
rect 17621 25033 17633 25036
rect 17667 25033 17679 25067
rect 17621 25027 17679 25033
rect 18262 25024 18268 25076
rect 18320 25024 18326 25076
rect 19366 25064 19372 25076
rect 19327 25036 19372 25064
rect 19366 25024 19372 25036
rect 19424 25024 19430 25076
rect 21850 25024 21856 25076
rect 21908 25064 21914 25076
rect 22313 25067 22371 25073
rect 22313 25064 22325 25067
rect 21908 25036 22325 25064
rect 21908 25024 21914 25036
rect 22313 25033 22325 25036
rect 22359 25033 22371 25067
rect 22313 25027 22371 25033
rect 14950 24996 14956 25008
rect 13352 24968 13524 24996
rect 14911 24968 14956 24996
rect 13352 24956 13358 24968
rect 14950 24956 14956 24968
rect 15008 24956 15014 25008
rect 15594 24956 15600 25008
rect 15652 24996 15658 25008
rect 15965 24999 16023 25005
rect 15965 24996 15977 24999
rect 15652 24968 15977 24996
rect 15652 24956 15658 24968
rect 15965 24965 15977 24968
rect 16011 24965 16023 24999
rect 16974 24996 16980 25008
rect 16935 24968 16980 24996
rect 15965 24959 16023 24965
rect 16974 24956 16980 24968
rect 17032 24956 17038 25008
rect 17066 24956 17072 25008
rect 17124 24996 17130 25008
rect 17161 24999 17219 25005
rect 17161 24996 17173 24999
rect 17124 24968 17173 24996
rect 17124 24956 17130 24968
rect 17161 24965 17173 24968
rect 17207 24996 17219 24999
rect 17894 24996 17900 25008
rect 17207 24968 17900 24996
rect 17207 24965 17219 24968
rect 17161 24959 17219 24965
rect 17894 24956 17900 24968
rect 17952 24956 17958 25008
rect 22586 24956 22592 25008
rect 22644 24996 22650 25008
rect 23156 25005 23184 25104
rect 24337 25101 24349 25135
rect 24383 25132 24395 25135
rect 24518 25132 24524 25144
rect 24383 25104 24524 25132
rect 24383 25101 24395 25104
rect 24337 25095 24395 25101
rect 24518 25092 24524 25104
rect 24576 25092 24582 25144
rect 24702 25132 24708 25144
rect 24663 25104 24708 25132
rect 24702 25092 24708 25104
rect 24760 25092 24766 25144
rect 24904 25141 24932 25228
rect 24889 25135 24947 25141
rect 24889 25101 24901 25135
rect 24935 25101 24947 25135
rect 24889 25095 24947 25101
rect 25809 25135 25867 25141
rect 25809 25101 25821 25135
rect 25855 25132 25867 25135
rect 26174 25132 26180 25144
rect 25855 25104 26180 25132
rect 25855 25101 25867 25104
rect 25809 25095 25867 25101
rect 26174 25092 26180 25104
rect 26232 25132 26238 25144
rect 26468 25132 26496 25299
rect 27094 25296 27100 25308
rect 27152 25296 27158 25348
rect 27189 25339 27247 25345
rect 27189 25305 27201 25339
rect 27235 25336 27247 25339
rect 27554 25336 27560 25348
rect 27235 25308 27560 25336
rect 27235 25305 27247 25308
rect 27189 25299 27247 25305
rect 27554 25296 27560 25308
rect 27612 25296 27618 25348
rect 28017 25203 28075 25209
rect 28017 25169 28029 25203
rect 28063 25200 28075 25203
rect 28566 25200 28572 25212
rect 28063 25172 28572 25200
rect 28063 25169 28075 25172
rect 28017 25163 28075 25169
rect 28566 25160 28572 25172
rect 28624 25160 28630 25212
rect 26232 25104 26496 25132
rect 26232 25092 26238 25104
rect 26726 25092 26732 25144
rect 26784 25132 26790 25144
rect 26913 25135 26971 25141
rect 26913 25132 26925 25135
rect 26784 25104 26925 25132
rect 26784 25092 26790 25104
rect 26913 25101 26925 25104
rect 26959 25101 26971 25135
rect 26913 25095 26971 25101
rect 24426 25024 24432 25076
rect 24484 25064 24490 25076
rect 25165 25067 25223 25073
rect 25165 25064 25177 25067
rect 24484 25036 25177 25064
rect 24484 25024 24490 25036
rect 25165 25033 25177 25036
rect 25211 25033 25223 25067
rect 25165 25027 25223 25033
rect 25898 25024 25904 25076
rect 25956 25064 25962 25076
rect 26085 25067 26143 25073
rect 26085 25064 26097 25067
rect 25956 25036 26097 25064
rect 25956 25024 25962 25036
rect 26085 25033 26097 25036
rect 26131 25064 26143 25067
rect 28201 25067 28259 25073
rect 26131 25036 26588 25064
rect 26131 25033 26143 25036
rect 26085 25027 26143 25033
rect 26560 25008 26588 25036
rect 28201 25033 28213 25067
rect 28247 25064 28259 25067
rect 28382 25064 28388 25076
rect 28247 25036 28388 25064
rect 28247 25033 28259 25036
rect 28201 25027 28259 25033
rect 28382 25024 28388 25036
rect 28440 25064 28446 25076
rect 28845 25067 28903 25073
rect 28845 25064 28857 25067
rect 28440 25036 28857 25064
rect 28440 25024 28446 25036
rect 28845 25033 28857 25036
rect 28891 25033 28903 25067
rect 28845 25027 28903 25033
rect 29302 25024 29308 25076
rect 29360 25024 29366 25076
rect 30590 25064 30596 25076
rect 30551 25036 30596 25064
rect 30590 25024 30596 25036
rect 30648 25024 30654 25076
rect 23141 24999 23199 25005
rect 23141 24996 23153 24999
rect 22644 24968 23153 24996
rect 22644 24956 22650 24968
rect 23141 24965 23153 24968
rect 23187 24965 23199 24999
rect 26542 24996 26548 25008
rect 26503 24968 26548 24996
rect 23141 24959 23199 24965
rect 26542 24956 26548 24968
rect 26600 24956 26606 25008
rect 27830 24996 27836 25008
rect 27791 24968 27836 24996
rect 27830 24956 27836 24968
rect 27888 24956 27894 25008
rect 28293 24999 28351 25005
rect 28293 24965 28305 24999
rect 28339 24996 28351 24999
rect 28474 24996 28480 25008
rect 28339 24968 28480 24996
rect 28339 24965 28351 24968
rect 28293 24959 28351 24965
rect 28474 24956 28480 24968
rect 28532 24956 28538 25008
rect 400 24906 31680 24928
rect 400 24854 18870 24906
rect 18922 24854 18934 24906
rect 18986 24854 18998 24906
rect 19050 24854 19062 24906
rect 19114 24854 19126 24906
rect 19178 24854 31680 24906
rect 400 24832 31680 24854
rect 1797 24795 1855 24801
rect 1797 24761 1809 24795
rect 1843 24792 1855 24795
rect 1886 24792 1892 24804
rect 1843 24764 1892 24792
rect 1843 24761 1855 24764
rect 1797 24755 1855 24761
rect 1886 24752 1892 24764
rect 1944 24792 1950 24804
rect 2346 24792 2352 24804
rect 1944 24764 2352 24792
rect 1944 24752 1950 24764
rect 2346 24752 2352 24764
rect 2404 24752 2410 24804
rect 3358 24792 3364 24804
rect 3319 24764 3364 24792
rect 3358 24752 3364 24764
rect 3416 24752 3422 24804
rect 18170 24792 18176 24804
rect 18131 24764 18176 24792
rect 18170 24752 18176 24764
rect 18228 24752 18234 24804
rect 23601 24795 23659 24801
rect 23601 24761 23613 24795
rect 23647 24792 23659 24795
rect 24702 24792 24708 24804
rect 23647 24764 24708 24792
rect 23647 24761 23659 24764
rect 23601 24755 23659 24761
rect 24702 24752 24708 24764
rect 24760 24752 24766 24804
rect 28753 24795 28811 24801
rect 28753 24761 28765 24795
rect 28799 24792 28811 24795
rect 29302 24792 29308 24804
rect 28799 24764 29308 24792
rect 28799 24761 28811 24764
rect 28753 24755 28811 24761
rect 29302 24752 29308 24764
rect 29360 24752 29366 24804
rect 1150 24684 1156 24736
rect 1208 24724 1214 24736
rect 7774 24724 7780 24736
rect 1208 24696 7780 24724
rect 1208 24684 1214 24696
rect 4465 24659 4523 24665
rect 4465 24625 4477 24659
rect 4511 24625 4523 24659
rect 4465 24619 4523 24625
rect 3637 24591 3695 24597
rect 3637 24557 3649 24591
rect 3683 24588 3695 24591
rect 3910 24588 3916 24600
rect 3683 24560 3916 24588
rect 3683 24557 3695 24560
rect 3637 24551 3695 24557
rect 3910 24548 3916 24560
rect 3968 24548 3974 24600
rect 4189 24591 4247 24597
rect 4189 24557 4201 24591
rect 4235 24588 4247 24591
rect 4278 24588 4284 24600
rect 4235 24560 4284 24588
rect 4235 24557 4247 24560
rect 4189 24551 4247 24557
rect 4278 24548 4284 24560
rect 4336 24548 4342 24600
rect 4480 24588 4508 24619
rect 4646 24616 4652 24668
rect 4704 24656 4710 24668
rect 5382 24656 5388 24668
rect 4704 24628 5388 24656
rect 4704 24616 4710 24628
rect 5382 24616 5388 24628
rect 5440 24656 5446 24668
rect 5842 24656 5848 24668
rect 5440 24628 5848 24656
rect 5440 24616 5446 24628
rect 5842 24616 5848 24628
rect 5900 24616 5906 24668
rect 7608 24665 7636 24696
rect 7774 24684 7780 24696
rect 7832 24684 7838 24736
rect 16974 24684 16980 24736
rect 17032 24724 17038 24736
rect 17161 24727 17219 24733
rect 17161 24724 17173 24727
rect 17032 24696 17173 24724
rect 17032 24684 17038 24696
rect 17161 24693 17173 24696
rect 17207 24693 17219 24727
rect 17161 24687 17219 24693
rect 21666 24684 21672 24736
rect 21724 24684 21730 24736
rect 26174 24724 26180 24736
rect 26135 24696 26180 24724
rect 26174 24684 26180 24696
rect 26232 24684 26238 24736
rect 7593 24659 7651 24665
rect 7593 24625 7605 24659
rect 7639 24625 7651 24659
rect 9246 24656 9252 24668
rect 9207 24628 9252 24656
rect 7593 24619 7651 24625
rect 9246 24616 9252 24628
rect 9304 24616 9310 24668
rect 15594 24656 15600 24668
rect 15555 24628 15600 24656
rect 15594 24616 15600 24628
rect 15652 24616 15658 24668
rect 15778 24656 15784 24668
rect 15739 24628 15784 24656
rect 15778 24616 15784 24628
rect 15836 24616 15842 24668
rect 17894 24656 17900 24668
rect 17807 24628 17900 24656
rect 17894 24616 17900 24628
rect 17952 24656 17958 24668
rect 18722 24656 18728 24668
rect 17952 24628 18728 24656
rect 17952 24616 17958 24628
rect 18722 24616 18728 24628
rect 18780 24656 18786 24668
rect 19366 24656 19372 24668
rect 18780 24628 19372 24656
rect 18780 24616 18786 24628
rect 19366 24616 19372 24628
rect 19424 24616 19430 24668
rect 20930 24656 20936 24668
rect 20891 24628 20936 24656
rect 20930 24616 20936 24628
rect 20988 24616 20994 24668
rect 25898 24656 25904 24668
rect 25859 24628 25904 24656
rect 25898 24616 25904 24628
rect 25956 24616 25962 24668
rect 26266 24616 26272 24668
rect 26324 24656 26330 24668
rect 27189 24659 27247 24665
rect 27189 24656 27201 24659
rect 26324 24628 27201 24656
rect 26324 24616 26330 24628
rect 27189 24625 27201 24628
rect 27235 24656 27247 24659
rect 27370 24656 27376 24668
rect 27235 24628 27376 24656
rect 27235 24625 27247 24628
rect 27189 24619 27247 24625
rect 27370 24616 27376 24628
rect 27428 24616 27434 24668
rect 27554 24656 27560 24668
rect 27515 24628 27560 24656
rect 27554 24616 27560 24628
rect 27612 24616 27618 24668
rect 28198 24656 28204 24668
rect 28159 24628 28204 24656
rect 28198 24616 28204 24628
rect 28256 24616 28262 24668
rect 29581 24659 29639 24665
rect 29581 24625 29593 24659
rect 29627 24656 29639 24659
rect 29854 24656 29860 24668
rect 29627 24628 29860 24656
rect 29627 24625 29639 24628
rect 29581 24619 29639 24625
rect 29854 24616 29860 24628
rect 29912 24616 29918 24668
rect 4554 24588 4560 24600
rect 4467 24560 4560 24588
rect 4554 24548 4560 24560
rect 4612 24588 4618 24600
rect 6210 24588 6216 24600
rect 4612 24560 6216 24588
rect 4612 24548 4618 24560
rect 6210 24548 6216 24560
rect 6268 24548 6274 24600
rect 7041 24591 7099 24597
rect 7041 24557 7053 24591
rect 7087 24588 7099 24591
rect 7682 24588 7688 24600
rect 7087 24560 7688 24588
rect 7087 24557 7099 24560
rect 7041 24551 7099 24557
rect 7682 24548 7688 24560
rect 7740 24588 7746 24600
rect 7777 24591 7835 24597
rect 7777 24588 7789 24591
rect 7740 24560 7789 24588
rect 7740 24548 7746 24560
rect 7777 24557 7789 24560
rect 7823 24557 7835 24591
rect 7777 24551 7835 24557
rect 16054 24548 16060 24600
rect 16112 24588 16118 24600
rect 16149 24591 16207 24597
rect 16149 24588 16161 24591
rect 16112 24560 16161 24588
rect 16112 24548 16118 24560
rect 16149 24557 16161 24560
rect 16195 24588 16207 24591
rect 17069 24591 17127 24597
rect 17069 24588 17081 24591
rect 16195 24560 17081 24588
rect 16195 24557 16207 24560
rect 16149 24551 16207 24557
rect 17069 24557 17081 24560
rect 17115 24588 17127 24591
rect 17710 24588 17716 24600
rect 17115 24560 17716 24588
rect 17115 24557 17127 24560
rect 17069 24551 17127 24557
rect 17710 24548 17716 24560
rect 17768 24548 17774 24600
rect 17986 24588 17992 24600
rect 17947 24560 17992 24588
rect 17986 24548 17992 24560
rect 18044 24548 18050 24600
rect 21206 24588 21212 24600
rect 21167 24560 21212 24588
rect 21206 24548 21212 24560
rect 21264 24548 21270 24600
rect 22954 24588 22960 24600
rect 22915 24560 22960 24588
rect 22954 24548 22960 24560
rect 23012 24548 23018 24600
rect 28477 24591 28535 24597
rect 28477 24557 28489 24591
rect 28523 24588 28535 24591
rect 29210 24588 29216 24600
rect 28523 24560 29216 24588
rect 28523 24557 28535 24560
rect 28477 24551 28535 24557
rect 29210 24548 29216 24560
rect 29268 24548 29274 24600
rect 29762 24588 29768 24600
rect 29723 24560 29768 24588
rect 29762 24548 29768 24560
rect 29820 24548 29826 24600
rect 28382 24520 28388 24532
rect 28343 24492 28388 24520
rect 28382 24480 28388 24492
rect 28440 24480 28446 24532
rect 2165 24455 2223 24461
rect 2165 24421 2177 24455
rect 2211 24452 2223 24455
rect 3082 24452 3088 24464
rect 2211 24424 3088 24452
rect 2211 24421 2223 24424
rect 2165 24415 2223 24421
rect 3082 24412 3088 24424
rect 3140 24412 3146 24464
rect 9522 24452 9528 24464
rect 9483 24424 9528 24452
rect 9522 24412 9528 24424
rect 9580 24412 9586 24464
rect 13297 24455 13355 24461
rect 13297 24421 13309 24455
rect 13343 24452 13355 24455
rect 13938 24452 13944 24464
rect 13343 24424 13944 24452
rect 13343 24421 13355 24424
rect 13297 24415 13355 24421
rect 13938 24412 13944 24424
rect 13996 24412 14002 24464
rect 18446 24452 18452 24464
rect 18359 24424 18452 24452
rect 18446 24412 18452 24424
rect 18504 24452 18510 24464
rect 21574 24452 21580 24464
rect 18504 24424 21580 24452
rect 18504 24412 18510 24424
rect 21574 24412 21580 24424
rect 21632 24412 21638 24464
rect 23414 24412 23420 24464
rect 23472 24452 23478 24464
rect 23601 24455 23659 24461
rect 23601 24452 23613 24455
rect 23472 24424 23613 24452
rect 23472 24412 23478 24424
rect 23601 24421 23613 24424
rect 23647 24452 23659 24455
rect 23693 24455 23751 24461
rect 23693 24452 23705 24455
rect 23647 24424 23705 24452
rect 23647 24421 23659 24424
rect 23601 24415 23659 24421
rect 23693 24421 23705 24424
rect 23739 24421 23751 24455
rect 23693 24415 23751 24421
rect 400 24362 31680 24384
rect 400 24310 3510 24362
rect 3562 24310 3574 24362
rect 3626 24310 3638 24362
rect 3690 24310 3702 24362
rect 3754 24310 3766 24362
rect 3818 24310 31680 24362
rect 400 24288 31680 24310
rect 3910 24208 3916 24260
rect 3968 24248 3974 24260
rect 4189 24251 4247 24257
rect 4189 24248 4201 24251
rect 3968 24220 4201 24248
rect 3968 24208 3974 24220
rect 4189 24217 4201 24220
rect 4235 24217 4247 24251
rect 4189 24211 4247 24217
rect 9062 24208 9068 24260
rect 9120 24248 9126 24260
rect 9522 24248 9528 24260
rect 9120 24220 9528 24248
rect 9120 24208 9126 24220
rect 9522 24208 9528 24220
rect 9580 24208 9586 24260
rect 10442 24248 10448 24260
rect 10403 24220 10448 24248
rect 10442 24208 10448 24220
rect 10500 24208 10506 24260
rect 12377 24251 12435 24257
rect 12377 24217 12389 24251
rect 12423 24248 12435 24251
rect 12558 24248 12564 24260
rect 12423 24220 12564 24248
rect 12423 24217 12435 24220
rect 12377 24211 12435 24217
rect 966 24140 972 24192
rect 1024 24180 1030 24192
rect 1981 24183 2039 24189
rect 1981 24180 1993 24183
rect 1024 24152 1993 24180
rect 1024 24140 1030 24152
rect 1981 24149 1993 24152
rect 2027 24180 2039 24183
rect 2441 24183 2499 24189
rect 2441 24180 2453 24183
rect 2027 24152 2453 24180
rect 2027 24149 2039 24152
rect 1981 24143 2039 24149
rect 2441 24149 2453 24152
rect 2487 24149 2499 24183
rect 2441 24143 2499 24149
rect 3729 24183 3787 24189
rect 3729 24149 3741 24183
rect 3775 24180 3787 24183
rect 4554 24180 4560 24192
rect 3775 24152 4560 24180
rect 3775 24149 3787 24152
rect 3729 24143 3787 24149
rect 4554 24140 4560 24152
rect 4612 24140 4618 24192
rect 1797 24115 1855 24121
rect 1797 24081 1809 24115
rect 1843 24112 1855 24115
rect 2993 24115 3051 24121
rect 2993 24112 3005 24115
rect 1843 24084 3005 24112
rect 1843 24081 1855 24084
rect 1797 24075 1855 24081
rect 2993 24081 3005 24084
rect 3039 24112 3051 24115
rect 3913 24115 3971 24121
rect 3039 24084 3220 24112
rect 3039 24081 3051 24084
rect 2993 24075 3051 24081
rect 2625 24047 2683 24053
rect 2625 24013 2637 24047
rect 2671 24013 2683 24047
rect 2625 24007 2683 24013
rect 1613 23979 1671 23985
rect 1613 23945 1625 23979
rect 1659 23976 1671 23979
rect 2640 23976 2668 24007
rect 2714 24004 2720 24056
rect 2772 24044 2778 24056
rect 3082 24044 3088 24056
rect 2772 24016 2817 24044
rect 3043 24016 3088 24044
rect 2772 24004 2778 24016
rect 3082 24004 3088 24016
rect 3140 24004 3146 24056
rect 3192 24044 3220 24084
rect 3913 24081 3925 24115
rect 3959 24112 3971 24115
rect 4646 24112 4652 24124
rect 3959 24084 4652 24112
rect 3959 24081 3971 24084
rect 3913 24075 3971 24081
rect 4646 24072 4652 24084
rect 4704 24072 4710 24124
rect 6857 24115 6915 24121
rect 6857 24081 6869 24115
rect 6903 24112 6915 24115
rect 8973 24115 9031 24121
rect 8973 24112 8985 24115
rect 6903 24084 8985 24112
rect 6903 24081 6915 24084
rect 6857 24075 6915 24081
rect 8973 24081 8985 24084
rect 9019 24112 9031 24115
rect 9246 24112 9252 24124
rect 9019 24084 9252 24112
rect 9019 24081 9031 24084
rect 8973 24075 9031 24081
rect 9246 24072 9252 24084
rect 9304 24072 9310 24124
rect 9614 24072 9620 24124
rect 9672 24112 9678 24124
rect 9985 24115 10043 24121
rect 9985 24112 9997 24115
rect 9672 24084 9997 24112
rect 9672 24072 9678 24084
rect 9985 24081 9997 24084
rect 10031 24112 10043 24115
rect 10629 24115 10687 24121
rect 10629 24112 10641 24115
rect 10031 24084 10641 24112
rect 10031 24081 10043 24084
rect 9985 24075 10043 24081
rect 10629 24081 10641 24084
rect 10675 24081 10687 24115
rect 10629 24075 10687 24081
rect 4738 24044 4744 24056
rect 3192 24016 4744 24044
rect 4738 24004 4744 24016
rect 4796 24044 4802 24056
rect 5750 24044 5756 24056
rect 4796 24016 5756 24044
rect 4796 24004 4802 24016
rect 5750 24004 5756 24016
rect 5808 24004 5814 24056
rect 6302 24004 6308 24056
rect 6360 24044 6366 24056
rect 6489 24047 6547 24053
rect 6489 24044 6501 24047
rect 6360 24016 6501 24044
rect 6360 24004 6366 24016
rect 6489 24013 6501 24016
rect 6535 24044 6547 24047
rect 6946 24044 6952 24056
rect 6535 24016 6952 24044
rect 6535 24013 6547 24016
rect 6489 24007 6547 24013
rect 6946 24004 6952 24016
rect 7004 24004 7010 24056
rect 9801 24047 9859 24053
rect 9801 24013 9813 24047
rect 9847 24044 9859 24047
rect 10442 24044 10448 24056
rect 9847 24016 10448 24044
rect 9847 24013 9859 24016
rect 9801 24007 9859 24013
rect 10442 24004 10448 24016
rect 10500 24044 10506 24056
rect 11270 24044 11276 24056
rect 10500 24016 11276 24044
rect 10500 24004 10506 24016
rect 11270 24004 11276 24016
rect 11328 24004 11334 24056
rect 11733 24047 11791 24053
rect 11733 24013 11745 24047
rect 11779 24044 11791 24047
rect 11914 24044 11920 24056
rect 11779 24016 11920 24044
rect 11779 24013 11791 24016
rect 11733 24007 11791 24013
rect 11914 24004 11920 24016
rect 11972 24044 11978 24056
rect 12392 24044 12420 24211
rect 12558 24208 12564 24220
rect 12616 24208 12622 24260
rect 15689 24251 15747 24257
rect 15689 24217 15701 24251
rect 15735 24248 15747 24251
rect 15778 24248 15784 24260
rect 15735 24220 15784 24248
rect 15735 24217 15747 24220
rect 15689 24211 15747 24217
rect 15778 24208 15784 24220
rect 15836 24208 15842 24260
rect 16054 24248 16060 24260
rect 16015 24220 16060 24248
rect 16054 24208 16060 24220
rect 16112 24208 16118 24260
rect 16974 24208 16980 24260
rect 17032 24248 17038 24260
rect 17345 24251 17403 24257
rect 17345 24248 17357 24251
rect 17032 24220 17357 24248
rect 17032 24208 17038 24220
rect 17345 24217 17357 24220
rect 17391 24217 17403 24251
rect 17710 24248 17716 24260
rect 17671 24220 17716 24248
rect 17345 24211 17403 24217
rect 17710 24208 17716 24220
rect 17768 24208 17774 24260
rect 20930 24208 20936 24260
rect 20988 24248 20994 24260
rect 21301 24251 21359 24257
rect 21301 24248 21313 24251
rect 20988 24220 21313 24248
rect 20988 24208 20994 24220
rect 21301 24217 21313 24220
rect 21347 24217 21359 24251
rect 21301 24211 21359 24217
rect 21577 24251 21635 24257
rect 21577 24217 21589 24251
rect 21623 24248 21635 24251
rect 21666 24248 21672 24260
rect 21623 24220 21672 24248
rect 21623 24217 21635 24220
rect 21577 24211 21635 24217
rect 21666 24208 21672 24220
rect 21724 24208 21730 24260
rect 25898 24248 25904 24260
rect 25859 24220 25904 24248
rect 25898 24208 25904 24220
rect 25956 24208 25962 24260
rect 26085 24251 26143 24257
rect 26085 24217 26097 24251
rect 26131 24248 26143 24251
rect 26174 24248 26180 24260
rect 26131 24220 26180 24248
rect 26131 24217 26143 24220
rect 26085 24211 26143 24217
rect 26174 24208 26180 24220
rect 26232 24208 26238 24260
rect 27370 24248 27376 24260
rect 27331 24220 27376 24248
rect 27370 24208 27376 24220
rect 27428 24208 27434 24260
rect 27922 24208 27928 24260
rect 27980 24248 27986 24260
rect 28017 24251 28075 24257
rect 28017 24248 28029 24251
rect 27980 24220 28029 24248
rect 27980 24208 27986 24220
rect 28017 24217 28029 24220
rect 28063 24248 28075 24251
rect 28198 24248 28204 24260
rect 28063 24220 28204 24248
rect 28063 24217 28075 24220
rect 28017 24211 28075 24217
rect 28198 24208 28204 24220
rect 28256 24208 28262 24260
rect 29302 24208 29308 24260
rect 29360 24248 29366 24260
rect 29762 24248 29768 24260
rect 29360 24220 29768 24248
rect 29360 24208 29366 24220
rect 29762 24208 29768 24220
rect 29820 24208 29826 24260
rect 29854 24208 29860 24260
rect 29912 24248 29918 24260
rect 29912 24220 29957 24248
rect 29912 24208 29918 24220
rect 17066 24180 17072 24192
rect 17027 24152 17072 24180
rect 17066 24140 17072 24152
rect 17124 24140 17130 24192
rect 17621 24183 17679 24189
rect 17621 24149 17633 24183
rect 17667 24180 17679 24183
rect 17986 24180 17992 24192
rect 17667 24152 17992 24180
rect 17667 24149 17679 24152
rect 17621 24143 17679 24149
rect 13938 24072 13944 24124
rect 13996 24112 14002 24124
rect 13996 24084 15548 24112
rect 13996 24072 14002 24084
rect 13202 24044 13208 24056
rect 11972 24016 12420 24044
rect 13163 24016 13208 24044
rect 11972 24004 11978 24016
rect 13202 24004 13208 24016
rect 13260 24004 13266 24056
rect 15520 24044 15548 24084
rect 15594 24072 15600 24124
rect 15652 24112 15658 24124
rect 15873 24115 15931 24121
rect 15873 24112 15885 24115
rect 15652 24084 15885 24112
rect 15652 24072 15658 24084
rect 15873 24081 15885 24084
rect 15919 24112 15931 24115
rect 17636 24112 17664 24143
rect 17986 24140 17992 24152
rect 18044 24140 18050 24192
rect 21025 24183 21083 24189
rect 21025 24149 21037 24183
rect 21071 24180 21083 24183
rect 22954 24180 22960 24192
rect 21071 24152 22960 24180
rect 21071 24149 21083 24152
rect 21025 24143 21083 24149
rect 22954 24140 22960 24152
rect 23012 24140 23018 24192
rect 27281 24183 27339 24189
rect 27281 24149 27293 24183
rect 27327 24180 27339 24183
rect 28382 24180 28388 24192
rect 27327 24152 28388 24180
rect 27327 24149 27339 24152
rect 27281 24143 27339 24149
rect 28382 24140 28388 24152
rect 28440 24140 28446 24192
rect 29397 24183 29455 24189
rect 29397 24180 29409 24183
rect 28860 24152 29409 24180
rect 15919 24084 17664 24112
rect 15919 24081 15931 24084
rect 15873 24075 15931 24081
rect 19277 24047 19335 24053
rect 19277 24044 19289 24047
rect 15520 24016 19289 24044
rect 19277 24013 19289 24016
rect 19323 24044 19335 24047
rect 19829 24047 19887 24053
rect 19829 24044 19841 24047
rect 19323 24016 19841 24044
rect 19323 24013 19335 24016
rect 19277 24007 19335 24013
rect 19829 24013 19841 24016
rect 19875 24044 19887 24047
rect 20286 24044 20292 24056
rect 19875 24016 20292 24044
rect 19875 24013 19887 24016
rect 19829 24007 19887 24013
rect 20286 24004 20292 24016
rect 20344 24004 20350 24056
rect 27370 24004 27376 24056
rect 27428 24044 27434 24056
rect 28474 24044 28480 24056
rect 27428 24016 28480 24044
rect 27428 24004 27434 24016
rect 28474 24004 28480 24016
rect 28532 24044 28538 24056
rect 28860 24053 28888 24152
rect 29397 24149 29409 24152
rect 29443 24180 29455 24183
rect 30590 24180 30596 24192
rect 29443 24152 30596 24180
rect 29443 24149 29455 24152
rect 29397 24143 29455 24149
rect 30590 24140 30596 24152
rect 30648 24140 30654 24192
rect 29762 24072 29768 24124
rect 29820 24112 29826 24124
rect 31510 24112 31516 24124
rect 29820 24084 31516 24112
rect 29820 24072 29826 24084
rect 31510 24072 31516 24084
rect 31568 24072 31574 24124
rect 28845 24047 28903 24053
rect 28845 24044 28857 24047
rect 28532 24016 28857 24044
rect 28532 24004 28538 24016
rect 28845 24013 28857 24016
rect 28891 24013 28903 24047
rect 29210 24044 29216 24056
rect 29123 24016 29216 24044
rect 28845 24007 28903 24013
rect 29210 24004 29216 24016
rect 29268 24044 29274 24056
rect 29489 24047 29547 24053
rect 29489 24044 29501 24047
rect 29268 24016 29501 24044
rect 29268 24004 29274 24016
rect 29489 24013 29501 24016
rect 29535 24013 29547 24047
rect 29489 24007 29547 24013
rect 3910 23976 3916 23988
rect 1659 23948 3916 23976
rect 1659 23945 1671 23948
rect 1613 23939 1671 23945
rect 3910 23936 3916 23948
rect 3968 23936 3974 23988
rect 6578 23936 6584 23988
rect 6636 23976 6642 23988
rect 6673 23979 6731 23985
rect 6673 23976 6685 23979
rect 6636 23948 6685 23976
rect 6636 23936 6642 23948
rect 6673 23945 6685 23948
rect 6719 23976 6731 23979
rect 7225 23979 7283 23985
rect 7225 23976 7237 23979
rect 6719 23948 7237 23976
rect 6719 23945 6731 23948
rect 6673 23939 6731 23945
rect 7225 23945 7237 23948
rect 7271 23945 7283 23979
rect 7225 23939 7283 23945
rect 7682 23936 7688 23988
rect 7740 23936 7746 23988
rect 12006 23976 12012 23988
rect 11967 23948 12012 23976
rect 12006 23936 12012 23948
rect 12064 23936 12070 23988
rect 12098 23936 12104 23988
rect 12156 23976 12162 23988
rect 12929 23979 12987 23985
rect 12929 23976 12941 23979
rect 12156 23948 12941 23976
rect 12156 23936 12162 23948
rect 12929 23945 12941 23948
rect 12975 23976 12987 23979
rect 13481 23979 13539 23985
rect 13481 23976 13493 23979
rect 12975 23948 13493 23976
rect 12975 23945 12987 23948
rect 12929 23939 12987 23945
rect 13481 23945 13493 23948
rect 13527 23945 13539 23979
rect 13481 23939 13539 23945
rect 13938 23936 13944 23988
rect 13996 23936 14002 23988
rect 15229 23979 15287 23985
rect 15229 23976 15241 23979
rect 15152 23948 15241 23976
rect 4097 23911 4155 23917
rect 4097 23877 4109 23911
rect 4143 23908 4155 23911
rect 4278 23908 4284 23920
rect 4143 23880 4284 23908
rect 4143 23877 4155 23880
rect 4097 23871 4155 23877
rect 4278 23868 4284 23880
rect 4336 23868 4342 23920
rect 12558 23908 12564 23920
rect 12519 23880 12564 23908
rect 12558 23868 12564 23880
rect 12616 23868 12622 23920
rect 12650 23868 12656 23920
rect 12708 23908 12714 23920
rect 13113 23911 13171 23917
rect 13113 23908 13125 23911
rect 12708 23880 13125 23908
rect 12708 23868 12714 23880
rect 13113 23877 13125 23880
rect 13159 23908 13171 23911
rect 15152 23908 15180 23948
rect 15229 23945 15241 23948
rect 15275 23945 15287 23979
rect 15229 23939 15287 23945
rect 19366 23936 19372 23988
rect 19424 23976 19430 23988
rect 19553 23979 19611 23985
rect 19553 23976 19565 23979
rect 19424 23948 19565 23976
rect 19424 23936 19430 23948
rect 19553 23945 19565 23948
rect 19599 23945 19611 23979
rect 21206 23976 21212 23988
rect 21119 23948 21212 23976
rect 19553 23939 19611 23945
rect 21206 23936 21212 23948
rect 21264 23976 21270 23988
rect 21942 23976 21948 23988
rect 21264 23948 21948 23976
rect 21264 23936 21270 23948
rect 21942 23936 21948 23948
rect 22000 23936 22006 23988
rect 25898 23936 25904 23988
rect 25956 23976 25962 23988
rect 27554 23976 27560 23988
rect 25956 23948 27560 23976
rect 25956 23936 25962 23948
rect 27554 23936 27560 23948
rect 27612 23936 27618 23988
rect 27833 23979 27891 23985
rect 27833 23945 27845 23979
rect 27879 23976 27891 23979
rect 29228 23976 29256 24004
rect 27879 23948 29256 23976
rect 27879 23945 27891 23948
rect 27833 23939 27891 23945
rect 20010 23908 20016 23920
rect 13159 23880 15180 23908
rect 19971 23880 20016 23908
rect 13159 23877 13171 23880
rect 13113 23871 13171 23877
rect 20010 23868 20016 23880
rect 20068 23868 20074 23920
rect 400 23818 31680 23840
rect 400 23766 18870 23818
rect 18922 23766 18934 23818
rect 18986 23766 18998 23818
rect 19050 23766 19062 23818
rect 19114 23766 19126 23818
rect 19178 23766 31680 23818
rect 400 23744 31680 23766
rect 2165 23707 2223 23713
rect 2165 23673 2177 23707
rect 2211 23704 2223 23707
rect 2622 23704 2628 23716
rect 2211 23676 2628 23704
rect 2211 23673 2223 23676
rect 2165 23667 2223 23673
rect 2622 23664 2628 23676
rect 2680 23664 2686 23716
rect 7682 23704 7688 23716
rect 7643 23676 7688 23704
rect 7682 23664 7688 23676
rect 7740 23664 7746 23716
rect 7774 23664 7780 23716
rect 7832 23704 7838 23716
rect 9982 23704 9988 23716
rect 7832 23676 9988 23704
rect 7832 23664 7838 23676
rect 9982 23664 9988 23676
rect 10040 23664 10046 23716
rect 13202 23704 13208 23716
rect 13163 23676 13208 23704
rect 13202 23664 13208 23676
rect 13260 23664 13266 23716
rect 19366 23664 19372 23716
rect 19424 23704 19430 23716
rect 20010 23704 20016 23716
rect 19424 23676 20016 23704
rect 19424 23664 19430 23676
rect 20010 23664 20016 23676
rect 20068 23664 20074 23716
rect 24242 23704 24248 23716
rect 24203 23676 24248 23704
rect 24242 23664 24248 23676
rect 24300 23664 24306 23716
rect 29581 23639 29639 23645
rect 29581 23605 29593 23639
rect 29627 23636 29639 23639
rect 30222 23636 30228 23648
rect 29627 23608 30228 23636
rect 29627 23605 29639 23608
rect 29581 23599 29639 23605
rect 30222 23596 30228 23608
rect 30280 23596 30286 23648
rect 1150 23568 1156 23580
rect 1063 23540 1156 23568
rect 1150 23528 1156 23540
rect 1208 23568 1214 23580
rect 1334 23568 1340 23580
rect 1208 23540 1340 23568
rect 1208 23528 1214 23540
rect 1334 23528 1340 23540
rect 1392 23528 1398 23580
rect 3358 23568 3364 23580
rect 3319 23540 3364 23568
rect 3358 23528 3364 23540
rect 3416 23528 3422 23580
rect 6857 23571 6915 23577
rect 6857 23537 6869 23571
rect 6903 23568 6915 23571
rect 7130 23568 7136 23580
rect 6903 23540 7136 23568
rect 6903 23537 6915 23540
rect 6857 23531 6915 23537
rect 7130 23528 7136 23540
rect 7188 23528 7194 23580
rect 9062 23568 9068 23580
rect 9023 23540 9068 23568
rect 9062 23528 9068 23540
rect 9120 23528 9126 23580
rect 11086 23568 11092 23580
rect 11047 23540 11092 23568
rect 11086 23528 11092 23540
rect 11144 23528 11150 23580
rect 11178 23528 11184 23580
rect 11236 23568 11242 23580
rect 11549 23571 11607 23577
rect 11549 23568 11561 23571
rect 11236 23540 11561 23568
rect 11236 23528 11242 23540
rect 11549 23537 11561 23540
rect 11595 23537 11607 23571
rect 11549 23531 11607 23537
rect 18633 23571 18691 23577
rect 18633 23537 18645 23571
rect 18679 23568 18691 23571
rect 18722 23568 18728 23580
rect 18679 23540 18728 23568
rect 18679 23537 18691 23540
rect 18633 23531 18691 23537
rect 18722 23528 18728 23540
rect 18780 23528 18786 23580
rect 21574 23568 21580 23580
rect 21535 23540 21580 23568
rect 21574 23528 21580 23540
rect 21632 23528 21638 23580
rect 22954 23568 22960 23580
rect 22915 23540 22960 23568
rect 22954 23528 22960 23540
rect 23012 23528 23018 23580
rect 23141 23571 23199 23577
rect 23141 23537 23153 23571
rect 23187 23537 23199 23571
rect 23141 23531 23199 23537
rect 969 23503 1027 23509
rect 969 23469 981 23503
rect 1015 23500 1027 23503
rect 1426 23500 1432 23512
rect 1015 23472 1432 23500
rect 1015 23469 1027 23472
rect 969 23463 1027 23469
rect 1426 23460 1432 23472
rect 1484 23460 1490 23512
rect 7038 23500 7044 23512
rect 6999 23472 7044 23500
rect 7038 23460 7044 23472
rect 7096 23460 7102 23512
rect 9341 23503 9399 23509
rect 9341 23469 9353 23503
rect 9387 23500 9399 23503
rect 9522 23500 9528 23512
rect 9387 23472 9528 23500
rect 9387 23469 9399 23472
rect 9341 23463 9399 23469
rect 9522 23460 9528 23472
rect 9580 23460 9586 23512
rect 10902 23500 10908 23512
rect 10863 23472 10908 23500
rect 10902 23460 10908 23472
rect 10960 23460 10966 23512
rect 11454 23500 11460 23512
rect 11415 23472 11460 23500
rect 11454 23460 11460 23472
rect 11512 23460 11518 23512
rect 18262 23460 18268 23512
rect 18320 23500 18326 23512
rect 18541 23503 18599 23509
rect 18541 23500 18553 23503
rect 18320 23472 18553 23500
rect 18320 23460 18326 23472
rect 18541 23469 18553 23472
rect 18587 23469 18599 23503
rect 18541 23463 18599 23469
rect 22862 23460 22868 23512
rect 22920 23500 22926 23512
rect 23156 23500 23184 23531
rect 26910 23528 26916 23580
rect 26968 23568 26974 23580
rect 27278 23568 27284 23580
rect 26968 23540 27284 23568
rect 26968 23528 26974 23540
rect 27278 23528 27284 23540
rect 27336 23568 27342 23580
rect 27373 23571 27431 23577
rect 27373 23568 27385 23571
rect 27336 23540 27385 23568
rect 27336 23528 27342 23540
rect 27373 23537 27385 23540
rect 27419 23537 27431 23571
rect 27554 23568 27560 23580
rect 27515 23540 27560 23568
rect 27373 23531 27431 23537
rect 27554 23528 27560 23540
rect 27612 23528 27618 23580
rect 28293 23571 28351 23577
rect 28293 23537 28305 23571
rect 28339 23537 28351 23571
rect 28474 23568 28480 23580
rect 28435 23540 28480 23568
rect 28293 23531 28351 23537
rect 22920 23472 23184 23500
rect 22920 23460 22926 23472
rect 27462 23460 27468 23512
rect 27520 23500 27526 23512
rect 28308 23500 28336 23531
rect 28474 23528 28480 23540
rect 28532 23528 28538 23580
rect 29765 23571 29823 23577
rect 29765 23537 29777 23571
rect 29811 23568 29823 23571
rect 30038 23568 30044 23580
rect 29811 23540 30044 23568
rect 29811 23537 29823 23540
rect 29765 23531 29823 23537
rect 30038 23528 30044 23540
rect 30096 23528 30102 23580
rect 30133 23503 30191 23509
rect 30133 23500 30145 23503
rect 27520 23472 30145 23500
rect 27520 23460 27526 23472
rect 30133 23469 30145 23472
rect 30179 23500 30191 23503
rect 30406 23500 30412 23512
rect 30179 23472 30412 23500
rect 30179 23469 30191 23472
rect 30133 23463 30191 23469
rect 30406 23460 30412 23472
rect 30464 23460 30470 23512
rect 11917 23435 11975 23441
rect 11917 23401 11929 23435
rect 11963 23432 11975 23435
rect 12098 23432 12104 23444
rect 11963 23404 12104 23432
rect 11963 23401 11975 23404
rect 11917 23395 11975 23401
rect 12098 23392 12104 23404
rect 12156 23392 12162 23444
rect 12285 23435 12343 23441
rect 12285 23401 12297 23435
rect 12331 23432 12343 23435
rect 12834 23432 12840 23444
rect 12331 23404 12840 23432
rect 12331 23401 12343 23404
rect 12285 23395 12343 23401
rect 12834 23392 12840 23404
rect 12892 23392 12898 23444
rect 26821 23435 26879 23441
rect 26821 23401 26833 23435
rect 26867 23432 26879 23435
rect 27002 23432 27008 23444
rect 26867 23404 27008 23432
rect 26867 23401 26879 23404
rect 26821 23395 26879 23401
rect 27002 23392 27008 23404
rect 27060 23392 27066 23444
rect 27186 23432 27192 23444
rect 27147 23404 27192 23432
rect 27186 23392 27192 23404
rect 27244 23392 27250 23444
rect 785 23367 843 23373
rect 785 23333 797 23367
rect 831 23364 843 23367
rect 1978 23364 1984 23376
rect 831 23336 1984 23364
rect 831 23333 843 23336
rect 785 23327 843 23333
rect 1978 23324 1984 23336
rect 2036 23324 2042 23376
rect 3082 23324 3088 23376
rect 3140 23364 3146 23376
rect 3637 23367 3695 23373
rect 3637 23364 3649 23367
rect 3140 23336 3649 23364
rect 3140 23324 3146 23336
rect 3637 23333 3649 23336
rect 3683 23364 3695 23367
rect 4002 23364 4008 23376
rect 3683 23336 4008 23364
rect 3683 23333 3695 23336
rect 3637 23327 3695 23333
rect 4002 23324 4008 23336
rect 4060 23324 4066 23376
rect 6213 23367 6271 23373
rect 6213 23333 6225 23367
rect 6259 23364 6271 23367
rect 7314 23364 7320 23376
rect 6259 23336 7320 23364
rect 6259 23333 6271 23336
rect 6213 23327 6271 23333
rect 7314 23324 7320 23336
rect 7372 23324 7378 23376
rect 12374 23364 12380 23376
rect 12335 23336 12380 23364
rect 12374 23324 12380 23336
rect 12432 23324 12438 23376
rect 17986 23324 17992 23376
rect 18044 23364 18050 23376
rect 18817 23367 18875 23373
rect 18817 23364 18829 23367
rect 18044 23336 18829 23364
rect 18044 23324 18050 23336
rect 18817 23333 18829 23336
rect 18863 23364 18875 23367
rect 21482 23364 21488 23376
rect 18863 23336 21488 23364
rect 18863 23333 18875 23336
rect 18817 23327 18875 23333
rect 21482 23324 21488 23336
rect 21540 23324 21546 23376
rect 21666 23364 21672 23376
rect 21627 23336 21672 23364
rect 21666 23324 21672 23336
rect 21724 23324 21730 23376
rect 23138 23324 23144 23376
rect 23196 23364 23202 23376
rect 23233 23367 23291 23373
rect 23233 23364 23245 23367
rect 23196 23336 23245 23364
rect 23196 23324 23202 23336
rect 23233 23333 23245 23336
rect 23279 23333 23291 23367
rect 23233 23327 23291 23333
rect 24061 23367 24119 23373
rect 24061 23333 24073 23367
rect 24107 23364 24119 23367
rect 24794 23364 24800 23376
rect 24107 23336 24800 23364
rect 24107 23333 24119 23336
rect 24061 23327 24119 23333
rect 24794 23324 24800 23336
rect 24852 23324 24858 23376
rect 400 23274 31680 23296
rect 400 23222 3510 23274
rect 3562 23222 3574 23274
rect 3626 23222 3638 23274
rect 3690 23222 3702 23274
rect 3754 23222 3766 23274
rect 3818 23222 31680 23274
rect 400 23200 31680 23222
rect 3085 23163 3143 23169
rect 3085 23129 3097 23163
rect 3131 23160 3143 23163
rect 3821 23163 3879 23169
rect 3821 23160 3833 23163
rect 3131 23132 3833 23160
rect 3131 23129 3143 23132
rect 3085 23123 3143 23129
rect 3821 23129 3833 23132
rect 3867 23160 3879 23163
rect 4554 23160 4560 23172
rect 3867 23132 4560 23160
rect 3867 23129 3879 23132
rect 3821 23123 3879 23129
rect 4554 23120 4560 23132
rect 4612 23120 4618 23172
rect 5750 23160 5756 23172
rect 5711 23132 5756 23160
rect 5750 23120 5756 23132
rect 5808 23160 5814 23172
rect 5808 23132 7084 23160
rect 5808 23120 5814 23132
rect 5937 23095 5995 23101
rect 5937 23061 5949 23095
rect 5983 23092 5995 23095
rect 6489 23095 6547 23101
rect 6489 23092 6501 23095
rect 5983 23064 6501 23092
rect 5983 23061 5995 23064
rect 5937 23055 5995 23061
rect 6489 23061 6501 23064
rect 6535 23092 6547 23095
rect 6578 23092 6584 23104
rect 6535 23064 6584 23092
rect 6535 23061 6547 23064
rect 6489 23055 6547 23061
rect 6578 23052 6584 23064
rect 6636 23052 6642 23104
rect 7056 23092 7084 23132
rect 7130 23120 7136 23172
rect 7188 23160 7194 23172
rect 7685 23163 7743 23169
rect 7685 23160 7697 23163
rect 7188 23132 7697 23160
rect 7188 23120 7194 23132
rect 7685 23129 7697 23132
rect 7731 23160 7743 23163
rect 7866 23160 7872 23172
rect 7731 23132 7872 23160
rect 7731 23129 7743 23132
rect 7685 23123 7743 23129
rect 7866 23120 7872 23132
rect 7924 23160 7930 23172
rect 10258 23160 10264 23172
rect 7924 23132 10264 23160
rect 7924 23120 7930 23132
rect 10258 23120 10264 23132
rect 10316 23120 10322 23172
rect 10629 23163 10687 23169
rect 10629 23129 10641 23163
rect 10675 23160 10687 23163
rect 12098 23160 12104 23172
rect 10675 23132 12104 23160
rect 10675 23129 10687 23132
rect 10629 23123 10687 23129
rect 12098 23120 12104 23132
rect 12156 23120 12162 23172
rect 12374 23120 12380 23172
rect 12432 23160 12438 23172
rect 12469 23163 12527 23169
rect 12469 23160 12481 23163
rect 12432 23132 12481 23160
rect 12432 23120 12438 23132
rect 12469 23129 12481 23132
rect 12515 23129 12527 23163
rect 12469 23123 12527 23129
rect 13202 23120 13208 23172
rect 13260 23160 13266 23172
rect 14950 23160 14956 23172
rect 13260 23132 14214 23160
rect 14911 23132 14956 23160
rect 13260 23120 13266 23132
rect 11273 23095 11331 23101
rect 11273 23092 11285 23095
rect 7056 23064 11285 23092
rect 966 23024 972 23036
rect 927 22996 972 23024
rect 966 22984 972 22996
rect 1024 22984 1030 23036
rect 1978 22984 1984 23036
rect 2036 23024 2042 23036
rect 2717 23027 2775 23033
rect 2717 23024 2729 23027
rect 2036 22996 2729 23024
rect 2036 22984 2042 22996
rect 2717 22993 2729 22996
rect 2763 23024 2775 23027
rect 3358 23024 3364 23036
rect 2763 22996 3364 23024
rect 2763 22993 2775 22996
rect 2717 22987 2775 22993
rect 3358 22984 3364 22996
rect 3416 23024 3422 23036
rect 4189 23027 4247 23033
rect 4189 23024 4201 23027
rect 3416 22996 4201 23024
rect 3416 22984 3422 22996
rect 690 22956 696 22968
rect 651 22928 696 22956
rect 690 22916 696 22928
rect 748 22916 754 22968
rect 3744 22965 3772 22996
rect 4189 22993 4201 22996
rect 4235 22993 4247 23027
rect 6302 23024 6308 23036
rect 6263 22996 6308 23024
rect 4189 22987 4247 22993
rect 6302 22984 6308 22996
rect 6360 22984 6366 23036
rect 7056 23033 7084 23064
rect 11273 23061 11285 23064
rect 11319 23092 11331 23095
rect 11454 23092 11460 23104
rect 11319 23064 11460 23092
rect 11319 23061 11331 23064
rect 11273 23055 11331 23061
rect 11454 23052 11460 23064
rect 11512 23052 11518 23104
rect 7041 23027 7099 23033
rect 7041 22993 7053 23027
rect 7087 22993 7099 23027
rect 11086 23024 11092 23036
rect 11047 22996 11092 23024
rect 7041 22987 7099 22993
rect 11086 22984 11092 22996
rect 11144 22984 11150 23036
rect 11914 23024 11920 23036
rect 11827 22996 11920 23024
rect 11914 22984 11920 22996
rect 11972 23024 11978 23036
rect 13113 23027 13171 23033
rect 13113 23024 13125 23027
rect 11972 22996 13125 23024
rect 11972 22984 11978 22996
rect 13113 22993 13125 22996
rect 13159 22993 13171 23027
rect 13113 22987 13171 22993
rect 3729 22959 3787 22965
rect 3729 22925 3741 22959
rect 3775 22925 3787 22959
rect 3729 22919 3787 22925
rect 5569 22959 5627 22965
rect 5569 22925 5581 22959
rect 5615 22956 5627 22959
rect 6486 22956 6492 22968
rect 5615 22928 6492 22956
rect 5615 22925 5627 22928
rect 5569 22919 5627 22925
rect 6486 22916 6492 22928
rect 6544 22916 6550 22968
rect 7314 22956 7320 22968
rect 7227 22928 7320 22956
rect 7314 22916 7320 22928
rect 7372 22956 7378 22968
rect 7372 22928 7728 22956
rect 7372 22916 7378 22928
rect 1426 22848 1432 22900
rect 1484 22848 1490 22900
rect 2898 22848 2904 22900
rect 2956 22888 2962 22900
rect 3545 22891 3603 22897
rect 3545 22888 3557 22891
rect 2956 22860 3557 22888
rect 2956 22848 2962 22860
rect 3545 22857 3557 22860
rect 3591 22888 3603 22891
rect 4370 22888 4376 22900
rect 3591 22860 4376 22888
rect 3591 22857 3603 22860
rect 3545 22851 3603 22857
rect 4370 22848 4376 22860
rect 4428 22848 4434 22900
rect 3269 22823 3327 22829
rect 3269 22789 3281 22823
rect 3315 22820 3327 22823
rect 4002 22820 4008 22832
rect 3315 22792 4008 22820
rect 3315 22789 3327 22792
rect 3269 22783 3327 22789
rect 4002 22780 4008 22792
rect 4060 22780 4066 22832
rect 7700 22820 7728 22928
rect 8142 22916 8148 22968
rect 8200 22956 8206 22968
rect 12009 22959 12067 22965
rect 12009 22956 12021 22959
rect 8200 22928 12021 22956
rect 8200 22916 8206 22928
rect 12009 22925 12021 22928
rect 12055 22956 12067 22959
rect 12650 22956 12656 22968
rect 12055 22928 12656 22956
rect 12055 22925 12067 22928
rect 12009 22919 12067 22925
rect 12650 22916 12656 22928
rect 12708 22916 12714 22968
rect 12834 22956 12840 22968
rect 12795 22928 12840 22956
rect 12834 22916 12840 22928
rect 12892 22916 12898 22968
rect 13202 22956 13208 22968
rect 13163 22928 13208 22956
rect 13202 22916 13208 22928
rect 13260 22916 13266 22968
rect 14186 22956 14214 23132
rect 14950 23120 14956 23132
rect 15008 23120 15014 23172
rect 17986 23160 17992 23172
rect 17947 23132 17992 23160
rect 17986 23120 17992 23132
rect 18044 23120 18050 23172
rect 18541 23163 18599 23169
rect 18541 23129 18553 23163
rect 18587 23160 18599 23163
rect 18722 23160 18728 23172
rect 18587 23132 18728 23160
rect 18587 23129 18599 23132
rect 18541 23123 18599 23129
rect 18722 23120 18728 23132
rect 18780 23120 18786 23172
rect 21301 23163 21359 23169
rect 21301 23129 21313 23163
rect 21347 23160 21359 23163
rect 21666 23160 21672 23172
rect 21347 23132 21672 23160
rect 21347 23129 21359 23132
rect 21301 23123 21359 23129
rect 21666 23120 21672 23132
rect 21724 23160 21730 23172
rect 23601 23163 23659 23169
rect 23601 23160 23613 23163
rect 21724 23132 23613 23160
rect 21724 23120 21730 23132
rect 23601 23129 23613 23132
rect 23647 23160 23659 23163
rect 24242 23160 24248 23172
rect 23647 23132 23874 23160
rect 24203 23132 24248 23160
rect 23647 23129 23659 23132
rect 23601 23123 23659 23129
rect 23846 23092 23874 23132
rect 24242 23120 24248 23132
rect 24300 23120 24306 23172
rect 24518 23120 24524 23172
rect 24576 23160 24582 23172
rect 25809 23163 25867 23169
rect 25809 23160 25821 23163
rect 24576 23132 25821 23160
rect 24576 23120 24582 23132
rect 25809 23129 25821 23132
rect 25855 23129 25867 23163
rect 26910 23160 26916 23172
rect 26871 23132 26916 23160
rect 25809 23123 25867 23129
rect 24150 23092 24156 23104
rect 23846 23064 24156 23092
rect 24150 23052 24156 23064
rect 24208 23092 24214 23104
rect 24208 23064 24932 23092
rect 24208 23052 24214 23064
rect 18630 23024 18636 23036
rect 18591 22996 18636 23024
rect 18630 22984 18636 22996
rect 18688 22984 18694 23036
rect 21485 23027 21543 23033
rect 21485 22993 21497 23027
rect 21531 23024 21543 23027
rect 21853 23027 21911 23033
rect 21853 23024 21865 23027
rect 21531 22996 21865 23024
rect 21531 22993 21543 22996
rect 21485 22987 21543 22993
rect 21853 22993 21865 22996
rect 21899 23024 21911 23027
rect 22954 23024 22960 23036
rect 21899 22996 22960 23024
rect 21899 22993 21911 22996
rect 21853 22987 21911 22993
rect 22954 22984 22960 22996
rect 23012 23024 23018 23036
rect 23233 23027 23291 23033
rect 23233 23024 23245 23027
rect 23012 22996 23245 23024
rect 23012 22984 23018 22996
rect 23233 22993 23245 22996
rect 23279 23024 23291 23027
rect 23877 23027 23935 23033
rect 23877 23024 23889 23027
rect 23279 22996 23889 23024
rect 23279 22993 23291 22996
rect 23233 22987 23291 22993
rect 23877 22993 23889 22996
rect 23923 23024 23935 23027
rect 24426 23024 24432 23036
rect 23923 22996 24288 23024
rect 24387 22996 24432 23024
rect 23923 22993 23935 22996
rect 23877 22987 23935 22993
rect 14677 22959 14735 22965
rect 14677 22956 14689 22959
rect 14186 22928 14689 22956
rect 14677 22925 14689 22928
rect 14723 22956 14735 22959
rect 14769 22959 14827 22965
rect 14769 22956 14781 22959
rect 14723 22928 14781 22956
rect 14723 22925 14735 22928
rect 14677 22919 14735 22925
rect 14769 22925 14781 22928
rect 14815 22925 14827 22959
rect 21574 22956 21580 22968
rect 21535 22928 21580 22956
rect 14769 22919 14827 22925
rect 21574 22916 21580 22928
rect 21632 22956 21638 22968
rect 22129 22959 22187 22965
rect 22129 22956 22141 22959
rect 21632 22928 22141 22956
rect 21632 22916 21638 22928
rect 22129 22925 22141 22928
rect 22175 22956 22187 22959
rect 22313 22959 22371 22965
rect 22313 22956 22325 22959
rect 22175 22928 22325 22956
rect 22175 22925 22187 22928
rect 22129 22919 22187 22925
rect 22313 22925 22325 22928
rect 22359 22925 22371 22959
rect 22313 22919 22371 22925
rect 22678 22916 22684 22968
rect 22736 22956 22742 22968
rect 23138 22956 23144 22968
rect 22736 22928 23144 22956
rect 22736 22916 22742 22928
rect 23138 22916 23144 22928
rect 23196 22956 23202 22968
rect 23325 22959 23383 22965
rect 23325 22956 23337 22959
rect 23196 22928 23337 22956
rect 23196 22916 23202 22928
rect 23325 22925 23337 22928
rect 23371 22925 23383 22959
rect 24260 22956 24288 22996
rect 24426 22984 24432 22996
rect 24484 22984 24490 23036
rect 24904 23033 24932 23064
rect 24889 23027 24947 23033
rect 24889 22993 24901 23027
rect 24935 22993 24947 23027
rect 25824 23024 25852 23123
rect 26910 23120 26916 23132
rect 26968 23120 26974 23172
rect 27186 23120 27192 23172
rect 27244 23160 27250 23172
rect 27741 23163 27799 23169
rect 27741 23160 27753 23163
rect 27244 23132 27753 23160
rect 27244 23120 27250 23132
rect 27741 23129 27753 23132
rect 27787 23129 27799 23163
rect 27741 23123 27799 23129
rect 29949 23163 30007 23169
rect 29949 23129 29961 23163
rect 29995 23160 30007 23163
rect 30406 23160 30412 23172
rect 29995 23132 30176 23160
rect 30367 23132 30412 23160
rect 29995 23129 30007 23132
rect 29949 23123 30007 23129
rect 30148 23104 30176 23132
rect 30406 23120 30412 23132
rect 30464 23120 30470 23172
rect 27462 23092 27468 23104
rect 27423 23064 27468 23092
rect 27462 23052 27468 23064
rect 27520 23052 27526 23104
rect 27649 23095 27707 23101
rect 27649 23061 27661 23095
rect 27695 23092 27707 23095
rect 28474 23092 28480 23104
rect 27695 23064 28480 23092
rect 27695 23061 27707 23064
rect 27649 23055 27707 23061
rect 26177 23027 26235 23033
rect 26177 23024 26189 23027
rect 25824 22996 26189 23024
rect 24889 22987 24947 22993
rect 26177 22993 26189 22996
rect 26223 23024 26235 23027
rect 27097 23027 27155 23033
rect 26223 22996 27048 23024
rect 26223 22993 26235 22996
rect 26177 22987 26235 22993
rect 24610 22956 24616 22968
rect 24260 22928 24616 22956
rect 23325 22919 23383 22925
rect 24610 22916 24616 22928
rect 24668 22916 24674 22968
rect 24794 22916 24800 22968
rect 24852 22956 24858 22968
rect 24981 22959 25039 22965
rect 24981 22956 24993 22959
rect 24852 22928 24993 22956
rect 24852 22916 24858 22928
rect 24981 22925 24993 22928
rect 25027 22925 25039 22959
rect 25990 22956 25996 22968
rect 25903 22928 25996 22956
rect 24981 22919 25039 22925
rect 25990 22916 25996 22928
rect 26048 22956 26054 22968
rect 26545 22959 26603 22965
rect 26545 22956 26557 22959
rect 26048 22928 26557 22956
rect 26048 22916 26054 22928
rect 26545 22925 26557 22928
rect 26591 22925 26603 22959
rect 26545 22919 26603 22925
rect 27020 22956 27048 22996
rect 27097 22993 27109 23027
rect 27143 23024 27155 23027
rect 27554 23024 27560 23036
rect 27143 22996 27560 23024
rect 27143 22993 27155 22996
rect 27097 22987 27155 22993
rect 27554 22984 27560 22996
rect 27612 22984 27618 23036
rect 27186 22956 27192 22968
rect 27020 22928 27192 22956
rect 9062 22848 9068 22900
rect 9120 22888 9126 22900
rect 9157 22891 9215 22897
rect 9157 22888 9169 22891
rect 9120 22860 9169 22888
rect 9120 22848 9126 22860
rect 9157 22857 9169 22860
rect 9203 22888 9215 22891
rect 12852 22888 12880 22916
rect 9203 22860 12880 22888
rect 14309 22891 14367 22897
rect 9203 22857 9215 22860
rect 9157 22851 9215 22857
rect 14309 22857 14321 22891
rect 14355 22888 14367 22891
rect 14950 22888 14956 22900
rect 14355 22860 14956 22888
rect 14355 22857 14367 22860
rect 14309 22851 14367 22857
rect 14950 22848 14956 22860
rect 15008 22848 15014 22900
rect 18078 22848 18084 22900
rect 18136 22888 18142 22900
rect 18173 22891 18231 22897
rect 18173 22888 18185 22891
rect 18136 22860 18185 22888
rect 18136 22848 18142 22860
rect 18173 22857 18185 22860
rect 18219 22888 18231 22891
rect 18909 22891 18967 22897
rect 18909 22888 18921 22891
rect 18219 22860 18921 22888
rect 18219 22857 18231 22860
rect 18173 22851 18231 22857
rect 18909 22857 18921 22860
rect 18955 22857 18967 22891
rect 18909 22851 18967 22857
rect 19366 22848 19372 22900
rect 19424 22848 19430 22900
rect 20654 22888 20660 22900
rect 20615 22860 20660 22888
rect 20654 22848 20660 22860
rect 20712 22848 20718 22900
rect 23966 22848 23972 22900
rect 24024 22888 24030 22900
rect 26008 22888 26036 22916
rect 24024 22860 26036 22888
rect 27020 22888 27048 22928
rect 27186 22916 27192 22928
rect 27244 22916 27250 22968
rect 27278 22916 27284 22968
rect 27336 22956 27342 22968
rect 27664 22956 27692 23055
rect 28474 23052 28480 23064
rect 28532 23052 28538 23104
rect 29673 23095 29731 23101
rect 29673 23061 29685 23095
rect 29719 23092 29731 23095
rect 30038 23092 30044 23104
rect 29719 23064 30044 23092
rect 29719 23061 29731 23064
rect 29673 23055 29731 23061
rect 30038 23052 30044 23064
rect 30096 23052 30102 23104
rect 30130 23052 30136 23104
rect 30188 23092 30194 23104
rect 30188 23064 30233 23092
rect 30188 23052 30194 23064
rect 27336 22928 27692 22956
rect 27336 22916 27342 22928
rect 27922 22888 27928 22900
rect 27020 22860 27928 22888
rect 24024 22848 24030 22860
rect 27922 22848 27928 22860
rect 27980 22848 27986 22900
rect 9341 22823 9399 22829
rect 9341 22820 9353 22823
rect 7700 22792 9353 22820
rect 9341 22789 9353 22792
rect 9387 22820 9399 22823
rect 9522 22820 9528 22832
rect 9387 22792 9528 22820
rect 9387 22789 9399 22792
rect 9341 22783 9399 22789
rect 9522 22780 9528 22792
rect 9580 22780 9586 22832
rect 10813 22823 10871 22829
rect 10813 22789 10825 22823
rect 10859 22820 10871 22823
rect 10902 22820 10908 22832
rect 10859 22792 10908 22820
rect 10859 22789 10871 22792
rect 10813 22783 10871 22789
rect 10902 22780 10908 22792
rect 10960 22780 10966 22832
rect 10997 22823 11055 22829
rect 10997 22789 11009 22823
rect 11043 22820 11055 22823
rect 11178 22820 11184 22832
rect 11043 22792 11184 22820
rect 11043 22789 11055 22792
rect 10997 22783 11055 22789
rect 11178 22780 11184 22792
rect 11236 22780 11242 22832
rect 11914 22780 11920 22832
rect 11972 22820 11978 22832
rect 13018 22820 13024 22832
rect 11972 22792 13024 22820
rect 11972 22780 11978 22792
rect 13018 22780 13024 22792
rect 13076 22780 13082 22832
rect 18262 22820 18268 22832
rect 18223 22792 18268 22820
rect 18262 22780 18268 22792
rect 18320 22780 18326 22832
rect 22862 22780 22868 22832
rect 22920 22820 22926 22832
rect 22957 22823 23015 22829
rect 22957 22820 22969 22823
rect 22920 22792 22969 22820
rect 22920 22780 22926 22792
rect 22957 22789 22969 22792
rect 23003 22789 23015 22823
rect 22957 22783 23015 22789
rect 27002 22780 27008 22832
rect 27060 22820 27066 22832
rect 27189 22823 27247 22829
rect 27189 22820 27201 22823
rect 27060 22792 27201 22820
rect 27060 22780 27066 22792
rect 27189 22789 27201 22792
rect 27235 22789 27247 22823
rect 30222 22820 30228 22832
rect 30183 22792 30228 22820
rect 27189 22783 27247 22789
rect 30222 22780 30228 22792
rect 30280 22780 30286 22832
rect 400 22730 31680 22752
rect 400 22678 18870 22730
rect 18922 22678 18934 22730
rect 18986 22678 18998 22730
rect 19050 22678 19062 22730
rect 19114 22678 19126 22730
rect 19178 22678 31680 22730
rect 400 22656 31680 22678
rect 785 22619 843 22625
rect 785 22585 797 22619
rect 831 22616 843 22619
rect 966 22616 972 22628
rect 831 22588 972 22616
rect 831 22585 843 22588
rect 785 22579 843 22585
rect 966 22576 972 22588
rect 1024 22576 1030 22628
rect 1245 22619 1303 22625
rect 1245 22585 1257 22619
rect 1291 22616 1303 22619
rect 1426 22616 1432 22628
rect 1291 22588 1432 22616
rect 1291 22585 1303 22588
rect 1245 22579 1303 22585
rect 1426 22576 1432 22588
rect 1484 22576 1490 22628
rect 2622 22576 2628 22628
rect 2680 22616 2686 22628
rect 6121 22619 6179 22625
rect 6121 22616 6133 22619
rect 2680 22588 6133 22616
rect 2680 22576 2686 22588
rect 6121 22585 6133 22588
rect 6167 22616 6179 22619
rect 6302 22616 6308 22628
rect 6167 22588 6308 22616
rect 6167 22585 6179 22588
rect 6121 22579 6179 22585
rect 6302 22576 6308 22588
rect 6360 22576 6366 22628
rect 6486 22616 6492 22628
rect 6447 22588 6492 22616
rect 6486 22576 6492 22588
rect 6544 22576 6550 22628
rect 12285 22619 12343 22625
rect 12285 22585 12297 22619
rect 12331 22616 12343 22619
rect 13202 22616 13208 22628
rect 12331 22588 13208 22616
rect 12331 22585 12343 22588
rect 12285 22579 12343 22585
rect 13202 22576 13208 22588
rect 13260 22616 13266 22628
rect 15686 22616 15692 22628
rect 13260 22588 15692 22616
rect 13260 22576 13266 22588
rect 15686 22576 15692 22588
rect 15744 22576 15750 22628
rect 18630 22576 18636 22628
rect 18688 22616 18694 22628
rect 18817 22619 18875 22625
rect 18817 22616 18829 22619
rect 18688 22588 18829 22616
rect 18688 22576 18694 22588
rect 18817 22585 18829 22588
rect 18863 22585 18875 22619
rect 18817 22579 18875 22585
rect 19093 22619 19151 22625
rect 19093 22585 19105 22619
rect 19139 22616 19151 22619
rect 19366 22616 19372 22628
rect 19139 22588 19372 22616
rect 19139 22585 19151 22588
rect 19093 22579 19151 22585
rect 19366 22576 19372 22588
rect 19424 22576 19430 22628
rect 23966 22616 23972 22628
rect 22972 22588 23972 22616
rect 6946 22508 6952 22560
rect 7004 22548 7010 22560
rect 7004 22520 10028 22548
rect 7004 22508 7010 22520
rect 10000 22492 10028 22520
rect 10718 22508 10724 22560
rect 10776 22508 10782 22560
rect 21850 22508 21856 22560
rect 21908 22548 21914 22560
rect 22037 22551 22095 22557
rect 22037 22548 22049 22551
rect 21908 22520 22049 22548
rect 21908 22508 21914 22520
rect 22037 22517 22049 22520
rect 22083 22517 22095 22551
rect 22037 22511 22095 22517
rect 22972 22492 23000 22588
rect 23966 22576 23972 22588
rect 24024 22576 24030 22628
rect 24061 22619 24119 22625
rect 24061 22585 24073 22619
rect 24107 22616 24119 22619
rect 24426 22616 24432 22628
rect 24107 22588 24432 22616
rect 24107 22585 24119 22588
rect 24061 22579 24119 22585
rect 24426 22576 24432 22588
rect 24484 22576 24490 22628
rect 23230 22548 23236 22560
rect 23156 22520 23236 22548
rect 3266 22440 3272 22492
rect 3324 22480 3330 22492
rect 3913 22483 3971 22489
rect 3913 22480 3925 22483
rect 3324 22452 3925 22480
rect 3324 22440 3330 22452
rect 3913 22449 3925 22452
rect 3959 22449 3971 22483
rect 4094 22480 4100 22492
rect 4055 22452 4100 22480
rect 3913 22443 3971 22449
rect 4094 22440 4100 22452
rect 4152 22440 4158 22492
rect 4554 22440 4560 22492
rect 4612 22480 4618 22492
rect 4612 22452 4657 22480
rect 4612 22440 4618 22452
rect 4922 22440 4928 22492
rect 4980 22480 4986 22492
rect 5017 22483 5075 22489
rect 5017 22480 5029 22483
rect 4980 22452 5029 22480
rect 4980 22440 4986 22452
rect 5017 22449 5029 22452
rect 5063 22449 5075 22483
rect 5017 22443 5075 22449
rect 6118 22440 6124 22492
rect 6176 22480 6182 22492
rect 7409 22483 7467 22489
rect 7409 22480 7421 22483
rect 6176 22452 7421 22480
rect 6176 22440 6182 22452
rect 7409 22449 7421 22452
rect 7455 22480 7467 22483
rect 8142 22480 8148 22492
rect 7455 22452 8148 22480
rect 7455 22449 7467 22452
rect 7409 22443 7467 22449
rect 8142 22440 8148 22452
rect 8200 22440 8206 22492
rect 9982 22480 9988 22492
rect 9895 22452 9988 22480
rect 9982 22440 9988 22452
rect 10040 22440 10046 22492
rect 13018 22480 13024 22492
rect 12979 22452 13024 22480
rect 13018 22440 13024 22452
rect 13076 22440 13082 22492
rect 14677 22483 14735 22489
rect 14677 22449 14689 22483
rect 14723 22480 14735 22483
rect 15134 22480 15140 22492
rect 14723 22452 15140 22480
rect 14723 22449 14735 22452
rect 14677 22443 14735 22449
rect 15134 22440 15140 22452
rect 15192 22480 15198 22492
rect 15962 22480 15968 22492
rect 15192 22452 15968 22480
rect 15192 22440 15198 22452
rect 15962 22440 15968 22452
rect 16020 22440 16026 22492
rect 16330 22480 16336 22492
rect 16291 22452 16336 22480
rect 16330 22440 16336 22452
rect 16388 22440 16394 22492
rect 21758 22440 21764 22492
rect 21816 22480 21822 22492
rect 22497 22483 22555 22489
rect 22497 22480 22509 22483
rect 21816 22452 22509 22480
rect 21816 22440 21822 22452
rect 22497 22449 22509 22452
rect 22543 22449 22555 22483
rect 22678 22480 22684 22492
rect 22639 22452 22684 22480
rect 22497 22443 22555 22449
rect 22678 22440 22684 22452
rect 22736 22440 22742 22492
rect 22954 22480 22960 22492
rect 22915 22452 22960 22480
rect 22954 22440 22960 22452
rect 23012 22440 23018 22492
rect 23156 22489 23184 22520
rect 23230 22508 23236 22520
rect 23288 22508 23294 22560
rect 27094 22508 27100 22560
rect 27152 22548 27158 22560
rect 27152 22520 28704 22548
rect 27152 22508 27158 22520
rect 23141 22483 23199 22489
rect 23141 22449 23153 22483
rect 23187 22449 23199 22483
rect 23141 22443 23199 22449
rect 26174 22440 26180 22492
rect 26232 22480 26238 22492
rect 26361 22483 26419 22489
rect 26361 22480 26373 22483
rect 26232 22452 26373 22480
rect 26232 22440 26238 22452
rect 26361 22449 26373 22452
rect 26407 22449 26419 22483
rect 26361 22443 26419 22449
rect 26545 22483 26603 22489
rect 26545 22449 26557 22483
rect 26591 22449 26603 22483
rect 26545 22443 26603 22449
rect 4112 22412 4140 22440
rect 5934 22412 5940 22424
rect 4112 22384 5940 22412
rect 5934 22372 5940 22384
rect 5992 22372 5998 22424
rect 7590 22412 7596 22424
rect 7551 22384 7596 22412
rect 7590 22372 7596 22384
rect 7648 22372 7654 22424
rect 10353 22415 10411 22421
rect 10353 22381 10365 22415
rect 10399 22412 10411 22415
rect 10718 22412 10724 22424
rect 10399 22384 10724 22412
rect 10399 22381 10411 22384
rect 10353 22375 10411 22381
rect 10718 22372 10724 22384
rect 10776 22372 10782 22424
rect 10902 22372 10908 22424
rect 10960 22412 10966 22424
rect 11546 22412 11552 22424
rect 10960 22384 11552 22412
rect 10960 22372 10966 22384
rect 11546 22372 11552 22384
rect 11604 22412 11610 22424
rect 11733 22415 11791 22421
rect 11733 22412 11745 22415
rect 11604 22384 11745 22412
rect 11604 22372 11610 22384
rect 11733 22381 11745 22384
rect 11779 22381 11791 22415
rect 11733 22375 11791 22381
rect 13481 22415 13539 22421
rect 13481 22381 13493 22415
rect 13527 22412 13539 22415
rect 14766 22412 14772 22424
rect 13527 22384 14772 22412
rect 13527 22381 13539 22384
rect 13481 22375 13539 22381
rect 14766 22372 14772 22384
rect 14824 22412 14830 22424
rect 14861 22415 14919 22421
rect 14861 22412 14873 22415
rect 14824 22384 14873 22412
rect 14824 22372 14830 22384
rect 14861 22381 14873 22384
rect 14907 22381 14919 22415
rect 14861 22375 14919 22381
rect 23230 22372 23236 22424
rect 23288 22412 23294 22424
rect 23417 22415 23475 22421
rect 23417 22412 23429 22415
rect 23288 22384 23429 22412
rect 23288 22372 23294 22384
rect 23417 22381 23429 22384
rect 23463 22381 23475 22415
rect 23417 22375 23475 22381
rect 25990 22372 25996 22424
rect 26048 22412 26054 22424
rect 26560 22412 26588 22443
rect 26910 22440 26916 22492
rect 26968 22480 26974 22492
rect 27005 22483 27063 22489
rect 27005 22480 27017 22483
rect 26968 22452 27017 22480
rect 26968 22440 26974 22452
rect 27005 22449 27017 22452
rect 27051 22449 27063 22483
rect 27005 22443 27063 22449
rect 27465 22483 27523 22489
rect 27465 22449 27477 22483
rect 27511 22449 27523 22483
rect 28566 22480 28572 22492
rect 28527 22452 28572 22480
rect 27465 22443 27523 22449
rect 26048 22384 26588 22412
rect 26048 22372 26054 22384
rect 3174 22304 3180 22356
rect 3232 22344 3238 22356
rect 3361 22347 3419 22353
rect 3361 22344 3373 22347
rect 3232 22316 3373 22344
rect 3232 22304 3238 22316
rect 3361 22313 3373 22316
rect 3407 22313 3419 22347
rect 3361 22307 3419 22313
rect 3729 22347 3787 22353
rect 3729 22313 3741 22347
rect 3775 22344 3787 22347
rect 3910 22344 3916 22356
rect 3775 22316 3916 22344
rect 3775 22313 3787 22316
rect 3729 22307 3787 22313
rect 3910 22304 3916 22316
rect 3968 22344 3974 22356
rect 4186 22344 4192 22356
rect 3968 22316 4192 22344
rect 3968 22304 3974 22316
rect 4186 22304 4192 22316
rect 4244 22304 4250 22356
rect 5566 22304 5572 22356
rect 5624 22344 5630 22356
rect 6857 22347 6915 22353
rect 6857 22344 6869 22347
rect 5624 22316 6869 22344
rect 5624 22304 5630 22316
rect 6857 22313 6869 22316
rect 6903 22344 6915 22347
rect 7038 22344 7044 22356
rect 6903 22316 7044 22344
rect 6903 22313 6915 22316
rect 6857 22307 6915 22313
rect 7038 22304 7044 22316
rect 7096 22304 7102 22356
rect 15686 22304 15692 22356
rect 15744 22344 15750 22356
rect 25806 22344 25812 22356
rect 15744 22316 16652 22344
rect 25767 22316 25812 22344
rect 15744 22304 15750 22316
rect 16624 22288 16652 22316
rect 25806 22304 25812 22316
rect 25864 22304 25870 22356
rect 25898 22304 25904 22356
rect 25956 22344 25962 22356
rect 25956 22316 26001 22344
rect 25956 22304 25962 22316
rect 690 22236 696 22288
rect 748 22276 754 22288
rect 877 22279 935 22285
rect 877 22276 889 22279
rect 748 22248 889 22276
rect 748 22236 754 22248
rect 877 22245 889 22248
rect 923 22245 935 22279
rect 1334 22276 1340 22288
rect 1295 22248 1340 22276
rect 877 22239 935 22245
rect 1334 22236 1340 22248
rect 1392 22236 1398 22288
rect 6302 22276 6308 22288
rect 6263 22248 6308 22276
rect 6302 22236 6308 22248
rect 6360 22236 6366 22288
rect 12650 22236 12656 22288
rect 12708 22276 12714 22288
rect 13021 22279 13079 22285
rect 13021 22276 13033 22279
rect 12708 22248 13033 22276
rect 12708 22236 12714 22248
rect 13021 22245 13033 22248
rect 13067 22276 13079 22279
rect 16514 22276 16520 22288
rect 13067 22248 16520 22276
rect 13067 22245 13079 22248
rect 13021 22239 13079 22245
rect 16514 22236 16520 22248
rect 16572 22236 16578 22288
rect 16606 22236 16612 22288
rect 16664 22276 16670 22288
rect 17437 22279 17495 22285
rect 16664 22248 16709 22276
rect 16664 22236 16670 22248
rect 17437 22245 17449 22279
rect 17483 22276 17495 22279
rect 17618 22276 17624 22288
rect 17483 22248 17624 22276
rect 17483 22245 17495 22248
rect 17437 22239 17495 22245
rect 17618 22236 17624 22248
rect 17676 22236 17682 22288
rect 18725 22279 18783 22285
rect 18725 22245 18737 22279
rect 18771 22276 18783 22279
rect 20654 22276 20660 22288
rect 18771 22248 20660 22276
rect 18771 22245 18783 22248
rect 18725 22239 18783 22245
rect 20654 22236 20660 22248
rect 20712 22236 20718 22288
rect 25530 22236 25536 22288
rect 25588 22276 25594 22288
rect 26266 22276 26272 22288
rect 25588 22248 26272 22276
rect 25588 22236 25594 22248
rect 26266 22236 26272 22248
rect 26324 22276 26330 22288
rect 27480 22276 27508 22443
rect 28566 22440 28572 22452
rect 28624 22440 28630 22492
rect 28676 22489 28704 22520
rect 28661 22483 28719 22489
rect 28661 22449 28673 22483
rect 28707 22480 28719 22483
rect 28750 22480 28756 22492
rect 28707 22452 28756 22480
rect 28707 22449 28719 22452
rect 28661 22443 28719 22449
rect 28750 22440 28756 22452
rect 28808 22440 28814 22492
rect 28842 22276 28848 22288
rect 26324 22248 27508 22276
rect 28803 22248 28848 22276
rect 26324 22236 26330 22248
rect 28842 22236 28848 22248
rect 28900 22236 28906 22288
rect 400 22186 31680 22208
rect 400 22134 3510 22186
rect 3562 22134 3574 22186
rect 3626 22134 3638 22186
rect 3690 22134 3702 22186
rect 3754 22134 3766 22186
rect 3818 22134 31680 22186
rect 400 22112 31680 22134
rect 2349 22075 2407 22081
rect 2349 22041 2361 22075
rect 2395 22072 2407 22075
rect 2898 22072 2904 22084
rect 2395 22044 2904 22072
rect 2395 22041 2407 22044
rect 2349 22035 2407 22041
rect 2898 22032 2904 22044
rect 2956 22032 2962 22084
rect 3266 22072 3272 22084
rect 3227 22044 3272 22072
rect 3266 22032 3272 22044
rect 3324 22032 3330 22084
rect 3637 22075 3695 22081
rect 3637 22041 3649 22075
rect 3683 22072 3695 22075
rect 4094 22072 4100 22084
rect 3683 22044 4100 22072
rect 3683 22041 3695 22044
rect 3637 22035 3695 22041
rect 4094 22032 4100 22044
rect 4152 22032 4158 22084
rect 4186 22032 4192 22084
rect 4244 22072 4250 22084
rect 5017 22075 5075 22081
rect 5017 22072 5029 22075
rect 4244 22044 5029 22072
rect 4244 22032 4250 22044
rect 5017 22041 5029 22044
rect 5063 22041 5075 22075
rect 5934 22072 5940 22084
rect 5847 22044 5940 22072
rect 5017 22035 5075 22041
rect 5934 22032 5940 22044
rect 5992 22072 5998 22084
rect 8142 22072 8148 22084
rect 5992 22044 7176 22072
rect 8103 22044 8148 22072
rect 5992 22032 5998 22044
rect 3284 22004 3312 22032
rect 4738 22004 4744 22016
rect 3284 21976 4744 22004
rect 4738 21964 4744 21976
rect 4796 21964 4802 22016
rect 4922 22004 4928 22016
rect 4883 21976 4928 22004
rect 4922 21964 4928 21976
rect 4980 21964 4986 22016
rect 6486 22004 6492 22016
rect 6447 21976 6492 22004
rect 6486 21964 6492 21976
rect 6544 21964 6550 22016
rect 4278 21936 4284 21948
rect 3836 21908 4140 21936
rect 4239 21908 4284 21936
rect 3836 21877 3864 21908
rect 4112 21880 4140 21908
rect 4278 21896 4284 21908
rect 4336 21936 4342 21948
rect 4940 21936 4968 21964
rect 4336 21908 4968 21936
rect 5385 21939 5443 21945
rect 4336 21896 4342 21908
rect 5385 21905 5397 21939
rect 5431 21936 5443 21939
rect 7148 21936 7176 22044
rect 8142 22032 8148 22044
rect 8200 22032 8206 22084
rect 10445 22075 10503 22081
rect 10445 22041 10457 22075
rect 10491 22072 10503 22075
rect 10810 22072 10816 22084
rect 10491 22044 10816 22072
rect 10491 22041 10503 22044
rect 10445 22035 10503 22041
rect 10810 22032 10816 22044
rect 10868 22032 10874 22084
rect 16514 22032 16520 22084
rect 16572 22072 16578 22084
rect 16885 22075 16943 22081
rect 16885 22072 16897 22075
rect 16572 22044 16897 22072
rect 16572 22032 16578 22044
rect 16885 22041 16897 22044
rect 16931 22041 16943 22075
rect 21758 22072 21764 22084
rect 21719 22044 21764 22072
rect 16885 22035 16943 22041
rect 10077 22007 10135 22013
rect 10077 21973 10089 22007
rect 10123 22004 10135 22007
rect 10902 22004 10908 22016
rect 10123 21976 10908 22004
rect 10123 21973 10135 21976
rect 10077 21967 10135 21973
rect 10902 21964 10908 21976
rect 10960 21964 10966 22016
rect 11454 21964 11460 22016
rect 11512 22004 11518 22016
rect 13205 22007 13263 22013
rect 13205 22004 13217 22007
rect 11512 21976 13217 22004
rect 11512 21964 11518 21976
rect 13205 21973 13217 21976
rect 13251 22004 13263 22007
rect 16606 22004 16612 22016
rect 13251 21976 13524 22004
rect 16567 21976 16612 22004
rect 13251 21973 13263 21976
rect 13205 21967 13263 21973
rect 10994 21936 11000 21948
rect 5431 21908 6440 21936
rect 5431 21905 5443 21908
rect 5385 21899 5443 21905
rect 2533 21871 2591 21877
rect 2533 21837 2545 21871
rect 2579 21868 2591 21871
rect 2625 21871 2683 21877
rect 2625 21868 2637 21871
rect 2579 21840 2637 21868
rect 2579 21837 2591 21840
rect 2533 21831 2591 21837
rect 2625 21837 2637 21840
rect 2671 21868 2683 21871
rect 3821 21871 3879 21877
rect 3821 21868 3833 21871
rect 2671 21840 3833 21868
rect 2671 21837 2683 21840
rect 2625 21831 2683 21837
rect 3821 21837 3833 21840
rect 3867 21837 3879 21871
rect 4002 21868 4008 21880
rect 3915 21840 4008 21868
rect 3821 21831 3879 21837
rect 2714 21692 2720 21744
rect 2772 21732 2778 21744
rect 3174 21732 3180 21744
rect 2772 21704 3180 21732
rect 2772 21692 2778 21704
rect 3174 21692 3180 21704
rect 3232 21732 3238 21744
rect 3361 21735 3419 21741
rect 3361 21732 3373 21735
rect 3232 21704 3373 21732
rect 3232 21692 3238 21704
rect 3361 21701 3373 21704
rect 3407 21701 3419 21735
rect 3928 21732 3956 21840
rect 4002 21828 4008 21840
rect 4060 21828 4066 21880
rect 4094 21828 4100 21880
rect 4152 21868 4158 21880
rect 4649 21871 4707 21877
rect 4649 21868 4661 21871
rect 4152 21840 4661 21868
rect 4152 21828 4158 21840
rect 4649 21837 4661 21840
rect 4695 21837 4707 21871
rect 4649 21831 4707 21837
rect 4738 21828 4744 21880
rect 4796 21868 4802 21880
rect 5400 21868 5428 21899
rect 6412 21880 6440 21908
rect 7148 21908 11000 21936
rect 4796 21840 5428 21868
rect 5753 21871 5811 21877
rect 4796 21828 4802 21840
rect 5753 21837 5765 21871
rect 5799 21868 5811 21871
rect 6118 21868 6124 21880
rect 5799 21840 6124 21868
rect 5799 21837 5811 21840
rect 5753 21831 5811 21837
rect 6118 21828 6124 21840
rect 6176 21828 6182 21880
rect 6394 21828 6400 21880
rect 6452 21868 6458 21880
rect 7148 21877 7176 21908
rect 10994 21896 11000 21908
rect 11052 21896 11058 21948
rect 13294 21896 13300 21948
rect 13352 21936 13358 21948
rect 13389 21939 13447 21945
rect 13389 21936 13401 21939
rect 13352 21908 13401 21936
rect 13352 21896 13358 21908
rect 13389 21905 13401 21908
rect 13435 21905 13447 21939
rect 13496 21936 13524 21976
rect 16606 21964 16612 21976
rect 16664 21964 16670 22016
rect 15413 21939 15471 21945
rect 15413 21936 15425 21939
rect 13496 21908 15425 21936
rect 13389 21899 13447 21905
rect 15413 21905 15425 21908
rect 15459 21905 15471 21939
rect 16900 21936 16928 22035
rect 21758 22032 21764 22044
rect 21816 22032 21822 22084
rect 21850 22032 21856 22084
rect 21908 22072 21914 22084
rect 22221 22075 22279 22081
rect 22221 22072 22233 22075
rect 21908 22044 22233 22072
rect 21908 22032 21914 22044
rect 22221 22041 22233 22044
rect 22267 22041 22279 22075
rect 22221 22035 22279 22041
rect 25349 22075 25407 22081
rect 25349 22041 25361 22075
rect 25395 22072 25407 22075
rect 25898 22072 25904 22084
rect 25395 22044 25904 22072
rect 25395 22041 25407 22044
rect 25349 22035 25407 22041
rect 25898 22032 25904 22044
rect 25956 22032 25962 22084
rect 28566 22072 28572 22084
rect 28527 22044 28572 22072
rect 28566 22032 28572 22044
rect 28624 22032 28630 22084
rect 28750 22072 28756 22084
rect 28711 22044 28756 22072
rect 28750 22032 28756 22044
rect 28808 22032 28814 22084
rect 28842 22032 28848 22084
rect 28900 22072 28906 22084
rect 28937 22075 28995 22081
rect 28937 22072 28949 22075
rect 28900 22044 28949 22072
rect 28900 22032 28906 22044
rect 28937 22041 28949 22044
rect 28983 22041 28995 22075
rect 28937 22035 28995 22041
rect 17161 22007 17219 22013
rect 17161 21973 17173 22007
rect 17207 22004 17219 22007
rect 21945 22007 22003 22013
rect 17207 21976 18124 22004
rect 17207 21973 17219 21976
rect 17161 21967 17219 21973
rect 18096 21948 18124 21976
rect 21945 21973 21957 22007
rect 21991 22004 22003 22007
rect 22678 22004 22684 22016
rect 21991 21976 22684 22004
rect 21991 21973 22003 21976
rect 21945 21967 22003 21973
rect 22678 21964 22684 21976
rect 22736 21964 22742 22016
rect 25530 22004 25536 22016
rect 25491 21976 25536 22004
rect 25530 21964 25536 21976
rect 25588 21964 25594 22016
rect 25809 22007 25867 22013
rect 25809 21973 25821 22007
rect 25855 22004 25867 22007
rect 26174 22004 26180 22016
rect 25855 21976 26180 22004
rect 25855 21973 25867 21976
rect 25809 21967 25867 21973
rect 26174 21964 26180 21976
rect 26232 21964 26238 22016
rect 26358 21964 26364 22016
rect 26416 22004 26422 22016
rect 27281 22007 27339 22013
rect 27281 22004 27293 22007
rect 26416 21976 27293 22004
rect 26416 21964 26422 21976
rect 27281 21973 27293 21976
rect 27327 22004 27339 22007
rect 28658 22004 28664 22016
rect 27327 21976 28664 22004
rect 27327 21973 27339 21976
rect 27281 21967 27339 21973
rect 28658 21964 28664 21976
rect 28716 22004 28722 22016
rect 30222 22004 30228 22016
rect 28716 21976 30228 22004
rect 28716 21964 28722 21976
rect 30222 21964 30228 21976
rect 30280 21964 30286 22016
rect 18078 21936 18084 21948
rect 16900 21908 17572 21936
rect 18039 21908 18084 21936
rect 15413 21899 15471 21905
rect 6673 21871 6731 21877
rect 6673 21868 6685 21871
rect 6452 21840 6685 21868
rect 6452 21828 6458 21840
rect 6673 21837 6685 21840
rect 6719 21837 6731 21871
rect 6673 21831 6731 21837
rect 7133 21871 7191 21877
rect 7133 21837 7145 21871
rect 7179 21837 7191 21871
rect 7133 21831 7191 21837
rect 7409 21871 7467 21877
rect 7409 21837 7421 21871
rect 7455 21837 7467 21871
rect 7774 21868 7780 21880
rect 7735 21840 7780 21868
rect 7409 21831 7467 21837
rect 4557 21735 4615 21741
rect 4557 21732 4569 21735
rect 3928 21704 4569 21732
rect 3361 21695 3419 21701
rect 4557 21701 4569 21704
rect 4603 21732 4615 21735
rect 4830 21732 4836 21744
rect 4603 21704 4836 21732
rect 4603 21701 4615 21704
rect 4557 21695 4615 21701
rect 4830 21692 4836 21704
rect 4888 21692 4894 21744
rect 5569 21735 5627 21741
rect 5569 21701 5581 21735
rect 5615 21732 5627 21735
rect 7424 21732 7452 21831
rect 7774 21828 7780 21840
rect 7832 21828 7838 21880
rect 9982 21828 9988 21880
rect 10040 21868 10046 21880
rect 10537 21871 10595 21877
rect 10537 21868 10549 21871
rect 10040 21840 10549 21868
rect 10040 21828 10046 21840
rect 10537 21837 10549 21840
rect 10583 21868 10595 21871
rect 12190 21868 12196 21880
rect 10583 21840 12196 21868
rect 10583 21837 10595 21840
rect 10537 21831 10595 21837
rect 12190 21828 12196 21840
rect 12248 21828 12254 21880
rect 14766 21828 14772 21880
rect 14824 21828 14830 21880
rect 15428 21868 15456 21899
rect 17544 21877 17572 21908
rect 18078 21896 18084 21908
rect 18136 21896 18142 21948
rect 22129 21939 22187 21945
rect 22129 21905 22141 21939
rect 22175 21936 22187 21939
rect 22770 21936 22776 21948
rect 22175 21908 22776 21936
rect 22175 21905 22187 21908
rect 22129 21899 22187 21905
rect 22770 21896 22776 21908
rect 22828 21936 22834 21948
rect 23138 21936 23144 21948
rect 22828 21908 23144 21936
rect 22828 21896 22834 21908
rect 23138 21896 23144 21908
rect 23196 21896 23202 21948
rect 25717 21939 25775 21945
rect 25717 21905 25729 21939
rect 25763 21936 25775 21939
rect 26269 21939 26327 21945
rect 26269 21936 26281 21939
rect 25763 21908 26281 21936
rect 25763 21905 25775 21908
rect 25717 21899 25775 21905
rect 26269 21905 26281 21908
rect 26315 21936 26327 21939
rect 26910 21936 26916 21948
rect 26315 21908 26916 21936
rect 26315 21905 26327 21908
rect 26269 21899 26327 21905
rect 26910 21896 26916 21908
rect 26968 21896 26974 21948
rect 17345 21871 17403 21877
rect 17345 21868 17357 21871
rect 15428 21840 17357 21868
rect 17345 21837 17357 21840
rect 17391 21837 17403 21871
rect 17345 21831 17403 21837
rect 17529 21871 17587 21877
rect 17529 21837 17541 21871
rect 17575 21837 17587 21871
rect 17529 21831 17587 21837
rect 10261 21803 10319 21809
rect 10261 21769 10273 21803
rect 10307 21800 10319 21803
rect 10718 21800 10724 21812
rect 10307 21772 10724 21800
rect 10307 21769 10319 21772
rect 10261 21763 10319 21769
rect 10718 21760 10724 21772
rect 10776 21760 10782 21812
rect 12006 21760 12012 21812
rect 12064 21800 12070 21812
rect 13113 21803 13171 21809
rect 13113 21800 13125 21803
rect 12064 21772 13125 21800
rect 12064 21760 12070 21772
rect 13113 21769 13125 21772
rect 13159 21800 13171 21803
rect 13665 21803 13723 21809
rect 13665 21800 13677 21803
rect 13159 21772 13677 21800
rect 13159 21769 13171 21772
rect 13113 21763 13171 21769
rect 13665 21769 13677 21772
rect 13711 21769 13723 21803
rect 17360 21800 17388 21831
rect 17618 21828 17624 21880
rect 17676 21868 17682 21880
rect 17676 21840 17721 21868
rect 17676 21828 17682 21840
rect 18354 21828 18360 21880
rect 18412 21868 18418 21880
rect 19093 21871 19151 21877
rect 19093 21868 19105 21871
rect 18412 21840 19105 21868
rect 18412 21828 18418 21840
rect 19093 21837 19105 21840
rect 19139 21868 19151 21871
rect 19553 21871 19611 21877
rect 19553 21868 19565 21871
rect 19139 21840 19565 21868
rect 19139 21837 19151 21840
rect 19093 21831 19151 21837
rect 19553 21837 19565 21840
rect 19599 21837 19611 21871
rect 19553 21831 19611 21837
rect 21482 21828 21488 21880
rect 21540 21868 21546 21880
rect 22405 21871 22463 21877
rect 22405 21868 22417 21871
rect 21540 21840 22417 21868
rect 21540 21828 21546 21840
rect 22405 21837 22417 21840
rect 22451 21868 22463 21871
rect 22954 21868 22960 21880
rect 22451 21840 22960 21868
rect 22451 21837 22463 21840
rect 22405 21831 22463 21837
rect 22954 21828 22960 21840
rect 23012 21828 23018 21880
rect 26358 21868 26364 21880
rect 26319 21840 26364 21868
rect 26358 21828 26364 21840
rect 26416 21828 26422 21880
rect 26450 21828 26456 21880
rect 26508 21868 26514 21880
rect 26545 21871 26603 21877
rect 26545 21868 26557 21871
rect 26508 21840 26557 21868
rect 26508 21828 26514 21840
rect 26545 21837 26557 21840
rect 26591 21868 26603 21871
rect 26591 21840 27140 21868
rect 26591 21837 26603 21840
rect 26545 21831 26603 21837
rect 18173 21803 18231 21809
rect 18173 21800 18185 21803
rect 17360 21772 18185 21800
rect 13665 21763 13723 21769
rect 18173 21769 18185 21772
rect 18219 21800 18231 21803
rect 18262 21800 18268 21812
rect 18219 21772 18268 21800
rect 18219 21769 18231 21772
rect 18173 21763 18231 21769
rect 18262 21760 18268 21772
rect 18320 21760 18326 21812
rect 18909 21803 18967 21809
rect 18909 21769 18921 21803
rect 18955 21800 18967 21803
rect 19829 21803 19887 21809
rect 19829 21800 19841 21803
rect 18955 21772 19841 21800
rect 18955 21769 18967 21772
rect 18909 21763 18967 21769
rect 19829 21769 19841 21772
rect 19875 21800 19887 21803
rect 24518 21800 24524 21812
rect 19875 21772 24524 21800
rect 19875 21769 19887 21772
rect 19829 21763 19887 21769
rect 24518 21760 24524 21772
rect 24576 21760 24582 21812
rect 27112 21744 27140 21840
rect 8694 21732 8700 21744
rect 5615 21704 8700 21732
rect 5615 21701 5627 21704
rect 5569 21695 5627 21701
rect 8694 21692 8700 21704
rect 8752 21692 8758 21744
rect 12650 21732 12656 21744
rect 12611 21704 12656 21732
rect 12650 21692 12656 21704
rect 12708 21692 12714 21744
rect 12929 21735 12987 21741
rect 12929 21701 12941 21735
rect 12975 21732 12987 21735
rect 13018 21732 13024 21744
rect 12975 21704 13024 21732
rect 12975 21701 12987 21704
rect 12929 21695 12987 21701
rect 13018 21692 13024 21704
rect 13076 21692 13082 21744
rect 15134 21692 15140 21744
rect 15192 21732 15198 21744
rect 15505 21735 15563 21741
rect 15505 21732 15517 21735
rect 15192 21704 15517 21732
rect 15192 21692 15198 21704
rect 15505 21701 15517 21704
rect 15551 21701 15563 21735
rect 16330 21732 16336 21744
rect 16291 21704 16336 21732
rect 15505 21695 15563 21701
rect 16330 21692 16336 21704
rect 16388 21692 16394 21744
rect 18722 21732 18728 21744
rect 18683 21704 18728 21732
rect 18722 21692 18728 21704
rect 18780 21732 18786 21744
rect 19185 21735 19243 21741
rect 19185 21732 19197 21735
rect 18780 21704 19197 21732
rect 18780 21692 18786 21704
rect 19185 21701 19197 21704
rect 19231 21701 19243 21735
rect 19185 21695 19243 21701
rect 22681 21735 22739 21741
rect 22681 21701 22693 21735
rect 22727 21732 22739 21735
rect 23230 21732 23236 21744
rect 22727 21704 23236 21732
rect 22727 21701 22739 21704
rect 22681 21695 22739 21701
rect 23230 21692 23236 21704
rect 23288 21692 23294 21744
rect 25990 21732 25996 21744
rect 25951 21704 25996 21732
rect 25990 21692 25996 21704
rect 26048 21692 26054 21744
rect 27094 21732 27100 21744
rect 27055 21704 27100 21732
rect 27094 21692 27100 21704
rect 27152 21692 27158 21744
rect 400 21642 31680 21664
rect 400 21590 18870 21642
rect 18922 21590 18934 21642
rect 18986 21590 18998 21642
rect 19050 21590 19062 21642
rect 19114 21590 19126 21642
rect 19178 21590 31680 21642
rect 400 21568 31680 21590
rect 3453 21531 3511 21537
rect 3453 21497 3465 21531
rect 3499 21528 3511 21531
rect 4554 21528 4560 21540
rect 3499 21500 4560 21528
rect 3499 21497 3511 21500
rect 3453 21491 3511 21497
rect 4554 21488 4560 21500
rect 4612 21488 4618 21540
rect 7222 21488 7228 21540
rect 7280 21528 7286 21540
rect 7501 21531 7559 21537
rect 7501 21528 7513 21531
rect 7280 21500 7513 21528
rect 7280 21488 7286 21500
rect 7501 21497 7513 21500
rect 7547 21528 7559 21531
rect 7590 21528 7596 21540
rect 7547 21500 7596 21528
rect 7547 21497 7559 21500
rect 7501 21491 7559 21497
rect 7590 21488 7596 21500
rect 7648 21488 7654 21540
rect 13294 21488 13300 21540
rect 13352 21528 13358 21540
rect 13389 21531 13447 21537
rect 13389 21528 13401 21531
rect 13352 21500 13401 21528
rect 13352 21488 13358 21500
rect 13389 21497 13401 21500
rect 13435 21497 13447 21531
rect 14766 21528 14772 21540
rect 14727 21500 14772 21528
rect 13389 21491 13447 21497
rect 14766 21488 14772 21500
rect 14824 21488 14830 21540
rect 16977 21531 17035 21537
rect 16977 21497 16989 21531
rect 17023 21528 17035 21531
rect 17342 21528 17348 21540
rect 17023 21500 17348 21528
rect 17023 21497 17035 21500
rect 16977 21491 17035 21497
rect 17342 21488 17348 21500
rect 17400 21488 17406 21540
rect 23414 21528 23420 21540
rect 23375 21500 23420 21528
rect 23414 21488 23420 21500
rect 23472 21488 23478 21540
rect 27554 21488 27560 21540
rect 27612 21528 27618 21540
rect 27612 21500 27784 21528
rect 27612 21488 27618 21500
rect 3637 21463 3695 21469
rect 3637 21429 3649 21463
rect 3683 21460 3695 21463
rect 4278 21460 4284 21472
rect 3683 21432 4284 21460
rect 3683 21429 3695 21432
rect 3637 21423 3695 21429
rect 4278 21420 4284 21432
rect 4336 21420 4342 21472
rect 7038 21460 7044 21472
rect 4756 21432 7044 21460
rect 4756 21404 4784 21432
rect 7038 21420 7044 21432
rect 7096 21420 7102 21472
rect 16422 21420 16428 21472
rect 16480 21460 16486 21472
rect 21761 21463 21819 21469
rect 16480 21432 21620 21460
rect 16480 21420 16486 21432
rect 1153 21395 1211 21401
rect 1153 21361 1165 21395
rect 1199 21392 1211 21395
rect 1334 21392 1340 21404
rect 1199 21364 1340 21392
rect 1199 21361 1211 21364
rect 1153 21355 1211 21361
rect 1334 21352 1340 21364
rect 1392 21352 1398 21404
rect 3910 21352 3916 21404
rect 3968 21392 3974 21404
rect 4370 21392 4376 21404
rect 3968 21364 4376 21392
rect 3968 21352 3974 21364
rect 4370 21352 4376 21364
rect 4428 21352 4434 21404
rect 4738 21392 4744 21404
rect 4651 21364 4744 21392
rect 4738 21352 4744 21364
rect 4796 21352 4802 21404
rect 5842 21352 5848 21404
rect 5900 21392 5906 21404
rect 6581 21395 6639 21401
rect 6581 21392 6593 21395
rect 5900 21364 6593 21392
rect 5900 21352 5906 21364
rect 6581 21361 6593 21364
rect 6627 21392 6639 21395
rect 7590 21392 7596 21404
rect 6627 21364 7596 21392
rect 6627 21361 6639 21364
rect 6581 21355 6639 21361
rect 7590 21352 7596 21364
rect 7648 21352 7654 21404
rect 10902 21352 10908 21404
rect 10960 21392 10966 21404
rect 10997 21395 11055 21401
rect 10997 21392 11009 21395
rect 10960 21364 11009 21392
rect 10960 21352 10966 21364
rect 10997 21361 11009 21364
rect 11043 21361 11055 21395
rect 10997 21355 11055 21361
rect 11086 21352 11092 21404
rect 11144 21392 11150 21404
rect 11181 21395 11239 21401
rect 11181 21392 11193 21395
rect 11144 21364 11193 21392
rect 11144 21352 11150 21364
rect 11181 21361 11193 21364
rect 11227 21361 11239 21395
rect 11454 21392 11460 21404
rect 11415 21364 11460 21392
rect 11181 21355 11239 21361
rect 11454 21352 11460 21364
rect 11512 21352 11518 21404
rect 12834 21392 12840 21404
rect 12747 21364 12840 21392
rect 12834 21352 12840 21364
rect 12892 21392 12898 21404
rect 15318 21392 15324 21404
rect 12892 21364 15324 21392
rect 12892 21352 12898 21364
rect 15318 21352 15324 21364
rect 15376 21352 15382 21404
rect 16514 21352 16520 21404
rect 16572 21392 16578 21404
rect 17728 21401 17756 21432
rect 17529 21395 17587 21401
rect 17529 21392 17541 21395
rect 16572 21364 17541 21392
rect 16572 21352 16578 21364
rect 17529 21361 17541 21364
rect 17575 21361 17587 21395
rect 17529 21355 17587 21361
rect 17713 21395 17771 21401
rect 17713 21361 17725 21395
rect 17759 21361 17771 21395
rect 17713 21355 17771 21361
rect 17897 21395 17955 21401
rect 17897 21361 17909 21395
rect 17943 21361 17955 21395
rect 18354 21392 18360 21404
rect 18267 21364 18360 21392
rect 17897 21355 17955 21361
rect 969 21327 1027 21333
rect 969 21293 981 21327
rect 1015 21324 1027 21327
rect 1426 21324 1432 21336
rect 1015 21296 1432 21324
rect 1015 21293 1027 21296
rect 969 21287 1027 21293
rect 1426 21284 1432 21296
rect 1484 21284 1490 21336
rect 3358 21284 3364 21336
rect 3416 21324 3422 21336
rect 3729 21327 3787 21333
rect 3729 21324 3741 21327
rect 3416 21296 3741 21324
rect 3416 21284 3422 21296
rect 3729 21293 3741 21296
rect 3775 21293 3787 21327
rect 3729 21287 3787 21293
rect 4465 21327 4523 21333
rect 4465 21293 4477 21327
rect 4511 21293 4523 21327
rect 4465 21287 4523 21293
rect 4186 21216 4192 21268
rect 4244 21256 4250 21268
rect 4480 21256 4508 21287
rect 4554 21284 4560 21336
rect 4612 21324 4618 21336
rect 4649 21327 4707 21333
rect 4649 21324 4661 21327
rect 4612 21296 4661 21324
rect 4612 21284 4618 21296
rect 4649 21293 4661 21296
rect 4695 21324 4707 21327
rect 5566 21324 5572 21336
rect 4695 21296 5572 21324
rect 4695 21293 4707 21296
rect 4649 21287 4707 21293
rect 5566 21284 5572 21296
rect 5624 21284 5630 21336
rect 5750 21324 5756 21336
rect 5711 21296 5756 21324
rect 5750 21284 5756 21296
rect 5808 21284 5814 21336
rect 6302 21324 6308 21336
rect 6215 21296 6308 21324
rect 6302 21284 6308 21296
rect 6360 21284 6366 21336
rect 6394 21284 6400 21336
rect 6452 21324 6458 21336
rect 6765 21327 6823 21333
rect 6765 21324 6777 21327
rect 6452 21296 6777 21324
rect 6452 21284 6458 21296
rect 6765 21293 6777 21296
rect 6811 21293 6823 21327
rect 6765 21287 6823 21293
rect 10537 21327 10595 21333
rect 10537 21293 10549 21327
rect 10583 21324 10595 21327
rect 10718 21324 10724 21336
rect 10583 21296 10724 21324
rect 10583 21293 10595 21296
rect 10537 21287 10595 21293
rect 10718 21284 10724 21296
rect 10776 21284 10782 21336
rect 10810 21284 10816 21336
rect 10868 21324 10874 21336
rect 11641 21327 11699 21333
rect 11641 21324 11653 21327
rect 10868 21296 11653 21324
rect 10868 21284 10874 21296
rect 11641 21293 11653 21296
rect 11687 21324 11699 21327
rect 11822 21324 11828 21336
rect 11687 21296 11828 21324
rect 11687 21293 11699 21296
rect 11641 21287 11699 21293
rect 11822 21284 11828 21296
rect 11880 21284 11886 21336
rect 11917 21327 11975 21333
rect 11917 21293 11929 21327
rect 11963 21324 11975 21327
rect 13018 21324 13024 21336
rect 11963 21296 13024 21324
rect 11963 21293 11975 21296
rect 11917 21287 11975 21293
rect 5768 21256 5796 21284
rect 4244 21228 5796 21256
rect 6320 21256 6348 21284
rect 7774 21256 7780 21268
rect 6320 21228 7780 21256
rect 4244 21216 4250 21228
rect 7774 21216 7780 21228
rect 7832 21216 7838 21268
rect 11178 21216 11184 21268
rect 11236 21256 11242 21268
rect 11932 21256 11960 21287
rect 13018 21284 13024 21296
rect 13076 21284 13082 21336
rect 17066 21324 17072 21336
rect 17027 21296 17072 21324
rect 17066 21284 17072 21296
rect 17124 21284 17130 21336
rect 17434 21284 17440 21336
rect 17492 21324 17498 21336
rect 17912 21324 17940 21355
rect 18354 21352 18360 21364
rect 18412 21392 18418 21404
rect 19366 21392 19372 21404
rect 18412 21364 19372 21392
rect 18412 21352 18418 21364
rect 19366 21352 19372 21364
rect 19424 21352 19430 21404
rect 21592 21392 21620 21432
rect 21761 21429 21773 21463
rect 21807 21460 21819 21463
rect 21942 21460 21948 21472
rect 21807 21432 21948 21460
rect 21807 21429 21819 21432
rect 21761 21423 21819 21429
rect 21942 21420 21948 21432
rect 22000 21420 22006 21472
rect 22144 21432 22448 21460
rect 22144 21404 22172 21432
rect 22126 21392 22132 21404
rect 21592 21364 22132 21392
rect 22126 21352 22132 21364
rect 22184 21352 22190 21404
rect 22310 21392 22316 21404
rect 22271 21364 22316 21392
rect 22310 21352 22316 21364
rect 22368 21352 22374 21404
rect 22420 21401 22448 21432
rect 27756 21404 27784 21500
rect 22405 21395 22463 21401
rect 22405 21361 22417 21395
rect 22451 21361 22463 21395
rect 22586 21392 22592 21404
rect 22547 21364 22592 21392
rect 22405 21355 22463 21361
rect 22586 21352 22592 21364
rect 22644 21352 22650 21404
rect 23230 21392 23236 21404
rect 23191 21364 23236 21392
rect 23230 21352 23236 21364
rect 23288 21352 23294 21404
rect 24150 21352 24156 21404
rect 24208 21392 24214 21404
rect 24245 21395 24303 21401
rect 24245 21392 24257 21395
rect 24208 21364 24257 21392
rect 24208 21352 24214 21364
rect 24245 21361 24257 21364
rect 24291 21361 24303 21395
rect 27002 21392 27008 21404
rect 24245 21355 24303 21361
rect 25824 21364 27008 21392
rect 25824 21336 25852 21364
rect 27002 21352 27008 21364
rect 27060 21352 27066 21404
rect 27462 21352 27468 21404
rect 27520 21392 27526 21404
rect 27557 21395 27615 21401
rect 27557 21392 27569 21395
rect 27520 21364 27569 21392
rect 27520 21352 27526 21364
rect 27557 21361 27569 21364
rect 27603 21361 27615 21395
rect 27738 21392 27744 21404
rect 27651 21364 27744 21392
rect 27557 21355 27615 21361
rect 27738 21352 27744 21364
rect 27796 21352 27802 21404
rect 28477 21395 28535 21401
rect 28477 21361 28489 21395
rect 28523 21361 28535 21395
rect 28477 21355 28535 21361
rect 17492 21296 17940 21324
rect 18449 21327 18507 21333
rect 17492 21284 17498 21296
rect 18449 21293 18461 21327
rect 18495 21324 18507 21327
rect 18722 21324 18728 21336
rect 18495 21296 18728 21324
rect 18495 21293 18507 21296
rect 18449 21287 18507 21293
rect 11236 21228 11960 21256
rect 11236 21216 11242 21228
rect 16238 21216 16244 21268
rect 16296 21256 16302 21268
rect 18464 21256 18492 21287
rect 18722 21284 18728 21296
rect 18780 21284 18786 21336
rect 22862 21324 22868 21336
rect 22823 21296 22868 21324
rect 22862 21284 22868 21296
rect 22920 21284 22926 21336
rect 24518 21324 24524 21336
rect 24479 21296 24524 21324
rect 24518 21284 24524 21296
rect 24576 21324 24582 21336
rect 25806 21324 25812 21336
rect 24576 21296 25812 21324
rect 24576 21284 24582 21296
rect 25806 21284 25812 21296
rect 25864 21284 25870 21336
rect 26726 21284 26732 21336
rect 26784 21324 26790 21336
rect 26784 21296 27140 21324
rect 26784 21284 26790 21296
rect 27112 21265 27140 21296
rect 27646 21284 27652 21336
rect 27704 21324 27710 21336
rect 28492 21324 28520 21355
rect 28566 21352 28572 21404
rect 28624 21392 28630 21404
rect 28661 21395 28719 21401
rect 28661 21392 28673 21395
rect 28624 21364 28673 21392
rect 28624 21352 28630 21364
rect 28661 21361 28673 21364
rect 28707 21361 28719 21395
rect 28661 21355 28719 21361
rect 29578 21324 29584 21336
rect 27704 21296 29584 21324
rect 27704 21284 27710 21296
rect 29578 21284 29584 21296
rect 29636 21284 29642 21336
rect 16296 21228 18492 21256
rect 27097 21259 27155 21265
rect 16296 21216 16302 21228
rect 27097 21225 27109 21259
rect 27143 21225 27155 21259
rect 27097 21219 27155 21225
rect 785 21191 843 21197
rect 785 21157 797 21191
rect 831 21188 843 21191
rect 2714 21188 2720 21200
rect 831 21160 2720 21188
rect 831 21157 843 21160
rect 785 21151 843 21157
rect 2714 21148 2720 21160
rect 2772 21148 2778 21200
rect 4002 21148 4008 21200
rect 4060 21188 4066 21200
rect 4554 21188 4560 21200
rect 4060 21160 4560 21188
rect 4060 21148 4066 21160
rect 4554 21148 4560 21160
rect 4612 21148 4618 21200
rect 6946 21188 6952 21200
rect 6907 21160 6952 21188
rect 6946 21148 6952 21160
rect 7004 21148 7010 21200
rect 8789 21191 8847 21197
rect 8789 21157 8801 21191
rect 8835 21188 8847 21191
rect 9062 21188 9068 21200
rect 8835 21160 9068 21188
rect 8835 21157 8847 21160
rect 8789 21151 8847 21157
rect 9062 21148 9068 21160
rect 9120 21148 9126 21200
rect 22770 21148 22776 21200
rect 22828 21188 22834 21200
rect 23782 21188 23788 21200
rect 22828 21160 23788 21188
rect 22828 21148 22834 21160
rect 23782 21148 23788 21160
rect 23840 21148 23846 21200
rect 25162 21148 25168 21200
rect 25220 21188 25226 21200
rect 28290 21188 28296 21200
rect 25220 21160 28296 21188
rect 25220 21148 25226 21160
rect 28290 21148 28296 21160
rect 28348 21148 28354 21200
rect 28566 21148 28572 21200
rect 28624 21188 28630 21200
rect 29029 21191 29087 21197
rect 29029 21188 29041 21191
rect 28624 21160 29041 21188
rect 28624 21148 28630 21160
rect 29029 21157 29041 21160
rect 29075 21157 29087 21191
rect 29029 21151 29087 21157
rect 400 21098 31680 21120
rect 400 21046 3510 21098
rect 3562 21046 3574 21098
rect 3626 21046 3638 21098
rect 3690 21046 3702 21098
rect 3754 21046 3766 21098
rect 3818 21046 31680 21098
rect 400 21024 31680 21046
rect 3358 20984 3364 20996
rect 3319 20956 3364 20984
rect 3358 20944 3364 20956
rect 3416 20944 3422 20996
rect 3637 20987 3695 20993
rect 3637 20953 3649 20987
rect 3683 20984 3695 20987
rect 3910 20984 3916 20996
rect 3683 20956 3916 20984
rect 3683 20953 3695 20956
rect 3637 20947 3695 20953
rect 3910 20944 3916 20956
rect 3968 20944 3974 20996
rect 4005 20987 4063 20993
rect 4005 20953 4017 20987
rect 4051 20984 4063 20987
rect 4370 20984 4376 20996
rect 4051 20956 4376 20984
rect 4051 20953 4063 20956
rect 4005 20947 4063 20953
rect 4370 20944 4376 20956
rect 4428 20944 4434 20996
rect 4741 20987 4799 20993
rect 4741 20953 4753 20987
rect 4787 20953 4799 20987
rect 4741 20947 4799 20953
rect 4756 20916 4784 20947
rect 4922 20944 4928 20996
rect 4980 20984 4986 20996
rect 5201 20987 5259 20993
rect 5201 20984 5213 20987
rect 4980 20956 5213 20984
rect 4980 20944 4986 20956
rect 5201 20953 5213 20956
rect 5247 20984 5259 20987
rect 5842 20984 5848 20996
rect 5247 20956 5848 20984
rect 5247 20953 5259 20956
rect 5201 20947 5259 20953
rect 5842 20944 5848 20956
rect 5900 20944 5906 20996
rect 6581 20987 6639 20993
rect 6581 20953 6593 20987
rect 6627 20984 6639 20987
rect 7866 20984 7872 20996
rect 6627 20956 7872 20984
rect 6627 20953 6639 20956
rect 6581 20947 6639 20953
rect 7866 20944 7872 20956
rect 7924 20944 7930 20996
rect 10718 20984 10724 20996
rect 10679 20956 10724 20984
rect 10718 20944 10724 20956
rect 10776 20944 10782 20996
rect 11086 20984 11092 20996
rect 11047 20956 11092 20984
rect 11086 20944 11092 20956
rect 11144 20944 11150 20996
rect 11362 20944 11368 20996
rect 11420 20984 11426 20996
rect 12834 20984 12840 20996
rect 11420 20956 12840 20984
rect 11420 20944 11426 20956
rect 12834 20944 12840 20956
rect 12892 20944 12898 20996
rect 13018 20984 13024 20996
rect 12979 20956 13024 20984
rect 13018 20944 13024 20956
rect 13076 20944 13082 20996
rect 16238 20984 16244 20996
rect 16199 20956 16244 20984
rect 16238 20944 16244 20956
rect 16296 20944 16302 20996
rect 16422 20984 16428 20996
rect 16383 20956 16428 20984
rect 16422 20944 16428 20956
rect 16480 20944 16486 20996
rect 16793 20987 16851 20993
rect 16793 20953 16805 20987
rect 16839 20984 16851 20987
rect 17066 20984 17072 20996
rect 16839 20956 17072 20984
rect 16839 20953 16851 20956
rect 16793 20947 16851 20953
rect 17066 20944 17072 20956
rect 17124 20944 17130 20996
rect 17158 20944 17164 20996
rect 17216 20984 17222 20996
rect 18354 20984 18360 20996
rect 17216 20956 18360 20984
rect 17216 20944 17222 20956
rect 18354 20944 18360 20956
rect 18412 20944 18418 20996
rect 21942 20984 21948 20996
rect 21903 20956 21948 20984
rect 21942 20944 21948 20956
rect 22000 20944 22006 20996
rect 22126 20984 22132 20996
rect 22087 20956 22132 20984
rect 22126 20944 22132 20956
rect 22184 20984 22190 20996
rect 22497 20987 22555 20993
rect 22497 20984 22509 20987
rect 22184 20956 22509 20984
rect 22184 20944 22190 20956
rect 22497 20953 22509 20956
rect 22543 20984 22555 20987
rect 23233 20987 23291 20993
rect 22543 20956 23184 20984
rect 22543 20953 22555 20956
rect 22497 20947 22555 20953
rect 4388 20888 4784 20916
rect 5385 20919 5443 20925
rect 2714 20848 2720 20860
rect 2675 20820 2720 20848
rect 2714 20808 2720 20820
rect 2772 20808 2778 20860
rect 3821 20851 3879 20857
rect 3821 20817 3833 20851
rect 3867 20848 3879 20851
rect 4002 20848 4008 20860
rect 3867 20820 4008 20848
rect 3867 20817 3879 20820
rect 3821 20811 3879 20817
rect 4002 20808 4008 20820
rect 4060 20808 4066 20860
rect 4186 20848 4192 20860
rect 4147 20820 4192 20848
rect 4186 20808 4192 20820
rect 4244 20808 4250 20860
rect 4388 20848 4416 20888
rect 5385 20885 5397 20919
rect 5431 20916 5443 20919
rect 5661 20919 5719 20925
rect 5661 20916 5673 20919
rect 5431 20888 5673 20916
rect 5431 20885 5443 20888
rect 5385 20879 5443 20885
rect 5661 20885 5673 20888
rect 5707 20916 5719 20919
rect 6302 20916 6308 20928
rect 5707 20888 6308 20916
rect 5707 20885 5719 20888
rect 5661 20879 5719 20885
rect 4296 20820 4416 20848
rect 690 20780 696 20792
rect 651 20752 696 20780
rect 690 20740 696 20752
rect 748 20740 754 20792
rect 4094 20740 4100 20792
rect 4152 20780 4158 20792
rect 4296 20789 4324 20820
rect 4462 20808 4468 20860
rect 4520 20848 4526 20860
rect 4738 20848 4744 20860
rect 4520 20820 4744 20848
rect 4520 20808 4526 20820
rect 4738 20808 4744 20820
rect 4796 20808 4802 20860
rect 4281 20783 4339 20789
rect 4281 20780 4293 20783
rect 4152 20752 4293 20780
rect 4152 20740 4158 20752
rect 4281 20749 4293 20752
rect 4327 20749 4339 20783
rect 4281 20743 4339 20749
rect 4649 20783 4707 20789
rect 4649 20749 4661 20783
rect 4695 20780 4707 20783
rect 4922 20780 4928 20792
rect 4695 20752 4928 20780
rect 4695 20749 4707 20752
rect 4649 20743 4707 20749
rect 4922 20740 4928 20752
rect 4980 20740 4986 20792
rect 969 20715 1027 20721
rect 969 20681 981 20715
rect 1015 20681 1027 20715
rect 969 20675 1027 20681
rect 782 20604 788 20656
rect 840 20644 846 20656
rect 984 20644 1012 20675
rect 1426 20672 1432 20724
rect 1484 20672 1490 20724
rect 4465 20715 4523 20721
rect 4465 20681 4477 20715
rect 4511 20712 4523 20715
rect 5400 20712 5428 20879
rect 6302 20876 6308 20888
rect 6360 20876 6366 20928
rect 8694 20876 8700 20928
rect 8752 20916 8758 20928
rect 9525 20919 9583 20925
rect 9525 20916 9537 20919
rect 8752 20888 9537 20916
rect 8752 20876 8758 20888
rect 9525 20885 9537 20888
rect 9571 20885 9583 20919
rect 9525 20879 9583 20885
rect 6397 20851 6455 20857
rect 6397 20817 6409 20851
rect 6443 20848 6455 20851
rect 7222 20848 7228 20860
rect 6443 20820 7228 20848
rect 6443 20817 6455 20820
rect 6397 20811 6455 20817
rect 7222 20808 7228 20820
rect 7280 20808 7286 20860
rect 8421 20851 8479 20857
rect 8421 20817 8433 20851
rect 8467 20848 8479 20851
rect 11104 20848 11132 20944
rect 11733 20851 11791 20857
rect 11733 20848 11745 20851
rect 8467 20820 9568 20848
rect 11104 20820 11745 20848
rect 8467 20817 8479 20820
rect 8421 20811 8479 20817
rect 6210 20780 6216 20792
rect 6123 20752 6216 20780
rect 6210 20740 6216 20752
rect 6268 20780 6274 20792
rect 7317 20783 7375 20789
rect 7317 20780 7329 20783
rect 6268 20752 7329 20780
rect 6268 20740 6274 20752
rect 7317 20749 7329 20752
rect 7363 20749 7375 20783
rect 7682 20780 7688 20792
rect 7643 20752 7688 20780
rect 7317 20743 7375 20749
rect 7682 20740 7688 20752
rect 7740 20740 7746 20792
rect 7866 20780 7872 20792
rect 7827 20752 7872 20780
rect 7866 20740 7872 20752
rect 7924 20740 7930 20792
rect 4511 20684 5428 20712
rect 4511 20681 4523 20684
rect 4465 20675 4523 20681
rect 7038 20672 7044 20724
rect 7096 20712 7102 20724
rect 8436 20712 8464 20811
rect 9540 20792 9568 20820
rect 11733 20817 11745 20820
rect 11779 20848 11791 20851
rect 12377 20851 12435 20857
rect 12377 20848 12389 20851
rect 11779 20820 12389 20848
rect 11779 20817 11791 20820
rect 11733 20811 11791 20817
rect 12377 20817 12389 20820
rect 12423 20848 12435 20851
rect 12650 20848 12656 20860
rect 12423 20820 12656 20848
rect 12423 20817 12435 20820
rect 12377 20811 12435 20817
rect 12650 20808 12656 20820
rect 12708 20808 12714 20860
rect 17084 20848 17112 20944
rect 21485 20919 21543 20925
rect 21485 20885 21497 20919
rect 21531 20916 21543 20919
rect 22586 20916 22592 20928
rect 21531 20888 22592 20916
rect 21531 20885 21543 20888
rect 21485 20879 21543 20885
rect 22586 20876 22592 20888
rect 22644 20876 22650 20928
rect 22770 20916 22776 20928
rect 22731 20888 22776 20916
rect 22770 20876 22776 20888
rect 22828 20876 22834 20928
rect 23156 20916 23184 20956
rect 23233 20953 23245 20987
rect 23279 20984 23291 20987
rect 23414 20984 23420 20996
rect 23279 20956 23420 20984
rect 23279 20953 23291 20956
rect 23233 20947 23291 20953
rect 23414 20944 23420 20956
rect 23472 20944 23478 20996
rect 24150 20944 24156 20996
rect 24208 20984 24214 20996
rect 24245 20987 24303 20993
rect 24245 20984 24257 20987
rect 24208 20956 24257 20984
rect 24208 20944 24214 20956
rect 24245 20953 24257 20956
rect 24291 20953 24303 20987
rect 24518 20984 24524 20996
rect 24479 20956 24524 20984
rect 24245 20947 24303 20953
rect 24518 20944 24524 20956
rect 24576 20944 24582 20996
rect 26726 20944 26732 20996
rect 26784 20984 26790 20996
rect 26821 20987 26879 20993
rect 26821 20984 26833 20987
rect 26784 20956 26833 20984
rect 26784 20944 26790 20956
rect 26821 20953 26833 20956
rect 26867 20953 26879 20987
rect 26821 20947 26879 20953
rect 27097 20987 27155 20993
rect 27097 20953 27109 20987
rect 27143 20984 27155 20987
rect 27462 20984 27468 20996
rect 27143 20956 27468 20984
rect 27143 20953 27155 20956
rect 27097 20947 27155 20953
rect 27462 20944 27468 20956
rect 27520 20944 27526 20996
rect 27646 20984 27652 20996
rect 27607 20956 27652 20984
rect 27646 20944 27652 20956
rect 27704 20944 27710 20996
rect 28017 20987 28075 20993
rect 28017 20953 28029 20987
rect 28063 20984 28075 20987
rect 29302 20984 29308 20996
rect 28063 20956 29308 20984
rect 28063 20953 28075 20956
rect 28017 20947 28075 20953
rect 29302 20944 29308 20956
rect 29360 20944 29366 20996
rect 23156 20888 23736 20916
rect 17621 20851 17679 20857
rect 17621 20848 17633 20851
rect 17084 20820 17633 20848
rect 17621 20817 17633 20820
rect 17667 20817 17679 20851
rect 17621 20811 17679 20817
rect 17710 20808 17716 20860
rect 17768 20848 17774 20860
rect 20013 20851 20071 20857
rect 20013 20848 20025 20851
rect 17768 20820 20025 20848
rect 17768 20808 17774 20820
rect 20013 20817 20025 20820
rect 20059 20848 20071 20851
rect 20657 20851 20715 20857
rect 20657 20848 20669 20851
rect 20059 20820 20669 20848
rect 20059 20817 20071 20820
rect 20013 20811 20071 20817
rect 20657 20817 20669 20820
rect 20703 20817 20715 20851
rect 20657 20811 20715 20817
rect 21669 20851 21727 20857
rect 21669 20817 21681 20851
rect 21715 20848 21727 20851
rect 23230 20848 23236 20860
rect 21715 20820 23236 20848
rect 21715 20817 21727 20820
rect 21669 20811 21727 20817
rect 23230 20808 23236 20820
rect 23288 20808 23294 20860
rect 8697 20783 8755 20789
rect 8697 20780 8709 20783
rect 7096 20684 8464 20712
rect 8528 20752 8709 20780
rect 8528 20712 8556 20752
rect 8697 20749 8709 20752
rect 8743 20749 8755 20783
rect 9062 20780 9068 20792
rect 9023 20752 9068 20780
rect 8697 20743 8755 20749
rect 9062 20740 9068 20752
rect 9120 20740 9126 20792
rect 9522 20780 9528 20792
rect 9483 20752 9528 20780
rect 9522 20740 9528 20752
rect 9580 20740 9586 20792
rect 10534 20740 10540 20792
rect 10592 20780 10598 20792
rect 10629 20783 10687 20789
rect 10629 20780 10641 20783
rect 10592 20752 10641 20780
rect 10592 20740 10598 20752
rect 10629 20749 10641 20752
rect 10675 20780 10687 20783
rect 11454 20780 11460 20792
rect 10675 20752 11460 20780
rect 10675 20749 10687 20752
rect 10629 20743 10687 20749
rect 11454 20740 11460 20752
rect 11512 20740 11518 20792
rect 11825 20783 11883 20789
rect 11825 20780 11837 20783
rect 11564 20752 11837 20780
rect 10902 20712 10908 20724
rect 8528 20684 10908 20712
rect 7096 20672 7102 20684
rect 6946 20644 6952 20656
rect 840 20616 1012 20644
rect 6907 20616 6952 20644
rect 840 20604 846 20616
rect 6946 20604 6952 20616
rect 7004 20604 7010 20656
rect 7130 20604 7136 20656
rect 7188 20644 7194 20656
rect 8528 20653 8556 20684
rect 10902 20672 10908 20684
rect 10960 20712 10966 20724
rect 11273 20715 11331 20721
rect 11273 20712 11285 20715
rect 10960 20684 11285 20712
rect 10960 20672 10966 20684
rect 11273 20681 11285 20684
rect 11319 20712 11331 20715
rect 11564 20712 11592 20752
rect 11825 20749 11837 20752
rect 11871 20780 11883 20783
rect 12561 20783 12619 20789
rect 12561 20780 12573 20783
rect 11871 20752 12573 20780
rect 11871 20749 11883 20752
rect 11825 20743 11883 20749
rect 12561 20749 12573 20752
rect 12607 20749 12619 20783
rect 12561 20743 12619 20749
rect 16977 20783 17035 20789
rect 16977 20749 16989 20783
rect 17023 20780 17035 20783
rect 17158 20780 17164 20792
rect 17023 20752 17164 20780
rect 17023 20749 17035 20752
rect 16977 20743 17035 20749
rect 17158 20740 17164 20752
rect 17216 20740 17222 20792
rect 17342 20780 17348 20792
rect 17303 20752 17348 20780
rect 17342 20740 17348 20752
rect 17400 20740 17406 20792
rect 20381 20783 20439 20789
rect 20381 20749 20393 20783
rect 20427 20780 20439 20783
rect 21853 20783 21911 20789
rect 20427 20752 21160 20780
rect 20427 20749 20439 20752
rect 20381 20743 20439 20749
rect 12285 20715 12343 20721
rect 12285 20712 12297 20715
rect 11319 20684 11592 20712
rect 11656 20684 12297 20712
rect 11319 20681 11331 20684
rect 11273 20675 11331 20681
rect 11656 20656 11684 20684
rect 12285 20681 12297 20684
rect 12331 20681 12343 20715
rect 12285 20675 12343 20681
rect 18078 20672 18084 20724
rect 18136 20672 18142 20724
rect 19366 20712 19372 20724
rect 19279 20684 19372 20712
rect 19366 20672 19372 20684
rect 19424 20712 19430 20724
rect 20197 20715 20255 20721
rect 20197 20712 20209 20715
rect 19424 20684 20209 20712
rect 19424 20672 19430 20684
rect 20197 20681 20209 20684
rect 20243 20712 20255 20715
rect 20841 20715 20899 20721
rect 20841 20712 20853 20715
rect 20243 20684 20853 20712
rect 20243 20681 20255 20684
rect 20197 20675 20255 20681
rect 20841 20681 20853 20684
rect 20887 20681 20899 20715
rect 20841 20675 20899 20681
rect 8513 20647 8571 20653
rect 8513 20644 8525 20647
rect 7188 20616 8525 20644
rect 7188 20604 7194 20616
rect 8513 20613 8525 20616
rect 8559 20613 8571 20647
rect 8513 20607 8571 20613
rect 9798 20604 9804 20656
rect 9856 20644 9862 20656
rect 10258 20644 10264 20656
rect 9856 20616 10264 20644
rect 9856 20604 9862 20616
rect 10258 20604 10264 20616
rect 10316 20644 10322 20656
rect 10353 20647 10411 20653
rect 10353 20644 10365 20647
rect 10316 20616 10365 20644
rect 10316 20604 10322 20616
rect 10353 20613 10365 20616
rect 10399 20644 10411 20647
rect 10810 20644 10816 20656
rect 10399 20616 10816 20644
rect 10399 20613 10411 20616
rect 10353 20607 10411 20613
rect 10810 20604 10816 20616
rect 10868 20604 10874 20656
rect 10997 20647 11055 20653
rect 10997 20613 11009 20647
rect 11043 20644 11055 20647
rect 11178 20644 11184 20656
rect 11043 20616 11184 20644
rect 11043 20613 11055 20616
rect 10997 20607 11055 20613
rect 11178 20604 11184 20616
rect 11236 20604 11242 20656
rect 11549 20647 11607 20653
rect 11549 20613 11561 20647
rect 11595 20644 11607 20647
rect 11638 20644 11644 20656
rect 11595 20616 11644 20644
rect 11595 20613 11607 20616
rect 11549 20607 11607 20613
rect 11638 20604 11644 20616
rect 11696 20604 11702 20656
rect 16514 20644 16520 20656
rect 16475 20616 16520 20644
rect 16514 20604 16520 20616
rect 16572 20604 16578 20656
rect 21132 20653 21160 20752
rect 21853 20749 21865 20783
rect 21899 20780 21911 20783
rect 22862 20780 22868 20792
rect 21899 20752 22868 20780
rect 21899 20749 21911 20752
rect 21853 20743 21911 20749
rect 22862 20740 22868 20752
rect 22920 20740 22926 20792
rect 23414 20780 23420 20792
rect 23375 20752 23420 20780
rect 23414 20740 23420 20752
rect 23472 20740 23478 20792
rect 23598 20780 23604 20792
rect 23559 20752 23604 20780
rect 23598 20740 23604 20752
rect 23656 20740 23662 20792
rect 22310 20712 22316 20724
rect 22271 20684 22316 20712
rect 22310 20672 22316 20684
rect 22368 20672 22374 20724
rect 21117 20647 21175 20653
rect 21117 20613 21129 20647
rect 21163 20644 21175 20647
rect 22126 20644 22132 20656
rect 21163 20616 22132 20644
rect 21163 20613 21175 20616
rect 21117 20607 21175 20613
rect 22126 20604 22132 20616
rect 22184 20604 22190 20656
rect 23708 20644 23736 20888
rect 27554 20876 27560 20928
rect 27612 20916 27618 20928
rect 27833 20919 27891 20925
rect 27833 20916 27845 20919
rect 27612 20888 27845 20916
rect 27612 20876 27618 20888
rect 27833 20885 27845 20888
rect 27879 20916 27891 20919
rect 28474 20916 28480 20928
rect 27879 20888 28480 20916
rect 27879 20885 27891 20888
rect 27833 20879 27891 20885
rect 28474 20876 28480 20888
rect 28532 20876 28538 20928
rect 23782 20808 23788 20860
rect 23840 20848 23846 20860
rect 23877 20851 23935 20857
rect 23877 20848 23889 20851
rect 23840 20820 23889 20848
rect 23840 20808 23846 20820
rect 23877 20817 23889 20820
rect 23923 20817 23935 20851
rect 23877 20811 23935 20817
rect 27002 20808 27008 20860
rect 27060 20848 27066 20860
rect 27373 20851 27431 20857
rect 27373 20848 27385 20851
rect 27060 20820 27385 20848
rect 27060 20808 27066 20820
rect 27373 20817 27385 20820
rect 27419 20817 27431 20851
rect 28566 20848 28572 20860
rect 28527 20820 28572 20848
rect 27373 20811 27431 20817
rect 28566 20808 28572 20820
rect 28624 20808 28630 20860
rect 23969 20783 24027 20789
rect 23969 20749 23981 20783
rect 24015 20749 24027 20783
rect 23969 20743 24027 20749
rect 23984 20712 24012 20743
rect 24610 20740 24616 20792
rect 24668 20780 24674 20792
rect 24981 20783 25039 20789
rect 24981 20780 24993 20783
rect 24668 20752 24993 20780
rect 24668 20740 24674 20752
rect 24981 20749 24993 20752
rect 25027 20780 25039 20783
rect 25625 20783 25683 20789
rect 25625 20780 25637 20783
rect 25027 20752 25637 20780
rect 25027 20749 25039 20752
rect 24981 20743 25039 20749
rect 25625 20749 25637 20752
rect 25671 20780 25683 20783
rect 27281 20783 27339 20789
rect 27281 20780 27293 20783
rect 25671 20752 27293 20780
rect 25671 20749 25683 20752
rect 25625 20743 25683 20749
rect 27281 20749 27293 20752
rect 27327 20780 27339 20783
rect 27738 20780 27744 20792
rect 27327 20752 27744 20780
rect 27327 20749 27339 20752
rect 27281 20743 27339 20749
rect 27738 20740 27744 20752
rect 27796 20740 27802 20792
rect 25257 20715 25315 20721
rect 25257 20712 25269 20715
rect 23846 20684 25269 20712
rect 23846 20644 23874 20684
rect 25257 20681 25269 20684
rect 25303 20712 25315 20715
rect 25809 20715 25867 20721
rect 25809 20712 25821 20715
rect 25303 20684 25821 20712
rect 25303 20681 25315 20684
rect 25257 20675 25315 20681
rect 25809 20681 25821 20684
rect 25855 20712 25867 20715
rect 25990 20712 25996 20724
rect 25855 20684 25996 20712
rect 25855 20681 25867 20684
rect 25809 20675 25867 20681
rect 25990 20672 25996 20684
rect 26048 20712 26054 20724
rect 27646 20712 27652 20724
rect 26048 20684 27652 20712
rect 26048 20672 26054 20684
rect 27646 20672 27652 20684
rect 27704 20672 27710 20724
rect 28845 20715 28903 20721
rect 28845 20712 28857 20715
rect 28124 20684 28857 20712
rect 28124 20656 28152 20684
rect 28845 20681 28857 20684
rect 28891 20681 28903 20715
rect 28845 20675 28903 20681
rect 29302 20672 29308 20724
rect 29360 20672 29366 20724
rect 30593 20715 30651 20721
rect 30593 20681 30605 20715
rect 30639 20681 30651 20715
rect 30593 20675 30651 20681
rect 28106 20644 28112 20656
rect 23708 20616 23874 20644
rect 28067 20616 28112 20644
rect 28106 20604 28112 20616
rect 28164 20604 28170 20656
rect 28290 20644 28296 20656
rect 28251 20616 28296 20644
rect 28290 20604 28296 20616
rect 28348 20644 28354 20656
rect 30608 20644 30636 20675
rect 28348 20616 30636 20644
rect 28348 20604 28354 20616
rect 400 20554 31680 20576
rect 400 20502 18870 20554
rect 18922 20502 18934 20554
rect 18986 20502 18998 20554
rect 19050 20502 19062 20554
rect 19114 20502 19126 20554
rect 19178 20502 31680 20554
rect 400 20480 31680 20502
rect 1245 20443 1303 20449
rect 1245 20409 1257 20443
rect 1291 20440 1303 20443
rect 1426 20440 1432 20452
rect 1291 20412 1432 20440
rect 1291 20409 1303 20412
rect 1245 20403 1303 20409
rect 1426 20400 1432 20412
rect 1484 20400 1490 20452
rect 2073 20443 2131 20449
rect 2073 20409 2085 20443
rect 2119 20440 2131 20443
rect 2622 20440 2628 20452
rect 2119 20412 2628 20440
rect 2119 20409 2131 20412
rect 2073 20403 2131 20409
rect 2622 20400 2628 20412
rect 2680 20400 2686 20452
rect 5750 20400 5756 20452
rect 5808 20440 5814 20452
rect 5937 20443 5995 20449
rect 5937 20440 5949 20443
rect 5808 20412 5949 20440
rect 5808 20400 5814 20412
rect 5937 20409 5949 20412
rect 5983 20409 5995 20443
rect 8694 20440 8700 20452
rect 8655 20412 8700 20440
rect 5937 20403 5995 20409
rect 8694 20400 8700 20412
rect 8752 20400 8758 20452
rect 9062 20400 9068 20452
rect 9120 20440 9126 20452
rect 9525 20443 9583 20449
rect 9525 20440 9537 20443
rect 9120 20412 9537 20440
rect 9120 20400 9126 20412
rect 9525 20409 9537 20412
rect 9571 20409 9583 20443
rect 9525 20403 9583 20409
rect 16514 20400 16520 20452
rect 16572 20440 16578 20452
rect 16572 20412 16836 20440
rect 16572 20400 16578 20412
rect 1334 20372 1340 20384
rect 1295 20344 1340 20372
rect 1334 20332 1340 20344
rect 1392 20332 1398 20384
rect 7774 20372 7780 20384
rect 7735 20344 7780 20372
rect 7774 20332 7780 20344
rect 7832 20332 7838 20384
rect 14677 20375 14735 20381
rect 9264 20344 11040 20372
rect 9264 20316 9292 20344
rect 2714 20264 2720 20316
rect 2772 20304 2778 20316
rect 3174 20304 3180 20316
rect 2772 20276 3180 20304
rect 2772 20264 2778 20276
rect 3174 20264 3180 20276
rect 3232 20304 3238 20316
rect 3361 20307 3419 20313
rect 3361 20304 3373 20307
rect 3232 20276 3373 20304
rect 3232 20264 3238 20276
rect 3361 20273 3373 20276
rect 3407 20273 3419 20307
rect 3361 20267 3419 20273
rect 5845 20307 5903 20313
rect 5845 20273 5857 20307
rect 5891 20304 5903 20307
rect 6394 20304 6400 20316
rect 5891 20276 6400 20304
rect 5891 20273 5903 20276
rect 5845 20267 5903 20273
rect 6394 20264 6400 20276
rect 6452 20264 6458 20316
rect 7038 20304 7044 20316
rect 6999 20276 7044 20304
rect 7038 20264 7044 20276
rect 7096 20264 7102 20316
rect 7188 20307 7246 20313
rect 7188 20273 7200 20307
rect 7234 20304 7246 20307
rect 7314 20304 7320 20316
rect 7234 20276 7320 20304
rect 7234 20273 7246 20276
rect 7188 20267 7246 20273
rect 7314 20264 7320 20276
rect 7372 20264 7378 20316
rect 9246 20304 9252 20316
rect 9207 20276 9252 20304
rect 9246 20264 9252 20276
rect 9304 20264 9310 20316
rect 11012 20313 11040 20344
rect 14677 20341 14689 20375
rect 14723 20372 14735 20375
rect 14950 20372 14956 20384
rect 14723 20344 14956 20372
rect 14723 20341 14735 20344
rect 14677 20335 14735 20341
rect 14950 20332 14956 20344
rect 15008 20332 15014 20384
rect 16808 20381 16836 20412
rect 17066 20400 17072 20452
rect 17124 20440 17130 20452
rect 17345 20443 17403 20449
rect 17345 20440 17357 20443
rect 17124 20412 17357 20440
rect 17124 20400 17130 20412
rect 17345 20409 17357 20412
rect 17391 20409 17403 20443
rect 17345 20403 17403 20409
rect 23049 20443 23107 20449
rect 23049 20409 23061 20443
rect 23095 20440 23107 20443
rect 23414 20440 23420 20452
rect 23095 20412 23420 20440
rect 23095 20409 23107 20412
rect 23049 20403 23107 20409
rect 23414 20400 23420 20412
rect 23472 20400 23478 20452
rect 27186 20400 27192 20452
rect 27244 20440 27250 20452
rect 28382 20440 28388 20452
rect 27244 20412 28388 20440
rect 27244 20400 27250 20412
rect 28382 20400 28388 20412
rect 28440 20400 28446 20452
rect 16793 20375 16851 20381
rect 16793 20341 16805 20375
rect 16839 20341 16851 20375
rect 16793 20335 16851 20341
rect 17621 20375 17679 20381
rect 17621 20341 17633 20375
rect 17667 20372 17679 20375
rect 18078 20372 18084 20384
rect 17667 20344 18084 20372
rect 17667 20341 17679 20344
rect 17621 20335 17679 20341
rect 18078 20332 18084 20344
rect 18136 20332 18142 20384
rect 20933 20375 20991 20381
rect 20933 20341 20945 20375
rect 20979 20372 20991 20375
rect 21390 20372 21396 20384
rect 20979 20344 21396 20372
rect 20979 20341 20991 20344
rect 20933 20335 20991 20341
rect 21390 20332 21396 20344
rect 21448 20372 21454 20384
rect 21758 20372 21764 20384
rect 21448 20344 21764 20372
rect 21448 20332 21454 20344
rect 21758 20332 21764 20344
rect 21816 20332 21822 20384
rect 21850 20332 21856 20384
rect 21908 20372 21914 20384
rect 23141 20375 23199 20381
rect 23141 20372 23153 20375
rect 21908 20344 23153 20372
rect 21908 20332 21914 20344
rect 23141 20341 23153 20344
rect 23187 20372 23199 20375
rect 23598 20372 23604 20384
rect 23187 20344 23604 20372
rect 23187 20341 23199 20344
rect 23141 20335 23199 20341
rect 23598 20332 23604 20344
rect 23656 20332 23662 20384
rect 28014 20372 28020 20384
rect 27664 20344 28020 20372
rect 9433 20307 9491 20313
rect 9433 20273 9445 20307
rect 9479 20273 9491 20307
rect 9433 20267 9491 20273
rect 10997 20307 11055 20313
rect 10997 20273 11009 20307
rect 11043 20304 11055 20307
rect 11178 20304 11184 20316
rect 11043 20276 11184 20304
rect 11043 20273 11055 20276
rect 10997 20267 11055 20273
rect 6670 20196 6676 20248
rect 6728 20236 6734 20248
rect 7409 20239 7467 20245
rect 7409 20236 7421 20239
rect 6728 20208 7421 20236
rect 6728 20196 6734 20208
rect 7409 20205 7421 20208
rect 7455 20205 7467 20239
rect 7409 20199 7467 20205
rect 8970 20196 8976 20248
rect 9028 20236 9034 20248
rect 9448 20236 9476 20267
rect 11178 20264 11184 20276
rect 11236 20264 11242 20316
rect 11638 20304 11644 20316
rect 11599 20276 11644 20304
rect 11638 20264 11644 20276
rect 11696 20264 11702 20316
rect 16422 20264 16428 20316
rect 16480 20304 16486 20316
rect 16517 20307 16575 20313
rect 16517 20304 16529 20307
rect 16480 20276 16529 20304
rect 16480 20264 16486 20276
rect 16517 20273 16529 20276
rect 16563 20273 16575 20307
rect 17069 20307 17127 20313
rect 17069 20304 17081 20307
rect 16517 20267 16575 20273
rect 16624 20276 17081 20304
rect 11086 20236 11092 20248
rect 9028 20208 9476 20236
rect 11047 20208 11092 20236
rect 9028 20196 9034 20208
rect 11086 20196 11092 20208
rect 11144 20196 11150 20248
rect 11730 20236 11736 20248
rect 11691 20208 11736 20236
rect 11730 20196 11736 20208
rect 11788 20196 11794 20248
rect 11822 20196 11828 20248
rect 11880 20236 11886 20248
rect 16624 20236 16652 20276
rect 17069 20273 17081 20276
rect 17115 20304 17127 20307
rect 17434 20304 17440 20316
rect 17115 20276 17440 20304
rect 17115 20273 17127 20276
rect 17069 20267 17127 20273
rect 17434 20264 17440 20276
rect 17492 20264 17498 20316
rect 17802 20304 17808 20316
rect 17763 20276 17808 20304
rect 17802 20264 17808 20276
rect 17860 20264 17866 20316
rect 21022 20264 21028 20316
rect 21080 20304 21086 20316
rect 21577 20307 21635 20313
rect 21577 20304 21589 20307
rect 21080 20276 21589 20304
rect 21080 20264 21086 20276
rect 21577 20273 21589 20276
rect 21623 20273 21635 20307
rect 21577 20267 21635 20273
rect 21666 20264 21672 20316
rect 21724 20304 21730 20316
rect 21945 20307 22003 20313
rect 21945 20304 21957 20307
rect 21724 20276 21957 20304
rect 21724 20264 21730 20276
rect 21945 20273 21957 20276
rect 21991 20273 22003 20307
rect 21945 20267 22003 20273
rect 23230 20264 23236 20316
rect 23288 20304 23294 20316
rect 26542 20304 26548 20316
rect 23288 20276 26548 20304
rect 23288 20264 23294 20276
rect 26542 20264 26548 20276
rect 26600 20304 26606 20316
rect 27370 20304 27376 20316
rect 26600 20276 27376 20304
rect 26600 20264 26606 20276
rect 27370 20264 27376 20276
rect 27428 20264 27434 20316
rect 27664 20313 27692 20344
rect 28014 20332 28020 20344
rect 28072 20372 28078 20384
rect 28842 20372 28848 20384
rect 28072 20344 28848 20372
rect 28072 20332 28078 20344
rect 28842 20332 28848 20344
rect 28900 20332 28906 20384
rect 27649 20307 27707 20313
rect 27649 20273 27661 20307
rect 27695 20273 27707 20307
rect 27830 20304 27836 20316
rect 27791 20276 27836 20304
rect 27649 20267 27707 20273
rect 27830 20264 27836 20276
rect 27888 20264 27894 20316
rect 28382 20313 28388 20316
rect 28109 20307 28167 20313
rect 28109 20273 28121 20307
rect 28155 20273 28167 20307
rect 28109 20267 28167 20273
rect 28362 20307 28388 20313
rect 28362 20273 28374 20307
rect 28362 20267 28388 20273
rect 21485 20239 21543 20245
rect 21485 20236 21497 20239
rect 11880 20208 16652 20236
rect 20764 20208 21497 20236
rect 11880 20196 11886 20208
rect 690 20128 696 20180
rect 748 20168 754 20180
rect 969 20171 1027 20177
rect 969 20168 981 20171
rect 748 20140 981 20168
rect 748 20128 754 20140
rect 969 20137 981 20140
rect 1015 20168 1027 20171
rect 6854 20168 6860 20180
rect 1015 20140 6860 20168
rect 1015 20137 1027 20140
rect 969 20131 1027 20137
rect 6854 20128 6860 20140
rect 6912 20128 6918 20180
rect 7314 20168 7320 20180
rect 7227 20140 7320 20168
rect 7314 20128 7320 20140
rect 7372 20168 7378 20180
rect 11362 20168 11368 20180
rect 7372 20140 11368 20168
rect 7372 20128 7378 20140
rect 11362 20128 11368 20140
rect 11420 20128 11426 20180
rect 12006 20168 12012 20180
rect 11967 20140 12012 20168
rect 12006 20128 12012 20140
rect 12064 20128 12070 20180
rect 12190 20128 12196 20180
rect 12248 20168 12254 20180
rect 14674 20168 14680 20180
rect 12248 20140 14680 20168
rect 12248 20128 12254 20140
rect 14674 20128 14680 20140
rect 14732 20168 14738 20180
rect 14953 20171 15011 20177
rect 14953 20168 14965 20171
rect 14732 20140 14965 20168
rect 14732 20128 14738 20140
rect 14953 20137 14965 20140
rect 14999 20168 15011 20171
rect 17342 20168 17348 20180
rect 14999 20140 17348 20168
rect 14999 20137 15011 20140
rect 14953 20131 15011 20137
rect 17342 20128 17348 20140
rect 17400 20128 17406 20180
rect 20764 20112 20792 20208
rect 21485 20205 21497 20208
rect 21531 20205 21543 20239
rect 22034 20236 22040 20248
rect 21995 20208 22040 20236
rect 21485 20199 21543 20205
rect 22034 20196 22040 20208
rect 22092 20196 22098 20248
rect 27462 20196 27468 20248
rect 27520 20236 27526 20248
rect 28124 20236 28152 20267
rect 28382 20264 28388 20267
rect 28440 20264 28446 20316
rect 27520 20208 28152 20236
rect 27520 20196 27526 20208
rect 28124 20168 28152 20208
rect 28198 20196 28204 20248
rect 28256 20236 28262 20248
rect 28661 20239 28719 20245
rect 28661 20236 28673 20239
rect 28256 20208 28673 20236
rect 28256 20196 28262 20208
rect 28661 20205 28673 20208
rect 28707 20205 28719 20239
rect 28661 20199 28719 20205
rect 29486 20196 29492 20248
rect 29544 20236 29550 20248
rect 30130 20236 30136 20248
rect 29544 20208 30136 20236
rect 29544 20196 29550 20208
rect 30130 20196 30136 20208
rect 30188 20196 30194 20248
rect 28290 20168 28296 20180
rect 28124 20140 28296 20168
rect 28290 20128 28296 20140
rect 28348 20128 28354 20180
rect 782 20100 788 20112
rect 743 20072 788 20100
rect 782 20060 788 20072
rect 840 20060 846 20112
rect 3266 20060 3272 20112
rect 3324 20100 3330 20112
rect 3453 20103 3511 20109
rect 3453 20100 3465 20103
rect 3324 20072 3465 20100
rect 3324 20060 3330 20072
rect 3453 20069 3465 20072
rect 3499 20069 3511 20103
rect 3453 20063 3511 20069
rect 4830 20060 4836 20112
rect 4888 20100 4894 20112
rect 6765 20103 6823 20109
rect 6765 20100 6777 20103
rect 4888 20072 6777 20100
rect 4888 20060 4894 20072
rect 6765 20069 6777 20072
rect 6811 20100 6823 20103
rect 7682 20100 7688 20112
rect 6811 20072 7688 20100
rect 6811 20069 6823 20072
rect 6765 20063 6823 20069
rect 7682 20060 7688 20072
rect 7740 20100 7746 20112
rect 7961 20103 8019 20109
rect 7961 20100 7973 20103
rect 7740 20072 7973 20100
rect 7740 20060 7746 20072
rect 7961 20069 7973 20072
rect 8007 20100 8019 20103
rect 8142 20100 8148 20112
rect 8007 20072 8148 20100
rect 8007 20069 8019 20072
rect 7961 20063 8019 20069
rect 8142 20060 8148 20072
rect 8200 20060 8206 20112
rect 9798 20060 9804 20112
rect 9856 20100 9862 20112
rect 9893 20103 9951 20109
rect 9893 20100 9905 20103
rect 9856 20072 9905 20100
rect 9856 20060 9862 20072
rect 9893 20069 9905 20072
rect 9939 20069 9951 20103
rect 12098 20100 12104 20112
rect 12059 20072 12104 20100
rect 9893 20063 9951 20069
rect 12098 20060 12104 20072
rect 12156 20060 12162 20112
rect 20289 20103 20347 20109
rect 20289 20069 20301 20103
rect 20335 20100 20347 20103
rect 20746 20100 20752 20112
rect 20335 20072 20752 20100
rect 20335 20069 20347 20072
rect 20289 20063 20347 20069
rect 20746 20060 20752 20072
rect 20804 20060 20810 20112
rect 400 20010 31680 20032
rect 400 19958 3510 20010
rect 3562 19958 3574 20010
rect 3626 19958 3638 20010
rect 3690 19958 3702 20010
rect 3754 19958 3766 20010
rect 3818 19958 31680 20010
rect 400 19936 31680 19958
rect 1150 19896 1156 19908
rect 1111 19868 1156 19896
rect 1150 19856 1156 19868
rect 1208 19896 1214 19908
rect 1245 19899 1303 19905
rect 1245 19896 1257 19899
rect 1208 19868 1257 19896
rect 1208 19856 1214 19868
rect 1245 19865 1257 19868
rect 1291 19865 1303 19899
rect 1245 19859 1303 19865
rect 3174 19856 3180 19908
rect 3232 19896 3238 19908
rect 3453 19899 3511 19905
rect 3453 19896 3465 19899
rect 3232 19868 3465 19896
rect 3232 19856 3238 19868
rect 3453 19865 3465 19868
rect 3499 19865 3511 19899
rect 3453 19859 3511 19865
rect 6302 19856 6308 19908
rect 6360 19896 6366 19908
rect 6489 19899 6547 19905
rect 6489 19896 6501 19899
rect 6360 19868 6501 19896
rect 6360 19856 6366 19868
rect 6489 19865 6501 19868
rect 6535 19865 6547 19899
rect 7222 19896 7228 19908
rect 7183 19868 7228 19896
rect 6489 19859 6547 19865
rect 7222 19856 7228 19868
rect 7280 19856 7286 19908
rect 9246 19896 9252 19908
rect 9207 19868 9252 19896
rect 9246 19856 9252 19868
rect 9304 19856 9310 19908
rect 9798 19896 9804 19908
rect 9759 19868 9804 19896
rect 9798 19856 9804 19868
rect 9856 19856 9862 19908
rect 10350 19856 10356 19908
rect 10408 19896 10414 19908
rect 10905 19899 10963 19905
rect 10408 19868 10856 19896
rect 10408 19856 10414 19868
rect 782 19788 788 19840
rect 840 19828 846 19840
rect 1889 19831 1947 19837
rect 1889 19828 1901 19831
rect 840 19800 1901 19828
rect 840 19788 846 19800
rect 1889 19797 1901 19800
rect 1935 19828 1947 19831
rect 2349 19831 2407 19837
rect 2349 19828 2361 19831
rect 1935 19800 2361 19828
rect 1935 19797 1947 19800
rect 1889 19791 1947 19797
rect 2349 19797 2361 19800
rect 2395 19797 2407 19831
rect 2349 19791 2407 19797
rect 7133 19831 7191 19837
rect 7133 19797 7145 19831
rect 7179 19828 7191 19831
rect 7314 19828 7320 19840
rect 7179 19800 7320 19828
rect 7179 19797 7191 19800
rect 7133 19791 7191 19797
rect 7314 19788 7320 19800
rect 7372 19788 7378 19840
rect 7409 19831 7467 19837
rect 7409 19797 7421 19831
rect 7455 19828 7467 19831
rect 7866 19828 7872 19840
rect 7455 19800 7872 19828
rect 7455 19797 7467 19800
rect 7409 19791 7467 19797
rect 7866 19788 7872 19800
rect 7924 19828 7930 19840
rect 8881 19831 8939 19837
rect 7924 19800 8464 19828
rect 7924 19788 7930 19800
rect 8436 19769 8464 19800
rect 8881 19797 8893 19831
rect 8927 19828 8939 19831
rect 9522 19828 9528 19840
rect 8927 19800 9528 19828
rect 8927 19797 8939 19800
rect 8881 19791 8939 19797
rect 9522 19788 9528 19800
rect 9580 19828 9586 19840
rect 9580 19800 10580 19828
rect 9580 19788 9586 19800
rect 1521 19763 1579 19769
rect 1521 19729 1533 19763
rect 1567 19760 1579 19763
rect 8421 19763 8479 19769
rect 8421 19760 8433 19763
rect 1567 19732 3220 19760
rect 8142 19734 8148 19746
rect 1567 19729 1579 19732
rect 1521 19723 1579 19729
rect 1705 19695 1763 19701
rect 1705 19661 1717 19695
rect 1751 19692 1763 19695
rect 2349 19695 2407 19701
rect 2349 19692 2361 19695
rect 1751 19664 2361 19692
rect 1751 19661 1763 19664
rect 1705 19655 1763 19661
rect 2349 19661 2361 19664
rect 2395 19661 2407 19695
rect 2622 19692 2628 19704
rect 2583 19664 2628 19692
rect 2349 19655 2407 19661
rect 2364 19624 2392 19655
rect 2622 19652 2628 19664
rect 2680 19652 2686 19704
rect 2714 19652 2720 19704
rect 2772 19692 2778 19704
rect 3192 19701 3220 19732
rect 8097 19706 8148 19734
rect 2901 19695 2959 19701
rect 2901 19692 2913 19695
rect 2772 19664 2913 19692
rect 2772 19652 2778 19664
rect 2901 19661 2913 19664
rect 2947 19661 2959 19695
rect 2901 19655 2959 19661
rect 3177 19695 3235 19701
rect 3177 19661 3189 19695
rect 3223 19692 3235 19695
rect 3358 19692 3364 19704
rect 3223 19664 3364 19692
rect 3223 19661 3235 19664
rect 3177 19655 3235 19661
rect 3358 19652 3364 19664
rect 3416 19652 3422 19704
rect 6670 19652 6676 19704
rect 6728 19692 6734 19704
rect 6857 19695 6915 19701
rect 6857 19692 6869 19695
rect 6728 19664 6869 19692
rect 6728 19652 6734 19664
rect 6857 19661 6869 19664
rect 6903 19661 6915 19695
rect 6857 19655 6915 19661
rect 7406 19652 7412 19704
rect 7464 19692 7470 19704
rect 7961 19695 8019 19701
rect 7961 19692 7973 19695
rect 7464 19664 7973 19692
rect 7464 19652 7470 19664
rect 7961 19661 7973 19664
rect 8007 19661 8019 19695
rect 8142 19694 8148 19706
rect 8200 19694 8206 19746
rect 8344 19732 8433 19760
rect 7961 19655 8019 19661
rect 8145 19661 8157 19694
rect 8191 19661 8203 19694
rect 8145 19655 8203 19661
rect 3266 19624 3272 19636
rect 2364 19596 3272 19624
rect 3266 19584 3272 19596
rect 3324 19624 3330 19636
rect 3637 19627 3695 19633
rect 3637 19624 3649 19627
rect 3324 19596 3649 19624
rect 3324 19584 3330 19596
rect 3637 19593 3649 19596
rect 3683 19593 3695 19627
rect 3637 19587 3695 19593
rect 6765 19627 6823 19633
rect 6765 19593 6777 19627
rect 6811 19624 6823 19627
rect 7130 19624 7136 19636
rect 6811 19596 7136 19624
rect 6811 19593 6823 19596
rect 6765 19587 6823 19593
rect 7130 19584 7136 19596
rect 7188 19624 7194 19636
rect 7225 19627 7283 19633
rect 7225 19624 7237 19627
rect 7188 19596 7237 19624
rect 7188 19584 7194 19596
rect 7225 19593 7237 19596
rect 7271 19593 7283 19627
rect 8344 19624 8372 19732
rect 8421 19729 8433 19732
rect 8467 19729 8479 19763
rect 8421 19723 8479 19729
rect 8528 19732 10212 19760
rect 8528 19704 8556 19732
rect 10184 19704 10212 19732
rect 10350 19720 10356 19772
rect 10408 19760 10414 19772
rect 10445 19763 10503 19769
rect 10445 19760 10457 19763
rect 10408 19732 10457 19760
rect 10408 19720 10414 19732
rect 10445 19729 10457 19732
rect 10491 19729 10503 19763
rect 10445 19723 10503 19729
rect 8510 19692 8516 19704
rect 8423 19664 8516 19692
rect 8510 19652 8516 19664
rect 8568 19652 8574 19704
rect 9341 19695 9399 19701
rect 9341 19692 9353 19695
rect 8896 19664 9353 19692
rect 8896 19624 8924 19664
rect 9341 19661 9353 19664
rect 9387 19692 9399 19695
rect 9522 19692 9528 19704
rect 9387 19664 9528 19692
rect 9387 19661 9399 19664
rect 9341 19655 9399 19661
rect 9522 19652 9528 19664
rect 9580 19652 9586 19704
rect 9982 19692 9988 19704
rect 9943 19664 9988 19692
rect 9982 19652 9988 19664
rect 10040 19652 10046 19704
rect 10166 19692 10172 19704
rect 10127 19664 10172 19692
rect 10166 19652 10172 19664
rect 10224 19652 10230 19704
rect 10552 19701 10580 19800
rect 10828 19760 10856 19868
rect 10905 19865 10917 19899
rect 10951 19896 10963 19899
rect 12006 19896 12012 19908
rect 10951 19868 12012 19896
rect 10951 19865 10963 19868
rect 10905 19859 10963 19865
rect 12006 19856 12012 19868
rect 12064 19856 12070 19908
rect 12193 19899 12251 19905
rect 12193 19865 12205 19899
rect 12239 19896 12251 19899
rect 12282 19896 12288 19908
rect 12239 19868 12288 19896
rect 12239 19865 12251 19868
rect 12193 19859 12251 19865
rect 12282 19856 12288 19868
rect 12340 19856 12346 19908
rect 14674 19896 14680 19908
rect 14635 19868 14680 19896
rect 14674 19856 14680 19868
rect 14732 19856 14738 19908
rect 14861 19899 14919 19905
rect 14861 19865 14873 19899
rect 14907 19896 14919 19899
rect 14950 19896 14956 19908
rect 14907 19868 14956 19896
rect 14907 19865 14919 19868
rect 14861 19859 14919 19865
rect 14950 19856 14956 19868
rect 15008 19856 15014 19908
rect 16514 19856 16520 19908
rect 16572 19896 16578 19908
rect 16701 19899 16759 19905
rect 16701 19896 16713 19899
rect 16572 19868 16713 19896
rect 16572 19856 16578 19868
rect 16701 19865 16713 19868
rect 16747 19865 16759 19899
rect 16701 19859 16759 19865
rect 17897 19899 17955 19905
rect 17897 19865 17909 19899
rect 17943 19896 17955 19899
rect 18078 19896 18084 19908
rect 17943 19868 18084 19896
rect 17943 19865 17955 19868
rect 17897 19859 17955 19865
rect 18078 19856 18084 19868
rect 18136 19856 18142 19908
rect 19737 19899 19795 19905
rect 19737 19865 19749 19899
rect 19783 19896 19795 19899
rect 20289 19899 20347 19905
rect 20289 19896 20301 19899
rect 19783 19868 20301 19896
rect 19783 19865 19795 19868
rect 19737 19859 19795 19865
rect 20289 19865 20301 19868
rect 20335 19896 20347 19899
rect 21850 19896 21856 19908
rect 20335 19868 21856 19896
rect 20335 19865 20347 19868
rect 20289 19859 20347 19865
rect 21850 19856 21856 19868
rect 21908 19856 21914 19908
rect 23693 19899 23751 19905
rect 23693 19865 23705 19899
rect 23739 19896 23751 19899
rect 24150 19896 24156 19908
rect 23739 19868 24156 19896
rect 23739 19865 23751 19868
rect 23693 19859 23751 19865
rect 11178 19828 11184 19840
rect 11139 19800 11184 19828
rect 11178 19788 11184 19800
rect 11236 19788 11242 19840
rect 17802 19788 17808 19840
rect 17860 19828 17866 19840
rect 17989 19831 18047 19837
rect 17989 19828 18001 19831
rect 17860 19800 18001 19828
rect 17860 19788 17866 19800
rect 17989 19797 18001 19800
rect 18035 19797 18047 19831
rect 17989 19791 18047 19797
rect 18538 19788 18544 19840
rect 18596 19828 18602 19840
rect 19918 19828 19924 19840
rect 18596 19800 19924 19828
rect 18596 19788 18602 19800
rect 19918 19788 19924 19800
rect 19976 19828 19982 19840
rect 20013 19831 20071 19837
rect 20013 19828 20025 19831
rect 19976 19800 20025 19828
rect 19976 19788 19982 19800
rect 20013 19797 20025 19800
rect 20059 19828 20071 19831
rect 21206 19828 21212 19840
rect 20059 19800 21212 19828
rect 20059 19797 20071 19800
rect 20013 19791 20071 19797
rect 21206 19788 21212 19800
rect 21264 19788 21270 19840
rect 21577 19831 21635 19837
rect 21577 19797 21589 19831
rect 21623 19828 21635 19831
rect 21666 19828 21672 19840
rect 21623 19800 21672 19828
rect 21623 19797 21635 19800
rect 21577 19791 21635 19797
rect 21666 19788 21672 19800
rect 21724 19788 21730 19840
rect 12561 19763 12619 19769
rect 12561 19760 12573 19763
rect 10828 19732 12573 19760
rect 10537 19695 10595 19701
rect 10537 19661 10549 19695
rect 10583 19661 10595 19695
rect 11086 19692 11092 19704
rect 11047 19664 11092 19692
rect 10537 19655 10595 19661
rect 11086 19652 11092 19664
rect 11144 19652 11150 19704
rect 11730 19692 11736 19704
rect 11643 19664 11736 19692
rect 11730 19652 11736 19664
rect 11788 19652 11794 19704
rect 11932 19701 11960 19732
rect 12561 19729 12573 19732
rect 12607 19729 12619 19763
rect 20746 19760 20752 19772
rect 20707 19732 20752 19760
rect 12561 19723 12619 19729
rect 20746 19720 20752 19732
rect 20804 19760 20810 19772
rect 22681 19763 22739 19769
rect 22681 19760 22693 19763
rect 20804 19732 22693 19760
rect 20804 19720 20810 19732
rect 22681 19729 22693 19732
rect 22727 19760 22739 19763
rect 23417 19763 23475 19769
rect 23417 19760 23429 19763
rect 22727 19732 23429 19760
rect 22727 19729 22739 19732
rect 22681 19723 22739 19729
rect 23417 19729 23429 19732
rect 23463 19729 23475 19763
rect 23417 19723 23475 19729
rect 11917 19695 11975 19701
rect 11917 19661 11929 19695
rect 11963 19661 11975 19695
rect 11917 19655 11975 19661
rect 12009 19695 12067 19701
rect 12009 19661 12021 19695
rect 12055 19692 12067 19695
rect 12098 19692 12104 19704
rect 12055 19664 12104 19692
rect 12055 19661 12067 19664
rect 12009 19655 12067 19661
rect 12098 19652 12104 19664
rect 12156 19652 12162 19704
rect 12374 19652 12380 19704
rect 12432 19692 12438 19704
rect 12834 19692 12840 19704
rect 12432 19664 12840 19692
rect 12432 19652 12438 19664
rect 12834 19652 12840 19664
rect 12892 19692 12898 19704
rect 13297 19695 13355 19701
rect 13297 19692 13309 19695
rect 12892 19664 13309 19692
rect 12892 19652 12898 19664
rect 13297 19661 13309 19664
rect 13343 19692 13355 19695
rect 13757 19695 13815 19701
rect 13757 19692 13769 19695
rect 13343 19664 13769 19692
rect 13343 19661 13355 19664
rect 13297 19655 13355 19661
rect 13757 19661 13769 19664
rect 13803 19661 13815 19695
rect 13757 19655 13815 19661
rect 20286 19652 20292 19704
rect 20344 19692 20350 19704
rect 20841 19695 20899 19701
rect 20841 19692 20853 19695
rect 20344 19664 20853 19692
rect 20344 19652 20350 19664
rect 20841 19661 20853 19664
rect 20887 19661 20899 19695
rect 21206 19692 21212 19704
rect 21167 19664 21212 19692
rect 20841 19655 20899 19661
rect 21206 19652 21212 19664
rect 21264 19652 21270 19704
rect 21301 19695 21359 19701
rect 21301 19661 21313 19695
rect 21347 19661 21359 19695
rect 21301 19655 21359 19661
rect 23141 19695 23199 19701
rect 23141 19661 23153 19695
rect 23187 19692 23199 19695
rect 23708 19692 23736 19859
rect 24150 19856 24156 19868
rect 24208 19856 24214 19908
rect 27186 19896 27192 19908
rect 27147 19868 27192 19896
rect 27186 19856 27192 19868
rect 27244 19856 27250 19908
rect 27649 19899 27707 19905
rect 27649 19865 27661 19899
rect 27695 19896 27707 19899
rect 28106 19896 28112 19908
rect 27695 19868 28112 19896
rect 27695 19865 27707 19868
rect 27649 19859 27707 19865
rect 28106 19856 28112 19868
rect 28164 19856 28170 19908
rect 27370 19788 27376 19840
rect 27428 19828 27434 19840
rect 27741 19831 27799 19837
rect 27741 19828 27753 19831
rect 27428 19800 27753 19828
rect 27428 19788 27434 19800
rect 27741 19797 27753 19800
rect 27787 19797 27799 19831
rect 28014 19828 28020 19840
rect 27975 19800 28020 19828
rect 27741 19791 27799 19797
rect 28014 19788 28020 19800
rect 28072 19788 28078 19840
rect 28566 19720 28572 19772
rect 28624 19760 28630 19772
rect 28845 19763 28903 19769
rect 28845 19760 28857 19763
rect 28624 19732 28857 19760
rect 28624 19720 28630 19732
rect 28845 19729 28857 19732
rect 28891 19760 28903 19763
rect 29397 19763 29455 19769
rect 29397 19760 29409 19763
rect 28891 19732 29409 19760
rect 28891 19729 28903 19732
rect 28845 19723 28903 19729
rect 29397 19729 29409 19732
rect 29443 19729 29455 19763
rect 29397 19723 29455 19729
rect 23187 19664 23736 19692
rect 23187 19661 23199 19664
rect 23141 19655 23199 19661
rect 11365 19627 11423 19633
rect 11365 19624 11377 19627
rect 8344 19596 8924 19624
rect 8988 19596 11377 19624
rect 7225 19587 7283 19593
rect 8988 19568 9016 19596
rect 11365 19593 11377 19596
rect 11411 19624 11423 19627
rect 11748 19624 11776 19652
rect 11411 19596 11776 19624
rect 11411 19593 11423 19596
rect 11365 19587 11423 19593
rect 12926 19584 12932 19636
rect 12984 19624 12990 19636
rect 13665 19627 13723 19633
rect 13665 19624 13677 19627
rect 12984 19596 13677 19624
rect 12984 19584 12990 19596
rect 13665 19593 13677 19596
rect 13711 19624 13723 19627
rect 13941 19627 13999 19633
rect 13941 19624 13953 19627
rect 13711 19596 13953 19624
rect 13711 19593 13723 19596
rect 13665 19587 13723 19593
rect 13941 19593 13953 19596
rect 13987 19593 13999 19627
rect 21316 19624 21344 19655
rect 27922 19652 27928 19704
rect 27980 19692 27986 19704
rect 28661 19695 28719 19701
rect 28661 19692 28673 19695
rect 27980 19664 28673 19692
rect 27980 19652 27986 19664
rect 28661 19661 28673 19664
rect 28707 19692 28719 19695
rect 29213 19695 29271 19701
rect 29213 19692 29225 19695
rect 28707 19664 29225 19692
rect 28707 19661 28719 19664
rect 28661 19655 28719 19661
rect 29213 19661 29225 19664
rect 29259 19661 29271 19695
rect 29213 19655 29271 19661
rect 21669 19627 21727 19633
rect 21669 19624 21681 19627
rect 13941 19587 13999 19593
rect 19844 19596 21681 19624
rect 19844 19568 19872 19596
rect 21669 19593 21681 19596
rect 21715 19624 21727 19627
rect 22034 19624 22040 19636
rect 21715 19596 22040 19624
rect 21715 19593 21727 19596
rect 21669 19587 21727 19593
rect 22034 19584 22040 19596
rect 22092 19584 22098 19636
rect 22957 19627 23015 19633
rect 22957 19593 22969 19627
rect 23003 19593 23015 19627
rect 22957 19587 23015 19593
rect 7777 19559 7835 19565
rect 7777 19525 7789 19559
rect 7823 19556 7835 19559
rect 7866 19556 7872 19568
rect 7823 19528 7872 19556
rect 7823 19525 7835 19528
rect 7777 19519 7835 19525
rect 7866 19516 7872 19528
rect 7924 19516 7930 19568
rect 8970 19556 8976 19568
rect 8931 19528 8976 19556
rect 8970 19516 8976 19528
rect 9028 19516 9034 19568
rect 9522 19516 9528 19568
rect 9580 19556 9586 19568
rect 10350 19556 10356 19568
rect 9580 19528 10356 19556
rect 9580 19516 9586 19528
rect 10350 19516 10356 19528
rect 10408 19516 10414 19568
rect 16422 19516 16428 19568
rect 16480 19556 16486 19568
rect 16609 19559 16667 19565
rect 16609 19556 16621 19559
rect 16480 19528 16621 19556
rect 16480 19516 16486 19528
rect 16609 19525 16621 19528
rect 16655 19556 16667 19559
rect 18078 19556 18084 19568
rect 16655 19528 18084 19556
rect 16655 19525 16667 19528
rect 16609 19519 16667 19525
rect 18078 19516 18084 19528
rect 18136 19516 18142 19568
rect 19826 19556 19832 19568
rect 19787 19528 19832 19556
rect 19826 19516 19832 19528
rect 19884 19516 19890 19568
rect 20194 19516 20200 19568
rect 20252 19556 20258 19568
rect 22972 19556 23000 19587
rect 26726 19584 26732 19636
rect 26784 19624 26790 19636
rect 27830 19624 27836 19636
rect 26784 19596 27836 19624
rect 26784 19584 26790 19596
rect 27830 19584 27836 19596
rect 27888 19624 27894 19636
rect 28109 19627 28167 19633
rect 28109 19624 28121 19627
rect 27888 19596 28121 19624
rect 27888 19584 27894 19596
rect 28109 19593 28121 19596
rect 28155 19593 28167 19627
rect 28109 19587 28167 19593
rect 23785 19559 23843 19565
rect 23785 19556 23797 19559
rect 20252 19528 23797 19556
rect 20252 19516 20258 19528
rect 23785 19525 23797 19528
rect 23831 19556 23843 19559
rect 26450 19556 26456 19568
rect 23831 19528 26456 19556
rect 23831 19525 23843 19528
rect 23785 19519 23843 19525
rect 26450 19516 26456 19528
rect 26508 19516 26514 19568
rect 27370 19556 27376 19568
rect 27331 19528 27376 19556
rect 27370 19516 27376 19528
rect 27428 19516 27434 19568
rect 400 19466 31680 19488
rect 400 19414 18870 19466
rect 18922 19414 18934 19466
rect 18986 19414 18998 19466
rect 19050 19414 19062 19466
rect 19114 19414 19126 19466
rect 19178 19414 31680 19466
rect 400 19392 31680 19414
rect 1886 19312 1892 19364
rect 1944 19352 1950 19364
rect 1981 19355 2039 19361
rect 1981 19352 1993 19355
rect 1944 19324 1993 19352
rect 1944 19312 1950 19324
rect 1981 19321 1993 19324
rect 2027 19352 2039 19355
rect 2622 19352 2628 19364
rect 2027 19324 2628 19352
rect 2027 19321 2039 19324
rect 1981 19315 2039 19321
rect 2622 19312 2628 19324
rect 2680 19312 2686 19364
rect 7038 19352 7044 19364
rect 6999 19324 7044 19352
rect 7038 19312 7044 19324
rect 7096 19312 7102 19364
rect 7590 19352 7596 19364
rect 7503 19324 7596 19352
rect 7590 19312 7596 19324
rect 7648 19352 7654 19364
rect 8510 19352 8516 19364
rect 7648 19324 8516 19352
rect 7648 19312 7654 19324
rect 8510 19312 8516 19324
rect 8568 19312 8574 19364
rect 9062 19312 9068 19364
rect 9120 19352 9126 19364
rect 9249 19355 9307 19361
rect 9249 19352 9261 19355
rect 9120 19324 9261 19352
rect 9120 19312 9126 19324
rect 9249 19321 9261 19324
rect 9295 19321 9307 19355
rect 9249 19315 9307 19321
rect 9617 19355 9675 19361
rect 9617 19321 9629 19355
rect 9663 19352 9675 19355
rect 10166 19352 10172 19364
rect 9663 19324 10172 19352
rect 9663 19321 9675 19324
rect 9617 19315 9675 19321
rect 10166 19312 10172 19324
rect 10224 19312 10230 19364
rect 10813 19355 10871 19361
rect 10813 19321 10825 19355
rect 10859 19352 10871 19355
rect 11638 19352 11644 19364
rect 10859 19324 11644 19352
rect 10859 19321 10871 19324
rect 10813 19315 10871 19321
rect 11638 19312 11644 19324
rect 11696 19312 11702 19364
rect 11730 19312 11736 19364
rect 11788 19352 11794 19364
rect 11917 19355 11975 19361
rect 11917 19352 11929 19355
rect 11788 19324 11929 19352
rect 11788 19312 11794 19324
rect 11917 19321 11929 19324
rect 11963 19321 11975 19355
rect 11917 19315 11975 19321
rect 12193 19355 12251 19361
rect 12193 19321 12205 19355
rect 12239 19352 12251 19355
rect 12282 19352 12288 19364
rect 12239 19324 12288 19352
rect 12239 19321 12251 19324
rect 12193 19315 12251 19321
rect 12282 19312 12288 19324
rect 12340 19312 12346 19364
rect 17802 19352 17808 19364
rect 15520 19324 17808 19352
rect 2714 19244 2720 19296
rect 2772 19284 2778 19296
rect 3266 19284 3272 19296
rect 2772 19256 3272 19284
rect 2772 19244 2778 19256
rect 3266 19244 3272 19256
rect 3324 19284 3330 19296
rect 3637 19287 3695 19293
rect 3637 19284 3649 19287
rect 3324 19256 3649 19284
rect 3324 19244 3330 19256
rect 3637 19253 3649 19256
rect 3683 19253 3695 19287
rect 3637 19247 3695 19253
rect 5382 19244 5388 19296
rect 5440 19284 5446 19296
rect 6486 19284 6492 19296
rect 5440 19256 6492 19284
rect 5440 19244 5446 19256
rect 6486 19244 6492 19256
rect 6544 19284 6550 19296
rect 6581 19287 6639 19293
rect 6581 19284 6593 19287
rect 6544 19256 6593 19284
rect 6544 19244 6550 19256
rect 6581 19253 6593 19256
rect 6627 19253 6639 19287
rect 6581 19247 6639 19253
rect 7406 19244 7412 19296
rect 7464 19284 7470 19296
rect 7685 19287 7743 19293
rect 7685 19284 7697 19287
rect 7464 19256 7697 19284
rect 7464 19244 7470 19256
rect 7685 19253 7697 19256
rect 7731 19284 7743 19287
rect 9709 19287 9767 19293
rect 9709 19284 9721 19287
rect 7731 19256 9721 19284
rect 7731 19253 7743 19256
rect 7685 19247 7743 19253
rect 9709 19253 9721 19256
rect 9755 19284 9767 19287
rect 9982 19284 9988 19296
rect 9755 19256 9988 19284
rect 9755 19253 9767 19256
rect 9709 19247 9767 19253
rect 9982 19244 9988 19256
rect 10040 19244 10046 19296
rect 11825 19287 11883 19293
rect 11825 19253 11837 19287
rect 11871 19284 11883 19287
rect 12098 19284 12104 19296
rect 11871 19256 12104 19284
rect 11871 19253 11883 19256
rect 11825 19247 11883 19253
rect 12098 19244 12104 19256
rect 12156 19244 12162 19296
rect 12742 19244 12748 19296
rect 12800 19284 12806 19296
rect 15226 19284 15232 19296
rect 12800 19256 13156 19284
rect 12800 19244 12806 19256
rect 3358 19216 3364 19228
rect 3271 19188 3364 19216
rect 3358 19176 3364 19188
rect 3416 19216 3422 19228
rect 4830 19216 4836 19228
rect 3416 19188 4836 19216
rect 3416 19176 3422 19188
rect 4830 19176 4836 19188
rect 4888 19216 4894 19228
rect 5017 19219 5075 19225
rect 5017 19216 5029 19219
rect 4888 19188 5029 19216
rect 4888 19176 4894 19188
rect 5017 19185 5029 19188
rect 5063 19185 5075 19219
rect 6302 19216 6308 19228
rect 6215 19188 6308 19216
rect 5017 19179 5075 19185
rect 6302 19176 6308 19188
rect 6360 19216 6366 19228
rect 7424 19216 7452 19244
rect 7866 19216 7872 19228
rect 6360 19188 7452 19216
rect 7827 19188 7872 19216
rect 6360 19176 6366 19188
rect 7866 19176 7872 19188
rect 7924 19176 7930 19228
rect 10534 19216 10540 19228
rect 10495 19188 10540 19216
rect 10534 19176 10540 19188
rect 10592 19176 10598 19228
rect 11546 19216 11552 19228
rect 11507 19188 11552 19216
rect 11546 19176 11552 19188
rect 11604 19176 11610 19228
rect 12834 19176 12840 19228
rect 12892 19216 12898 19228
rect 13128 19225 13156 19256
rect 14876 19256 15232 19284
rect 14876 19225 14904 19256
rect 15226 19244 15232 19256
rect 15284 19284 15290 19296
rect 15520 19284 15548 19324
rect 17802 19312 17808 19324
rect 17860 19312 17866 19364
rect 20286 19352 20292 19364
rect 20247 19324 20292 19352
rect 20286 19312 20292 19324
rect 20344 19312 20350 19364
rect 20746 19312 20752 19364
rect 20804 19352 20810 19364
rect 20933 19355 20991 19361
rect 20933 19352 20945 19355
rect 20804 19324 20945 19352
rect 20804 19312 20810 19324
rect 20933 19321 20945 19324
rect 20979 19321 20991 19355
rect 21390 19352 21396 19364
rect 21351 19324 21396 19352
rect 20933 19315 20991 19321
rect 21390 19312 21396 19324
rect 21448 19312 21454 19364
rect 23325 19355 23383 19361
rect 23325 19321 23337 19355
rect 23371 19352 23383 19355
rect 23414 19352 23420 19364
rect 23371 19324 23420 19352
rect 23371 19321 23383 19324
rect 23325 19315 23383 19321
rect 23414 19312 23420 19324
rect 23472 19312 23478 19364
rect 16882 19284 16888 19296
rect 15284 19256 15548 19284
rect 16795 19256 16888 19284
rect 15284 19244 15290 19256
rect 16882 19244 16888 19256
rect 16940 19284 16946 19296
rect 20304 19284 20332 19312
rect 16940 19256 20332 19284
rect 16940 19244 16946 19256
rect 28198 19244 28204 19296
rect 28256 19284 28262 19296
rect 28658 19284 28664 19296
rect 28256 19256 28664 19284
rect 28256 19244 28262 19256
rect 28658 19244 28664 19256
rect 28716 19284 28722 19296
rect 28937 19287 28995 19293
rect 28937 19284 28949 19287
rect 28716 19256 28949 19284
rect 28716 19244 28722 19256
rect 28937 19253 28949 19256
rect 28983 19284 28995 19287
rect 29394 19284 29400 19296
rect 28983 19256 29400 19284
rect 28983 19253 28995 19256
rect 28937 19247 28995 19253
rect 29394 19244 29400 19256
rect 29452 19244 29458 19296
rect 12929 19219 12987 19225
rect 12929 19216 12941 19219
rect 12892 19188 12941 19216
rect 12892 19176 12898 19188
rect 12929 19185 12941 19188
rect 12975 19185 12987 19219
rect 12929 19179 12987 19185
rect 13113 19219 13171 19225
rect 13113 19185 13125 19219
rect 13159 19185 13171 19219
rect 13113 19179 13171 19185
rect 14861 19219 14919 19225
rect 14861 19185 14873 19219
rect 14907 19185 14919 19219
rect 16146 19216 16152 19228
rect 16107 19188 16152 19216
rect 14861 19179 14919 19185
rect 16146 19176 16152 19188
rect 16204 19176 16210 19228
rect 16606 19216 16612 19228
rect 16567 19188 16612 19216
rect 16606 19176 16612 19188
rect 16664 19176 16670 19228
rect 20654 19176 20660 19228
rect 20712 19216 20718 19228
rect 21945 19219 22003 19225
rect 21945 19216 21957 19219
rect 20712 19188 21957 19216
rect 20712 19176 20718 19188
rect 21945 19185 21957 19188
rect 21991 19216 22003 19219
rect 22034 19216 22040 19228
rect 21991 19188 22040 19216
rect 21991 19185 22003 19188
rect 21945 19179 22003 19185
rect 22034 19176 22040 19188
rect 22092 19176 22098 19228
rect 23230 19216 23236 19228
rect 23191 19188 23236 19216
rect 23230 19176 23236 19188
rect 23288 19176 23294 19228
rect 26910 19176 26916 19228
rect 26968 19216 26974 19228
rect 27922 19216 27928 19228
rect 26968 19188 27928 19216
rect 26968 19176 26974 19188
rect 27922 19176 27928 19188
rect 27980 19176 27986 19228
rect 29118 19216 29124 19228
rect 29079 19188 29124 19216
rect 29118 19176 29124 19188
rect 29176 19176 29182 19228
rect 30498 19216 30504 19228
rect 30459 19188 30504 19216
rect 30498 19176 30504 19188
rect 30556 19176 30562 19228
rect 5290 19148 5296 19160
rect 5251 19120 5296 19148
rect 5290 19108 5296 19120
rect 5348 19108 5354 19160
rect 7884 19148 7912 19176
rect 11730 19148 11736 19160
rect 7884 19120 11736 19148
rect 11730 19108 11736 19120
rect 11788 19108 11794 19160
rect 13478 19148 13484 19160
rect 13439 19120 13484 19148
rect 13478 19108 13484 19120
rect 13536 19108 13542 19160
rect 15042 19148 15048 19160
rect 15003 19120 15048 19148
rect 15042 19108 15048 19120
rect 15100 19108 15106 19160
rect 22126 19148 22132 19160
rect 22087 19120 22132 19148
rect 22126 19108 22132 19120
rect 22184 19108 22190 19160
rect 26726 19108 26732 19160
rect 26784 19148 26790 19160
rect 27097 19151 27155 19157
rect 27097 19148 27109 19151
rect 26784 19120 27109 19148
rect 26784 19108 26790 19120
rect 27097 19117 27109 19120
rect 27143 19117 27155 19151
rect 27646 19148 27652 19160
rect 27607 19120 27652 19148
rect 27097 19111 27155 19117
rect 27646 19108 27652 19120
rect 27704 19108 27710 19160
rect 28106 19148 28112 19160
rect 28067 19120 28112 19148
rect 28106 19108 28112 19120
rect 28164 19148 28170 19160
rect 28569 19151 28627 19157
rect 28569 19148 28581 19151
rect 28164 19120 28581 19148
rect 28164 19108 28170 19120
rect 28569 19117 28581 19120
rect 28615 19117 28627 19151
rect 28569 19111 28627 19117
rect 29489 19151 29547 19157
rect 29489 19117 29501 19151
rect 29535 19148 29547 19151
rect 29578 19148 29584 19160
rect 29535 19120 29584 19148
rect 29535 19117 29547 19120
rect 29489 19111 29547 19117
rect 29578 19108 29584 19120
rect 29636 19108 29642 19160
rect 5308 19080 5336 19108
rect 10258 19080 10264 19092
rect 5308 19052 10264 19080
rect 10258 19040 10264 19052
rect 10316 19040 10322 19092
rect 10350 19012 10356 19024
rect 10311 18984 10356 19012
rect 10350 18972 10356 18984
rect 10408 18972 10414 19024
rect 21022 18972 21028 19024
rect 21080 19012 21086 19024
rect 21117 19015 21175 19021
rect 21117 19012 21129 19015
rect 21080 18984 21129 19012
rect 21080 18972 21086 18984
rect 21117 18981 21129 18984
rect 21163 18981 21175 19015
rect 21117 18975 21175 18981
rect 23877 19015 23935 19021
rect 23877 18981 23889 19015
rect 23923 19012 23935 19015
rect 24150 19012 24156 19024
rect 23923 18984 24156 19012
rect 23923 18981 23935 18984
rect 23877 18975 23935 18981
rect 24150 18972 24156 18984
rect 24208 18972 24214 19024
rect 24702 18972 24708 19024
rect 24760 19012 24766 19024
rect 25162 19012 25168 19024
rect 24760 18984 25168 19012
rect 24760 18972 24766 18984
rect 25162 18972 25168 18984
rect 25220 18972 25226 19024
rect 400 18922 31680 18944
rect 400 18870 3510 18922
rect 3562 18870 3574 18922
rect 3626 18870 3638 18922
rect 3690 18870 3702 18922
rect 3754 18870 3766 18922
rect 3818 18870 31680 18922
rect 400 18848 31680 18870
rect 3358 18808 3364 18820
rect 3319 18780 3364 18808
rect 3358 18768 3364 18780
rect 3416 18768 3422 18820
rect 5290 18808 5296 18820
rect 5251 18780 5296 18808
rect 5290 18768 5296 18780
rect 5348 18768 5354 18820
rect 6302 18808 6308 18820
rect 6263 18780 6308 18808
rect 6302 18768 6308 18780
rect 6360 18768 6366 18820
rect 6486 18808 6492 18820
rect 6447 18780 6492 18808
rect 6486 18768 6492 18780
rect 6544 18768 6550 18820
rect 10353 18811 10411 18817
rect 10353 18777 10365 18811
rect 10399 18808 10411 18811
rect 10534 18808 10540 18820
rect 10399 18780 10540 18808
rect 10399 18777 10411 18780
rect 10353 18771 10411 18777
rect 10534 18768 10540 18780
rect 10592 18768 10598 18820
rect 11270 18808 11276 18820
rect 11231 18780 11276 18808
rect 11270 18768 11276 18780
rect 11328 18768 11334 18820
rect 11546 18808 11552 18820
rect 11507 18780 11552 18808
rect 11546 18768 11552 18780
rect 11604 18768 11610 18820
rect 12098 18768 12104 18820
rect 12156 18808 12162 18820
rect 12285 18811 12343 18817
rect 12285 18808 12297 18811
rect 12156 18780 12297 18808
rect 12156 18768 12162 18780
rect 12285 18777 12297 18780
rect 12331 18808 12343 18811
rect 12469 18811 12527 18817
rect 12469 18808 12481 18811
rect 12331 18780 12481 18808
rect 12331 18777 12343 18780
rect 12285 18771 12343 18777
rect 12469 18777 12481 18780
rect 12515 18777 12527 18811
rect 12469 18771 12527 18777
rect 12742 18768 12748 18820
rect 12800 18808 12806 18820
rect 12837 18811 12895 18817
rect 12837 18808 12849 18811
rect 12800 18780 12849 18808
rect 12800 18768 12806 18780
rect 12837 18777 12849 18780
rect 12883 18777 12895 18811
rect 12837 18771 12895 18777
rect 13478 18768 13484 18820
rect 13536 18808 13542 18820
rect 13849 18811 13907 18817
rect 13849 18808 13861 18811
rect 13536 18780 13861 18808
rect 13536 18768 13542 18780
rect 13849 18777 13861 18780
rect 13895 18777 13907 18811
rect 14953 18811 15011 18817
rect 14953 18808 14965 18811
rect 13849 18771 13907 18777
rect 14186 18780 14965 18808
rect 3266 18700 3272 18752
rect 3324 18740 3330 18752
rect 3545 18743 3603 18749
rect 3545 18740 3557 18743
rect 3324 18712 3557 18740
rect 3324 18700 3330 18712
rect 3545 18709 3557 18712
rect 3591 18709 3603 18743
rect 3545 18703 3603 18709
rect 9798 18700 9804 18752
rect 9856 18740 9862 18752
rect 9856 18712 13064 18740
rect 9856 18700 9862 18712
rect 5474 18632 5480 18684
rect 5532 18672 5538 18684
rect 8970 18672 8976 18684
rect 5532 18644 8976 18672
rect 5532 18632 5538 18644
rect 8970 18632 8976 18644
rect 9028 18672 9034 18684
rect 9249 18675 9307 18681
rect 9249 18672 9261 18675
rect 9028 18644 9261 18672
rect 9028 18632 9034 18644
rect 9249 18641 9261 18644
rect 9295 18672 9307 18675
rect 9893 18675 9951 18681
rect 9893 18672 9905 18675
rect 9295 18644 9905 18672
rect 9295 18641 9307 18644
rect 9249 18635 9307 18641
rect 9893 18641 9905 18644
rect 9939 18641 9951 18675
rect 9893 18635 9951 18641
rect 11270 18632 11276 18684
rect 11328 18672 11334 18684
rect 11917 18675 11975 18681
rect 11917 18672 11929 18675
rect 11328 18644 11929 18672
rect 11328 18632 11334 18644
rect 11917 18641 11929 18644
rect 11963 18641 11975 18675
rect 11917 18635 11975 18641
rect 12745 18675 12803 18681
rect 12745 18641 12757 18675
rect 12791 18672 12803 18675
rect 12834 18672 12840 18684
rect 12791 18644 12840 18672
rect 12791 18641 12803 18644
rect 12745 18635 12803 18641
rect 12834 18632 12840 18644
rect 12892 18632 12898 18684
rect 6670 18564 6676 18616
rect 6728 18604 6734 18616
rect 9065 18607 9123 18613
rect 9065 18604 9077 18607
rect 6728 18576 9077 18604
rect 6728 18564 6734 18576
rect 9065 18573 9077 18576
rect 9111 18604 9123 18607
rect 9617 18607 9675 18613
rect 9617 18604 9629 18607
rect 9111 18576 9629 18604
rect 9111 18573 9123 18576
rect 9065 18567 9123 18573
rect 9617 18573 9629 18576
rect 9663 18604 9675 18607
rect 10350 18604 10356 18616
rect 9663 18576 10356 18604
rect 9663 18573 9675 18576
rect 9617 18567 9675 18573
rect 10350 18564 10356 18576
rect 10408 18604 10414 18616
rect 10445 18607 10503 18613
rect 10445 18604 10457 18607
rect 10408 18576 10457 18604
rect 10408 18564 10414 18576
rect 10445 18573 10457 18576
rect 10491 18573 10503 18607
rect 10445 18567 10503 18573
rect 11733 18607 11791 18613
rect 11733 18573 11745 18607
rect 11779 18604 11791 18607
rect 12098 18604 12104 18616
rect 11779 18576 12104 18604
rect 11779 18573 11791 18576
rect 11733 18567 11791 18573
rect 12098 18564 12104 18576
rect 12156 18564 12162 18616
rect 13036 18613 13064 18712
rect 13021 18607 13079 18613
rect 13021 18573 13033 18607
rect 13067 18604 13079 18607
rect 13110 18604 13116 18616
rect 13067 18576 13116 18604
rect 13067 18573 13079 18576
rect 13021 18567 13079 18573
rect 13110 18564 13116 18576
rect 13168 18604 13174 18616
rect 13481 18607 13539 18613
rect 13481 18604 13493 18607
rect 13168 18576 13493 18604
rect 13168 18564 13174 18576
rect 13481 18573 13493 18576
rect 13527 18573 13539 18607
rect 13481 18567 13539 18573
rect 5934 18536 5940 18548
rect 4526 18508 5940 18536
rect 1610 18428 1616 18480
rect 1668 18468 1674 18480
rect 4526 18468 4554 18508
rect 5934 18496 5940 18508
rect 5992 18496 5998 18548
rect 13389 18539 13447 18545
rect 13389 18505 13401 18539
rect 13435 18536 13447 18539
rect 13662 18536 13668 18548
rect 13435 18508 13668 18536
rect 13435 18505 13447 18508
rect 13389 18499 13447 18505
rect 13662 18496 13668 18508
rect 13720 18496 13726 18548
rect 1668 18440 4554 18468
rect 1668 18428 1674 18440
rect 4830 18428 4836 18480
rect 4888 18468 4894 18480
rect 5017 18471 5075 18477
rect 5017 18468 5029 18471
rect 4888 18440 5029 18468
rect 4888 18428 4894 18440
rect 5017 18437 5029 18440
rect 5063 18437 5075 18471
rect 13864 18468 13892 18771
rect 13938 18632 13944 18684
rect 13996 18672 14002 18684
rect 14186 18672 14214 18780
rect 14953 18777 14965 18780
rect 14999 18808 15011 18811
rect 15042 18808 15048 18820
rect 14999 18780 15048 18808
rect 14999 18777 15011 18780
rect 14953 18771 15011 18777
rect 15042 18768 15048 18780
rect 15100 18768 15106 18820
rect 15137 18811 15195 18817
rect 15137 18777 15149 18811
rect 15183 18808 15195 18811
rect 15226 18808 15232 18820
rect 15183 18780 15232 18808
rect 15183 18777 15195 18780
rect 15137 18771 15195 18777
rect 15226 18768 15232 18780
rect 15284 18768 15290 18820
rect 16146 18808 16152 18820
rect 16107 18780 16152 18808
rect 16146 18768 16152 18780
rect 16204 18768 16210 18820
rect 16609 18811 16667 18817
rect 16609 18777 16621 18811
rect 16655 18808 16667 18811
rect 16882 18808 16888 18820
rect 16655 18780 16888 18808
rect 16655 18777 16667 18780
rect 16609 18771 16667 18777
rect 16882 18768 16888 18780
rect 16940 18768 16946 18820
rect 23230 18808 23236 18820
rect 23191 18780 23236 18808
rect 23230 18768 23236 18780
rect 23288 18768 23294 18820
rect 23506 18808 23512 18820
rect 23467 18780 23512 18808
rect 23506 18768 23512 18780
rect 23564 18808 23570 18820
rect 25898 18808 25904 18820
rect 23564 18780 25904 18808
rect 23564 18768 23570 18780
rect 25898 18768 25904 18780
rect 25956 18768 25962 18820
rect 26726 18808 26732 18820
rect 26687 18780 26732 18808
rect 26726 18768 26732 18780
rect 26784 18768 26790 18820
rect 26910 18808 26916 18820
rect 26871 18780 26916 18808
rect 26910 18768 26916 18780
rect 26968 18768 26974 18820
rect 27097 18811 27155 18817
rect 27097 18777 27109 18811
rect 27143 18808 27155 18811
rect 28106 18808 28112 18820
rect 27143 18780 28112 18808
rect 27143 18777 27155 18780
rect 27097 18771 27155 18777
rect 28106 18768 28112 18780
rect 28164 18808 28170 18820
rect 28845 18811 28903 18817
rect 28845 18808 28857 18811
rect 28164 18780 28857 18808
rect 28164 18768 28170 18780
rect 28845 18777 28857 18780
rect 28891 18777 28903 18811
rect 28845 18771 28903 18777
rect 29118 18768 29124 18820
rect 29176 18808 29182 18820
rect 29486 18808 29492 18820
rect 29176 18780 29492 18808
rect 29176 18768 29182 18780
rect 29486 18768 29492 18780
rect 29544 18768 29550 18820
rect 29578 18768 29584 18820
rect 29636 18808 29642 18820
rect 29765 18811 29823 18817
rect 29765 18808 29777 18811
rect 29636 18780 29777 18808
rect 29636 18768 29642 18780
rect 29765 18777 29777 18780
rect 29811 18777 29823 18811
rect 29765 18771 29823 18777
rect 30409 18811 30467 18817
rect 30409 18777 30421 18811
rect 30455 18808 30467 18811
rect 30498 18808 30504 18820
rect 30455 18780 30504 18808
rect 30455 18777 30467 18780
rect 30409 18771 30467 18777
rect 30498 18768 30504 18780
rect 30556 18768 30562 18820
rect 14674 18700 14680 18752
rect 14732 18740 14738 18752
rect 23141 18743 23199 18749
rect 14732 18712 18124 18740
rect 14732 18700 14738 18712
rect 17989 18675 18047 18681
rect 17989 18672 18001 18675
rect 13996 18644 14214 18672
rect 17544 18644 18001 18672
rect 13996 18632 14002 18644
rect 15226 18564 15232 18616
rect 15284 18604 15290 18616
rect 16698 18604 16704 18616
rect 15284 18576 16704 18604
rect 15284 18564 15290 18576
rect 16698 18564 16704 18576
rect 16756 18604 16762 18616
rect 17544 18613 17572 18644
rect 17989 18641 18001 18644
rect 18035 18641 18047 18675
rect 18096 18672 18124 18712
rect 23141 18709 23153 18743
rect 23187 18740 23199 18743
rect 23414 18740 23420 18752
rect 23187 18712 23420 18740
rect 23187 18709 23199 18712
rect 23141 18703 23199 18709
rect 23414 18700 23420 18712
rect 23472 18700 23478 18752
rect 27646 18740 27652 18752
rect 27607 18712 27652 18740
rect 27646 18700 27652 18712
rect 27704 18700 27710 18752
rect 27925 18743 27983 18749
rect 27925 18709 27937 18743
rect 27971 18740 27983 18743
rect 28198 18740 28204 18752
rect 27971 18712 28204 18740
rect 27971 18709 27983 18712
rect 27925 18703 27983 18709
rect 28198 18700 28204 18712
rect 28256 18700 28262 18752
rect 29026 18740 29032 18752
rect 28584 18712 29032 18740
rect 24150 18672 24156 18684
rect 18096 18644 24012 18672
rect 24111 18644 24156 18672
rect 17989 18635 18047 18641
rect 17529 18607 17587 18613
rect 17529 18604 17541 18607
rect 16756 18576 17541 18604
rect 16756 18564 16762 18576
rect 17529 18573 17541 18576
rect 17575 18573 17587 18607
rect 18173 18607 18231 18613
rect 18173 18604 18185 18607
rect 17529 18567 17587 18573
rect 17636 18576 18185 18604
rect 17345 18539 17403 18545
rect 17345 18536 17357 18539
rect 17084 18508 17357 18536
rect 17084 18480 17112 18508
rect 17345 18505 17357 18508
rect 17391 18536 17403 18539
rect 17636 18536 17664 18576
rect 18173 18573 18185 18576
rect 18219 18573 18231 18607
rect 22034 18604 22040 18616
rect 21995 18576 22040 18604
rect 18173 18567 18231 18573
rect 22034 18564 22040 18576
rect 22092 18564 22098 18616
rect 23782 18604 23788 18616
rect 23743 18576 23788 18604
rect 23782 18564 23788 18576
rect 23840 18564 23846 18616
rect 23984 18604 24012 18644
rect 24150 18632 24156 18644
rect 24208 18632 24214 18684
rect 28584 18681 28612 18712
rect 29026 18700 29032 18712
rect 29084 18740 29090 18752
rect 29213 18743 29271 18749
rect 29213 18740 29225 18743
rect 29084 18712 29225 18740
rect 29084 18700 29090 18712
rect 29213 18709 29225 18712
rect 29259 18709 29271 18743
rect 29213 18703 29271 18709
rect 28569 18675 28627 18681
rect 28569 18672 28581 18675
rect 24260 18644 28581 18672
rect 24260 18604 24288 18644
rect 28569 18641 28581 18644
rect 28615 18641 28627 18675
rect 28569 18635 28627 18641
rect 29394 18632 29400 18684
rect 29452 18672 29458 18684
rect 29581 18675 29639 18681
rect 29581 18672 29593 18675
rect 29452 18644 29593 18672
rect 29452 18632 29458 18644
rect 29581 18641 29593 18644
rect 29627 18641 29639 18675
rect 29581 18635 29639 18641
rect 27465 18607 27523 18613
rect 27465 18604 27477 18607
rect 23984 18576 24288 18604
rect 25272 18576 27477 18604
rect 17391 18508 17664 18536
rect 17897 18539 17955 18545
rect 17391 18505 17403 18508
rect 17345 18499 17403 18505
rect 17897 18505 17909 18539
rect 17943 18536 17955 18539
rect 17943 18508 23874 18536
rect 17943 18505 17955 18508
rect 17897 18499 17955 18505
rect 14582 18468 14588 18480
rect 13864 18440 14588 18468
rect 5017 18431 5075 18437
rect 14582 18428 14588 18440
rect 14640 18428 14646 18480
rect 16425 18471 16483 18477
rect 16425 18437 16437 18471
rect 16471 18468 16483 18471
rect 16606 18468 16612 18480
rect 16471 18440 16612 18468
rect 16471 18437 16483 18440
rect 16425 18431 16483 18437
rect 16606 18428 16612 18440
rect 16664 18468 16670 18480
rect 17066 18468 17072 18480
rect 16664 18440 17072 18468
rect 16664 18428 16670 18440
rect 17066 18428 17072 18440
rect 17124 18428 17130 18480
rect 17161 18471 17219 18477
rect 17161 18437 17173 18471
rect 17207 18468 17219 18471
rect 17912 18468 17940 18499
rect 22126 18468 22132 18480
rect 17207 18440 17940 18468
rect 22087 18440 22132 18468
rect 17207 18437 17219 18440
rect 17161 18431 17219 18437
rect 22126 18428 22132 18440
rect 22184 18428 22190 18480
rect 23690 18468 23696 18480
rect 23651 18440 23696 18468
rect 23690 18428 23696 18440
rect 23748 18428 23754 18480
rect 23846 18468 23874 18508
rect 24702 18496 24708 18548
rect 24760 18496 24766 18548
rect 25272 18468 25300 18576
rect 27465 18573 27477 18576
rect 27511 18604 27523 18607
rect 27738 18604 27744 18616
rect 27511 18576 27744 18604
rect 27511 18573 27523 18576
rect 27465 18567 27523 18573
rect 27738 18564 27744 18576
rect 27796 18604 27802 18616
rect 28198 18604 28204 18616
rect 27796 18576 28204 18604
rect 27796 18564 27802 18576
rect 28198 18564 28204 18576
rect 28256 18564 28262 18616
rect 28661 18607 28719 18613
rect 28661 18573 28673 18607
rect 28707 18573 28719 18607
rect 28661 18567 28719 18573
rect 26634 18496 26640 18548
rect 26692 18536 26698 18548
rect 27557 18539 27615 18545
rect 27557 18536 27569 18539
rect 26692 18508 27569 18536
rect 26692 18496 26698 18508
rect 27557 18505 27569 18508
rect 27603 18536 27615 18539
rect 28676 18536 28704 18567
rect 27603 18508 28704 18536
rect 27603 18505 27615 18508
rect 27557 18499 27615 18505
rect 28124 18480 28152 18508
rect 28106 18468 28112 18480
rect 23846 18440 25300 18468
rect 28067 18440 28112 18468
rect 28106 18428 28112 18440
rect 28164 18468 28170 18480
rect 28293 18471 28351 18477
rect 28293 18468 28305 18471
rect 28164 18440 28305 18468
rect 28164 18428 28170 18440
rect 28293 18437 28305 18440
rect 28339 18437 28351 18471
rect 28293 18431 28351 18437
rect 29394 18428 29400 18480
rect 29452 18468 29458 18480
rect 29452 18440 29497 18468
rect 29452 18428 29458 18440
rect 400 18378 31680 18400
rect 400 18326 18870 18378
rect 18922 18326 18934 18378
rect 18986 18326 18998 18378
rect 19050 18326 19062 18378
rect 19114 18326 19126 18378
rect 19178 18326 31680 18378
rect 400 18304 31680 18326
rect 4002 18224 4008 18276
rect 4060 18264 4066 18276
rect 6118 18264 6124 18276
rect 4060 18236 6124 18264
rect 4060 18224 4066 18236
rect 6118 18224 6124 18236
rect 6176 18224 6182 18276
rect 4370 18156 4376 18208
rect 4428 18196 4434 18208
rect 6397 18199 6455 18205
rect 6397 18196 6409 18199
rect 4428 18168 6409 18196
rect 4428 18156 4434 18168
rect 6397 18165 6409 18168
rect 6443 18196 6455 18199
rect 6946 18196 6952 18208
rect 6443 18168 6952 18196
rect 6443 18165 6455 18168
rect 6397 18159 6455 18165
rect 6946 18156 6952 18168
rect 7004 18156 7010 18208
rect 14582 18196 14588 18208
rect 14495 18168 14588 18196
rect 14582 18156 14588 18168
rect 14640 18196 14646 18208
rect 16146 18196 16152 18208
rect 14640 18168 16152 18196
rect 14640 18156 14646 18168
rect 16146 18156 16152 18168
rect 16204 18156 16210 18208
rect 21114 18156 21120 18208
rect 21172 18156 21178 18208
rect 26634 18196 26640 18208
rect 26595 18168 26640 18196
rect 26634 18156 26640 18168
rect 26692 18156 26698 18208
rect 28293 18199 28351 18205
rect 28293 18165 28305 18199
rect 28339 18196 28351 18199
rect 28382 18196 28388 18208
rect 28339 18168 28388 18196
rect 28339 18165 28351 18168
rect 28293 18159 28351 18165
rect 28382 18156 28388 18168
rect 28440 18156 28446 18208
rect 28750 18156 28756 18208
rect 28808 18156 28814 18208
rect 4738 18088 4744 18140
rect 4796 18128 4802 18140
rect 4833 18131 4891 18137
rect 4833 18128 4845 18131
rect 4796 18100 4845 18128
rect 4796 18088 4802 18100
rect 4833 18097 4845 18100
rect 4879 18097 4891 18131
rect 4833 18091 4891 18097
rect 4980 18131 5038 18137
rect 4980 18097 4992 18131
rect 5026 18128 5038 18131
rect 6486 18128 6492 18140
rect 5026 18100 6492 18128
rect 5026 18097 5038 18100
rect 4980 18091 5038 18097
rect 6486 18088 6492 18100
rect 6544 18137 6550 18140
rect 6544 18131 6602 18137
rect 6544 18097 6556 18131
rect 6590 18128 6602 18131
rect 7314 18128 7320 18140
rect 6590 18100 7320 18128
rect 6590 18097 6602 18100
rect 6544 18091 6602 18097
rect 6544 18088 6550 18091
rect 7314 18088 7320 18100
rect 7372 18088 7378 18140
rect 12742 18088 12748 18140
rect 12800 18128 12806 18140
rect 12837 18131 12895 18137
rect 12837 18128 12849 18131
rect 12800 18100 12849 18128
rect 12800 18088 12806 18100
rect 12837 18097 12849 18100
rect 12883 18097 12895 18131
rect 12837 18091 12895 18097
rect 12926 18088 12932 18140
rect 12984 18128 12990 18140
rect 13110 18128 13116 18140
rect 12984 18100 13029 18128
rect 13071 18100 13116 18128
rect 12984 18088 12990 18100
rect 13110 18088 13116 18100
rect 13168 18088 13174 18140
rect 14766 18128 14772 18140
rect 14727 18100 14772 18128
rect 14766 18088 14772 18100
rect 14824 18088 14830 18140
rect 15137 18131 15195 18137
rect 15137 18097 15149 18131
rect 15183 18128 15195 18131
rect 15226 18128 15232 18140
rect 15183 18100 15232 18128
rect 15183 18097 15195 18100
rect 15137 18091 15195 18097
rect 15226 18088 15232 18100
rect 15284 18088 15290 18140
rect 16606 18128 16612 18140
rect 16567 18100 16612 18128
rect 16606 18088 16612 18100
rect 16664 18088 16670 18140
rect 17066 18128 17072 18140
rect 17027 18100 17072 18128
rect 17066 18088 17072 18100
rect 17124 18088 17130 18140
rect 17434 18088 17440 18140
rect 17492 18128 17498 18140
rect 18817 18131 18875 18137
rect 18817 18128 18829 18131
rect 17492 18100 18829 18128
rect 17492 18088 17498 18100
rect 18817 18097 18829 18100
rect 18863 18128 18875 18131
rect 19001 18131 19059 18137
rect 19001 18128 19013 18131
rect 18863 18100 19013 18128
rect 18863 18097 18875 18100
rect 18817 18091 18875 18097
rect 19001 18097 19013 18100
rect 19047 18097 19059 18131
rect 19001 18091 19059 18097
rect 26450 18088 26456 18140
rect 26508 18128 26514 18140
rect 26821 18131 26879 18137
rect 26821 18128 26833 18131
rect 26508 18100 26833 18128
rect 26508 18088 26514 18100
rect 26821 18097 26833 18100
rect 26867 18097 26879 18131
rect 28014 18128 28020 18140
rect 27975 18100 28020 18128
rect 26821 18091 26879 18097
rect 28014 18088 28020 18100
rect 28072 18088 28078 18140
rect 5201 18063 5259 18069
rect 5201 18029 5213 18063
rect 5247 18060 5259 18063
rect 5474 18060 5480 18072
rect 5247 18032 5480 18060
rect 5247 18029 5259 18032
rect 5201 18023 5259 18029
rect 5474 18020 5480 18032
rect 5532 18020 5538 18072
rect 6670 18020 6676 18072
rect 6728 18060 6734 18072
rect 6765 18063 6823 18069
rect 6765 18060 6777 18063
rect 6728 18032 6777 18060
rect 6728 18020 6734 18032
rect 6765 18029 6777 18032
rect 6811 18029 6823 18063
rect 13570 18060 13576 18072
rect 13483 18032 13576 18060
rect 6765 18023 6823 18029
rect 13570 18020 13576 18032
rect 13628 18060 13634 18072
rect 16624 18060 16652 18088
rect 17158 18060 17164 18072
rect 13628 18032 16652 18060
rect 17119 18032 17164 18060
rect 13628 18020 13634 18032
rect 17158 18020 17164 18032
rect 17216 18020 17222 18072
rect 17802 18020 17808 18072
rect 17860 18060 17866 18072
rect 20381 18063 20439 18069
rect 20381 18060 20393 18063
rect 17860 18032 20393 18060
rect 17860 18020 17866 18032
rect 20381 18029 20393 18032
rect 20427 18029 20439 18063
rect 20746 18060 20752 18072
rect 20707 18032 20752 18060
rect 20381 18023 20439 18029
rect 20746 18020 20752 18032
rect 20804 18020 20810 18072
rect 21666 18020 21672 18072
rect 21724 18060 21730 18072
rect 22129 18063 22187 18069
rect 22129 18060 22141 18063
rect 21724 18032 22141 18060
rect 21724 18020 21730 18032
rect 22129 18029 22141 18032
rect 22175 18029 22187 18063
rect 30038 18060 30044 18072
rect 29999 18032 30044 18060
rect 22129 18023 22187 18029
rect 30038 18020 30044 18032
rect 30096 18020 30102 18072
rect 5109 17995 5167 18001
rect 5109 17961 5121 17995
rect 5155 17992 5167 17995
rect 5382 17992 5388 18004
rect 5155 17964 5388 17992
rect 5155 17961 5167 17964
rect 5109 17955 5167 17961
rect 5382 17952 5388 17964
rect 5440 17952 5446 18004
rect 6302 17952 6308 18004
rect 6360 17992 6366 18004
rect 6360 17964 6716 17992
rect 6360 17952 6366 17964
rect 5290 17924 5296 17936
rect 5251 17896 5296 17924
rect 5290 17884 5296 17896
rect 5348 17884 5354 17936
rect 6688 17933 6716 17964
rect 6673 17927 6731 17933
rect 6673 17893 6685 17927
rect 6719 17924 6731 17927
rect 6762 17924 6768 17936
rect 6719 17896 6768 17924
rect 6719 17893 6731 17896
rect 6673 17887 6731 17893
rect 6762 17884 6768 17896
rect 6820 17884 6826 17936
rect 7041 17927 7099 17933
rect 7041 17893 7053 17927
rect 7087 17924 7099 17927
rect 7222 17924 7228 17936
rect 7087 17896 7228 17924
rect 7087 17893 7099 17896
rect 7041 17887 7099 17893
rect 7222 17884 7228 17896
rect 7280 17884 7286 17936
rect 17897 17927 17955 17933
rect 17897 17893 17909 17927
rect 17943 17924 17955 17927
rect 18170 17924 18176 17936
rect 17943 17896 18176 17924
rect 17943 17893 17955 17896
rect 17897 17887 17955 17893
rect 18170 17884 18176 17896
rect 18228 17884 18234 17936
rect 18817 17927 18875 17933
rect 18817 17893 18829 17927
rect 18863 17924 18875 17927
rect 19277 17927 19335 17933
rect 19277 17924 19289 17927
rect 18863 17896 19289 17924
rect 18863 17893 18875 17896
rect 18817 17887 18875 17893
rect 19277 17893 19289 17896
rect 19323 17924 19335 17927
rect 19826 17924 19832 17936
rect 19323 17896 19832 17924
rect 19323 17893 19335 17896
rect 19277 17887 19335 17893
rect 19826 17884 19832 17896
rect 19884 17924 19890 17936
rect 20930 17924 20936 17936
rect 19884 17896 20936 17924
rect 19884 17884 19890 17896
rect 20930 17884 20936 17896
rect 20988 17884 20994 17936
rect 23414 17884 23420 17936
rect 23472 17924 23478 17936
rect 23782 17924 23788 17936
rect 23472 17896 23788 17924
rect 23472 17884 23478 17896
rect 23782 17884 23788 17896
rect 23840 17924 23846 17936
rect 23966 17924 23972 17936
rect 23840 17896 23972 17924
rect 23840 17884 23846 17896
rect 23966 17884 23972 17896
rect 24024 17884 24030 17936
rect 24061 17927 24119 17933
rect 24061 17893 24073 17927
rect 24107 17924 24119 17927
rect 24242 17924 24248 17936
rect 24107 17896 24248 17924
rect 24107 17893 24119 17896
rect 24061 17887 24119 17893
rect 24242 17884 24248 17896
rect 24300 17884 24306 17936
rect 26910 17924 26916 17936
rect 26871 17896 26916 17924
rect 26910 17884 26916 17896
rect 26968 17884 26974 17936
rect 400 17834 31680 17856
rect 400 17782 3510 17834
rect 3562 17782 3574 17834
rect 3626 17782 3638 17834
rect 3690 17782 3702 17834
rect 3754 17782 3766 17834
rect 3818 17782 31680 17834
rect 400 17760 31680 17782
rect 3545 17723 3603 17729
rect 3545 17689 3557 17723
rect 3591 17720 3603 17723
rect 4281 17723 4339 17729
rect 4281 17720 4293 17723
rect 3591 17692 4293 17720
rect 3591 17689 3603 17692
rect 3545 17683 3603 17689
rect 4281 17689 4293 17692
rect 4327 17720 4339 17723
rect 5290 17720 5296 17732
rect 4327 17692 5296 17720
rect 4327 17689 4339 17692
rect 4281 17683 4339 17689
rect 1797 17519 1855 17525
rect 1797 17485 1809 17519
rect 1843 17516 1855 17519
rect 2346 17516 2352 17528
rect 1843 17488 2352 17516
rect 1843 17485 1855 17488
rect 1797 17479 1855 17485
rect 2346 17476 2352 17488
rect 2404 17476 2410 17528
rect 3269 17519 3327 17525
rect 3269 17485 3281 17519
rect 3315 17516 3327 17519
rect 3560 17516 3588 17683
rect 5290 17680 5296 17692
rect 5348 17680 5354 17732
rect 5569 17723 5627 17729
rect 5569 17689 5581 17723
rect 5615 17720 5627 17723
rect 6486 17720 6492 17732
rect 5615 17692 6492 17720
rect 5615 17689 5627 17692
rect 5569 17683 5627 17689
rect 6486 17680 6492 17692
rect 6544 17680 6550 17732
rect 6670 17720 6676 17732
rect 6631 17692 6676 17720
rect 6670 17680 6676 17692
rect 6728 17680 6734 17732
rect 6762 17680 6768 17732
rect 6820 17720 6826 17732
rect 6946 17720 6952 17732
rect 6820 17692 6865 17720
rect 6907 17692 6952 17720
rect 6820 17680 6826 17692
rect 6946 17680 6952 17692
rect 7004 17680 7010 17732
rect 9065 17723 9123 17729
rect 9065 17689 9077 17723
rect 9111 17720 9123 17723
rect 11546 17720 11552 17732
rect 9111 17692 11552 17720
rect 9111 17689 9123 17692
rect 9065 17683 9123 17689
rect 4649 17655 4707 17661
rect 4649 17621 4661 17655
rect 4695 17652 4707 17655
rect 4738 17652 4744 17664
rect 4695 17624 4744 17652
rect 4695 17621 4707 17624
rect 4649 17615 4707 17621
rect 4738 17612 4744 17624
rect 4796 17612 4802 17664
rect 5385 17587 5443 17593
rect 3315 17488 3588 17516
rect 4388 17556 4876 17584
rect 3315 17485 3327 17488
rect 3269 17479 3327 17485
rect 1610 17448 1616 17460
rect 1523 17420 1616 17448
rect 1610 17408 1616 17420
rect 1668 17448 1674 17460
rect 2533 17451 2591 17457
rect 2533 17448 2545 17451
rect 1668 17420 2545 17448
rect 1668 17408 1674 17420
rect 2533 17417 2545 17420
rect 2579 17448 2591 17451
rect 3361 17451 3419 17457
rect 3361 17448 3373 17451
rect 2579 17420 3373 17448
rect 2579 17417 2591 17420
rect 2533 17411 2591 17417
rect 3361 17417 3373 17420
rect 3407 17448 3419 17451
rect 3637 17451 3695 17457
rect 3637 17448 3649 17451
rect 3407 17420 3649 17448
rect 3407 17417 3419 17420
rect 3361 17411 3419 17417
rect 3637 17417 3649 17420
rect 3683 17417 3695 17451
rect 3637 17411 3695 17417
rect 1242 17340 1248 17392
rect 1300 17380 1306 17392
rect 1521 17383 1579 17389
rect 1521 17380 1533 17383
rect 1300 17352 1533 17380
rect 1300 17340 1306 17352
rect 1521 17349 1533 17352
rect 1567 17380 1579 17383
rect 1794 17380 1800 17392
rect 1567 17352 1800 17380
rect 1567 17349 1579 17352
rect 1521 17343 1579 17349
rect 1794 17340 1800 17352
rect 1852 17380 1858 17392
rect 1889 17383 1947 17389
rect 1889 17380 1901 17383
rect 1852 17352 1901 17380
rect 1852 17340 1858 17352
rect 1889 17349 1901 17352
rect 1935 17349 1947 17383
rect 2346 17380 2352 17392
rect 2307 17352 2352 17380
rect 1889 17343 1947 17349
rect 2346 17340 2352 17352
rect 2404 17340 2410 17392
rect 3910 17340 3916 17392
rect 3968 17380 3974 17392
rect 4388 17389 4416 17556
rect 4741 17519 4799 17525
rect 4741 17485 4753 17519
rect 4787 17485 4799 17519
rect 4741 17479 4799 17485
rect 4462 17408 4468 17460
rect 4520 17448 4526 17460
rect 4554 17448 4560 17460
rect 4520 17420 4560 17448
rect 4520 17408 4526 17420
rect 4554 17408 4560 17420
rect 4612 17408 4618 17460
rect 4373 17383 4431 17389
rect 4373 17380 4385 17383
rect 3968 17352 4385 17380
rect 3968 17340 3974 17352
rect 4373 17349 4385 17352
rect 4419 17349 4431 17383
rect 4756 17380 4784 17479
rect 4848 17460 4876 17556
rect 5385 17553 5397 17587
rect 5431 17584 5443 17587
rect 8329 17587 8387 17593
rect 8329 17584 8341 17587
rect 5431 17556 8341 17584
rect 5431 17553 5443 17556
rect 5385 17547 5443 17553
rect 8329 17553 8341 17556
rect 8375 17584 8387 17587
rect 9080 17584 9108 17683
rect 11546 17680 11552 17692
rect 11604 17680 11610 17732
rect 12742 17720 12748 17732
rect 12703 17692 12748 17720
rect 12742 17680 12748 17692
rect 12800 17680 12806 17732
rect 12837 17723 12895 17729
rect 12837 17689 12849 17723
rect 12883 17720 12895 17723
rect 13018 17720 13024 17732
rect 12883 17692 13024 17720
rect 12883 17689 12895 17692
rect 12837 17683 12895 17689
rect 13018 17680 13024 17692
rect 13076 17720 13082 17732
rect 13076 17692 13616 17720
rect 13076 17680 13082 17692
rect 9249 17655 9307 17661
rect 9249 17621 9261 17655
rect 9295 17652 9307 17655
rect 11914 17652 11920 17664
rect 9295 17624 11920 17652
rect 9295 17621 9307 17624
rect 9249 17615 9307 17621
rect 8375 17556 9108 17584
rect 8375 17553 8387 17556
rect 8329 17547 8387 17553
rect 4830 17408 4836 17460
rect 4888 17448 4894 17460
rect 5017 17451 5075 17457
rect 5017 17448 5029 17451
rect 4888 17420 5029 17448
rect 4888 17408 4894 17420
rect 5017 17417 5029 17420
rect 5063 17417 5075 17451
rect 5017 17411 5075 17417
rect 5198 17380 5204 17392
rect 4756 17352 5204 17380
rect 4373 17343 4431 17349
rect 5198 17340 5204 17352
rect 5256 17380 5262 17392
rect 5400 17380 5428 17547
rect 5474 17476 5480 17528
rect 5532 17516 5538 17528
rect 5661 17519 5719 17525
rect 5661 17516 5673 17519
rect 5532 17488 5673 17516
rect 5532 17476 5538 17488
rect 5661 17485 5673 17488
rect 5707 17485 5719 17519
rect 8418 17516 8424 17528
rect 8331 17488 8424 17516
rect 5661 17479 5719 17485
rect 8418 17476 8424 17488
rect 8476 17516 8482 17528
rect 9264 17516 9292 17615
rect 11914 17612 11920 17624
rect 11972 17612 11978 17664
rect 12561 17655 12619 17661
rect 12561 17621 12573 17655
rect 12607 17652 12619 17655
rect 12926 17652 12932 17664
rect 12607 17624 12932 17652
rect 12607 17621 12619 17624
rect 12561 17615 12619 17621
rect 12926 17612 12932 17624
rect 12984 17652 12990 17664
rect 13113 17655 13171 17661
rect 13113 17652 13125 17655
rect 12984 17624 13125 17652
rect 12984 17612 12990 17624
rect 13113 17621 13125 17624
rect 13159 17621 13171 17655
rect 13113 17615 13171 17621
rect 13588 17584 13616 17692
rect 13662 17680 13668 17732
rect 13720 17720 13726 17732
rect 13849 17723 13907 17729
rect 13849 17720 13861 17723
rect 13720 17692 13861 17720
rect 13720 17680 13726 17692
rect 13849 17689 13861 17692
rect 13895 17720 13907 17723
rect 14766 17720 14772 17732
rect 13895 17692 14772 17720
rect 13895 17689 13907 17692
rect 13849 17683 13907 17689
rect 14766 17680 14772 17692
rect 14824 17720 14830 17732
rect 15413 17723 15471 17729
rect 15413 17720 15425 17723
rect 14824 17692 15425 17720
rect 14824 17680 14830 17692
rect 15413 17689 15425 17692
rect 15459 17689 15471 17723
rect 15413 17683 15471 17689
rect 17069 17723 17127 17729
rect 17069 17689 17081 17723
rect 17115 17720 17127 17723
rect 17158 17720 17164 17732
rect 17115 17692 17164 17720
rect 17115 17689 17127 17692
rect 17069 17683 17127 17689
rect 17158 17680 17164 17692
rect 17216 17720 17222 17732
rect 20194 17720 20200 17732
rect 17216 17692 20200 17720
rect 17216 17680 17222 17692
rect 20194 17680 20200 17692
rect 20252 17680 20258 17732
rect 20289 17723 20347 17729
rect 20289 17689 20301 17723
rect 20335 17720 20347 17723
rect 20746 17720 20752 17732
rect 20335 17692 20752 17720
rect 20335 17689 20347 17692
rect 20289 17683 20347 17689
rect 20746 17680 20752 17692
rect 20804 17680 20810 17732
rect 20838 17680 20844 17732
rect 20896 17720 20902 17732
rect 21577 17723 21635 17729
rect 21577 17720 21589 17723
rect 20896 17692 21589 17720
rect 20896 17680 20902 17692
rect 21577 17689 21589 17692
rect 21623 17720 21635 17723
rect 22126 17720 22132 17732
rect 21623 17692 22132 17720
rect 21623 17689 21635 17692
rect 21577 17683 21635 17689
rect 22126 17680 22132 17692
rect 22184 17720 22190 17732
rect 23874 17720 23880 17732
rect 22184 17692 23880 17720
rect 22184 17680 22190 17692
rect 23874 17680 23880 17692
rect 23932 17680 23938 17732
rect 26361 17723 26419 17729
rect 26361 17689 26373 17723
rect 26407 17720 26419 17723
rect 26910 17720 26916 17732
rect 26407 17692 26916 17720
rect 26407 17689 26419 17692
rect 26361 17683 26419 17689
rect 26910 17680 26916 17692
rect 26968 17680 26974 17732
rect 28109 17723 28167 17729
rect 28109 17689 28121 17723
rect 28155 17720 28167 17723
rect 30038 17720 30044 17732
rect 28155 17692 30044 17720
rect 28155 17689 28167 17692
rect 28109 17683 28167 17689
rect 30038 17680 30044 17692
rect 30096 17680 30102 17732
rect 14309 17655 14367 17661
rect 14309 17621 14321 17655
rect 14355 17652 14367 17655
rect 14493 17655 14551 17661
rect 14493 17652 14505 17655
rect 14355 17624 14505 17652
rect 14355 17621 14367 17624
rect 14309 17615 14367 17621
rect 14493 17621 14505 17624
rect 14539 17652 14551 17655
rect 14582 17652 14588 17664
rect 14539 17624 14588 17652
rect 14539 17621 14551 17624
rect 14493 17615 14551 17621
rect 14582 17612 14588 17624
rect 14640 17612 14646 17664
rect 19918 17652 19924 17664
rect 19879 17624 19924 17652
rect 19918 17612 19924 17624
rect 19976 17612 19982 17664
rect 20657 17655 20715 17661
rect 20657 17621 20669 17655
rect 20703 17652 20715 17655
rect 21666 17652 21672 17664
rect 20703 17624 21672 17652
rect 20703 17621 20715 17624
rect 20657 17615 20715 17621
rect 21666 17612 21672 17624
rect 21724 17612 21730 17664
rect 26450 17612 26456 17664
rect 26508 17652 26514 17664
rect 26729 17655 26787 17661
rect 26729 17652 26741 17655
rect 26508 17624 26741 17652
rect 26508 17612 26514 17624
rect 26729 17621 26741 17624
rect 26775 17621 26787 17655
rect 26729 17615 26787 17621
rect 28014 17612 28020 17664
rect 28072 17652 28078 17664
rect 28753 17655 28811 17661
rect 28753 17652 28765 17655
rect 28072 17624 28765 17652
rect 28072 17612 28078 17624
rect 28753 17621 28765 17624
rect 28799 17621 28811 17655
rect 28753 17615 28811 17621
rect 18170 17584 18176 17596
rect 13588 17556 14214 17584
rect 18131 17556 18176 17584
rect 8476 17488 9292 17516
rect 8476 17476 8482 17488
rect 12742 17476 12748 17528
rect 12800 17516 12806 17528
rect 13021 17519 13079 17525
rect 13021 17516 13033 17519
rect 12800 17488 13033 17516
rect 12800 17476 12806 17488
rect 13021 17485 13033 17488
rect 13067 17485 13079 17519
rect 13021 17479 13079 17485
rect 13297 17519 13355 17525
rect 13297 17485 13309 17519
rect 13343 17516 13355 17519
rect 13662 17516 13668 17528
rect 13343 17488 13668 17516
rect 13343 17485 13355 17488
rect 13297 17479 13355 17485
rect 13662 17476 13668 17488
rect 13720 17476 13726 17528
rect 14186 17516 14214 17556
rect 18170 17544 18176 17556
rect 18228 17544 18234 17596
rect 23966 17584 23972 17596
rect 23927 17556 23972 17584
rect 23966 17544 23972 17556
rect 24024 17544 24030 17596
rect 24242 17544 24248 17596
rect 24300 17584 24306 17596
rect 24337 17587 24395 17593
rect 24337 17584 24349 17587
rect 24300 17556 24349 17584
rect 24300 17544 24306 17556
rect 24337 17553 24349 17556
rect 24383 17553 24395 17587
rect 24337 17547 24395 17553
rect 25530 17544 25536 17596
rect 25588 17584 25594 17596
rect 25717 17587 25775 17593
rect 25717 17584 25729 17587
rect 25588 17556 25729 17584
rect 25588 17544 25594 17556
rect 25717 17553 25729 17556
rect 25763 17553 25775 17587
rect 25717 17547 25775 17553
rect 26545 17587 26603 17593
rect 26545 17553 26557 17587
rect 26591 17584 26603 17587
rect 26634 17584 26640 17596
rect 26591 17556 26640 17584
rect 26591 17553 26603 17556
rect 26545 17547 26603 17553
rect 26634 17544 26640 17556
rect 26692 17544 26698 17596
rect 28293 17587 28351 17593
rect 28293 17553 28305 17587
rect 28339 17584 28351 17587
rect 28382 17584 28388 17596
rect 28339 17556 28388 17584
rect 28339 17553 28351 17556
rect 28293 17547 28351 17553
rect 28382 17544 28388 17556
rect 28440 17544 28446 17596
rect 14769 17519 14827 17525
rect 14769 17516 14781 17519
rect 14186 17488 14781 17516
rect 14769 17485 14781 17488
rect 14815 17516 14827 17519
rect 15229 17519 15287 17525
rect 15229 17516 15241 17519
rect 14815 17488 15241 17516
rect 14815 17485 14827 17488
rect 14769 17479 14827 17485
rect 15229 17485 15241 17488
rect 15275 17485 15287 17519
rect 17802 17516 17808 17528
rect 17763 17488 17808 17516
rect 15229 17479 15287 17485
rect 17802 17476 17808 17488
rect 17860 17476 17866 17528
rect 20838 17516 20844 17528
rect 20799 17488 20844 17516
rect 20838 17476 20844 17488
rect 20896 17476 20902 17528
rect 20930 17476 20936 17528
rect 20988 17516 20994 17528
rect 21669 17519 21727 17525
rect 21669 17516 21681 17519
rect 20988 17488 21681 17516
rect 20988 17476 20994 17488
rect 21669 17485 21681 17488
rect 21715 17516 21727 17519
rect 22494 17516 22500 17528
rect 21715 17488 22500 17516
rect 21715 17485 21727 17488
rect 21669 17479 21727 17485
rect 22494 17476 22500 17488
rect 22552 17476 22558 17528
rect 25898 17476 25904 17528
rect 25956 17516 25962 17528
rect 27097 17519 27155 17525
rect 27097 17516 27109 17519
rect 25956 17488 27109 17516
rect 25956 17476 25962 17488
rect 27097 17485 27109 17488
rect 27143 17516 27155 17519
rect 27557 17519 27615 17525
rect 27557 17516 27569 17519
rect 27143 17488 27569 17516
rect 27143 17485 27155 17488
rect 27097 17479 27155 17485
rect 27557 17485 27569 17488
rect 27603 17485 27615 17519
rect 27557 17479 27615 17485
rect 8237 17451 8295 17457
rect 8237 17417 8249 17451
rect 8283 17448 8295 17451
rect 8881 17451 8939 17457
rect 8881 17448 8893 17451
rect 8283 17420 8893 17448
rect 8283 17417 8295 17420
rect 8237 17411 8295 17417
rect 8881 17417 8893 17420
rect 8927 17448 8939 17451
rect 9062 17448 9068 17460
rect 8927 17420 9068 17448
rect 8927 17417 8939 17420
rect 8881 17411 8939 17417
rect 9062 17408 9068 17420
rect 9120 17408 9126 17460
rect 12377 17451 12435 17457
rect 12377 17417 12389 17451
rect 12423 17448 12435 17451
rect 13754 17448 13760 17460
rect 12423 17420 13760 17448
rect 12423 17417 12435 17420
rect 12377 17411 12435 17417
rect 13754 17408 13760 17420
rect 13812 17408 13818 17460
rect 14582 17448 14588 17460
rect 14543 17420 14588 17448
rect 14582 17408 14588 17420
rect 14640 17408 14646 17460
rect 16422 17408 16428 17460
rect 16480 17448 16486 17460
rect 16793 17451 16851 17457
rect 16793 17448 16805 17451
rect 16480 17420 16805 17448
rect 16480 17408 16486 17420
rect 16793 17417 16805 17420
rect 16839 17448 16851 17451
rect 17066 17448 17072 17460
rect 16839 17420 17072 17448
rect 16839 17417 16851 17420
rect 16793 17411 16851 17417
rect 17066 17408 17072 17420
rect 17124 17408 17130 17460
rect 20102 17448 20108 17460
rect 7222 17380 7228 17392
rect 5256 17352 5428 17380
rect 7183 17352 7228 17380
rect 5256 17340 5262 17352
rect 7222 17340 7228 17352
rect 7280 17340 7286 17392
rect 14122 17380 14128 17392
rect 14083 17352 14128 17380
rect 14122 17340 14128 17352
rect 14180 17340 14186 17392
rect 14306 17340 14312 17392
rect 14364 17380 14370 17392
rect 14861 17383 14919 17389
rect 14861 17380 14873 17383
rect 14364 17352 14873 17380
rect 14364 17340 14370 17352
rect 14861 17349 14873 17352
rect 14907 17380 14919 17383
rect 15597 17383 15655 17389
rect 15597 17380 15609 17383
rect 14907 17352 15609 17380
rect 14907 17349 14919 17352
rect 14861 17343 14919 17349
rect 15597 17349 15609 17352
rect 15643 17380 15655 17383
rect 15962 17380 15968 17392
rect 15643 17352 15968 17380
rect 15643 17349 15655 17352
rect 15597 17343 15655 17349
rect 15962 17340 15968 17352
rect 16020 17340 16026 17392
rect 16054 17340 16060 17392
rect 16112 17380 16118 17392
rect 16606 17380 16612 17392
rect 16112 17352 16612 17380
rect 16112 17340 16118 17352
rect 16606 17340 16612 17352
rect 16664 17340 16670 17392
rect 17526 17380 17532 17392
rect 17487 17352 17532 17380
rect 17526 17340 17532 17352
rect 17584 17340 17590 17392
rect 17713 17383 17771 17389
rect 17713 17349 17725 17383
rect 17759 17380 17771 17383
rect 19200 17380 19228 17448
rect 20015 17420 20108 17448
rect 20102 17408 20108 17420
rect 20160 17448 20166 17460
rect 21390 17448 21396 17460
rect 20160 17420 21396 17448
rect 20160 17408 20166 17420
rect 21390 17408 21396 17420
rect 21448 17408 21454 17460
rect 22586 17408 22592 17460
rect 22644 17448 22650 17460
rect 23690 17448 23696 17460
rect 22644 17420 23696 17448
rect 22644 17408 22650 17420
rect 23690 17408 23696 17420
rect 23748 17448 23754 17460
rect 23785 17451 23843 17457
rect 23785 17448 23797 17451
rect 23748 17420 23797 17448
rect 23748 17408 23754 17420
rect 23785 17417 23797 17420
rect 23831 17417 23843 17451
rect 23785 17411 23843 17417
rect 20194 17380 20200 17392
rect 17759 17352 20200 17380
rect 17759 17349 17771 17352
rect 17713 17343 17771 17349
rect 20194 17340 20200 17352
rect 20252 17380 20258 17392
rect 20381 17383 20439 17389
rect 20381 17380 20393 17383
rect 20252 17352 20393 17380
rect 20252 17340 20258 17352
rect 20381 17349 20393 17352
rect 20427 17380 20439 17383
rect 21114 17380 21120 17392
rect 20427 17352 21120 17380
rect 20427 17349 20439 17352
rect 20381 17343 20439 17349
rect 21114 17340 21120 17352
rect 21172 17340 21178 17392
rect 21850 17380 21856 17392
rect 21811 17352 21856 17380
rect 21850 17340 21856 17352
rect 21908 17380 21914 17392
rect 23414 17380 23420 17392
rect 21908 17352 23420 17380
rect 21908 17340 21914 17352
rect 23414 17340 23420 17352
rect 23472 17340 23478 17392
rect 23598 17380 23604 17392
rect 23559 17352 23604 17380
rect 23598 17340 23604 17352
rect 23656 17340 23662 17392
rect 23800 17380 23828 17411
rect 24702 17408 24708 17460
rect 24760 17408 24766 17460
rect 26913 17451 26971 17457
rect 26913 17417 26925 17451
rect 26959 17448 26971 17451
rect 27833 17451 27891 17457
rect 27833 17448 27845 17451
rect 26959 17420 27845 17448
rect 26959 17417 26971 17420
rect 26913 17411 26971 17417
rect 27833 17417 27845 17420
rect 27879 17448 27891 17451
rect 28474 17448 28480 17460
rect 27879 17420 28480 17448
rect 27879 17417 27891 17420
rect 27833 17411 27891 17417
rect 28474 17408 28480 17420
rect 28532 17408 28538 17460
rect 24720 17380 24748 17408
rect 27186 17380 27192 17392
rect 23800 17352 24748 17380
rect 27147 17352 27192 17380
rect 27186 17340 27192 17352
rect 27244 17340 27250 17392
rect 28566 17380 28572 17392
rect 28527 17352 28572 17380
rect 28566 17340 28572 17352
rect 28624 17340 28630 17392
rect 400 17290 31680 17312
rect 400 17238 18870 17290
rect 18922 17238 18934 17290
rect 18986 17238 18998 17290
rect 19050 17238 19062 17290
rect 19114 17238 19126 17290
rect 19178 17238 31680 17290
rect 400 17216 31680 17238
rect 1242 17176 1248 17188
rect 1203 17148 1248 17176
rect 1242 17136 1248 17148
rect 1300 17136 1306 17188
rect 4738 17136 4744 17188
rect 4796 17176 4802 17188
rect 12929 17179 12987 17185
rect 4796 17148 6348 17176
rect 4796 17136 4802 17148
rect 4925 17111 4983 17117
rect 4925 17077 4937 17111
rect 4971 17108 4983 17111
rect 4971 17080 5336 17108
rect 4971 17077 4983 17080
rect 4925 17071 4983 17077
rect 1610 17040 1616 17052
rect 1571 17012 1616 17040
rect 1610 17000 1616 17012
rect 1668 17000 1674 17052
rect 2073 17043 2131 17049
rect 2073 17009 2085 17043
rect 2119 17040 2131 17043
rect 2346 17040 2352 17052
rect 2119 17012 2352 17040
rect 2119 17009 2131 17012
rect 2073 17003 2131 17009
rect 2346 17000 2352 17012
rect 2404 17040 2410 17052
rect 4189 17043 4247 17049
rect 2404 17012 4140 17040
rect 2404 17000 2410 17012
rect 4112 16984 4140 17012
rect 4189 17009 4201 17043
rect 4235 17040 4247 17043
rect 4278 17040 4284 17052
rect 4235 17012 4284 17040
rect 4235 17009 4247 17012
rect 4189 17003 4247 17009
rect 4278 17000 4284 17012
rect 4336 17040 4342 17052
rect 4462 17040 4468 17052
rect 4336 17012 4468 17040
rect 4336 17000 4342 17012
rect 4462 17000 4468 17012
rect 4520 17000 4526 17052
rect 5198 17040 5204 17052
rect 5159 17012 5204 17040
rect 5198 17000 5204 17012
rect 5256 17000 5262 17052
rect 5308 17049 5336 17080
rect 5293 17043 5351 17049
rect 5293 17009 5305 17043
rect 5339 17040 5351 17043
rect 5382 17040 5388 17052
rect 5339 17012 5388 17040
rect 5339 17009 5351 17012
rect 5293 17003 5351 17009
rect 5382 17000 5388 17012
rect 5440 17000 5446 17052
rect 5474 17000 5480 17052
rect 5532 17040 5538 17052
rect 6320 17040 6348 17148
rect 12929 17145 12941 17179
rect 12975 17176 12987 17179
rect 13570 17176 13576 17188
rect 12975 17148 13576 17176
rect 12975 17145 12987 17148
rect 12929 17139 12987 17145
rect 13570 17136 13576 17148
rect 13628 17136 13634 17188
rect 14122 17136 14128 17188
rect 14180 17176 14186 17188
rect 15226 17176 15232 17188
rect 14180 17148 15232 17176
rect 14180 17136 14186 17148
rect 15226 17136 15232 17148
rect 15284 17136 15290 17188
rect 18170 17176 18176 17188
rect 18131 17148 18176 17176
rect 18170 17136 18176 17148
rect 18228 17136 18234 17188
rect 20473 17179 20531 17185
rect 20473 17145 20485 17179
rect 20519 17176 20531 17179
rect 20746 17176 20752 17188
rect 20519 17148 20752 17176
rect 20519 17145 20531 17148
rect 20473 17139 20531 17145
rect 20746 17136 20752 17148
rect 20804 17136 20810 17188
rect 27005 17179 27063 17185
rect 27005 17145 27017 17179
rect 27051 17176 27063 17179
rect 27186 17176 27192 17188
rect 27051 17148 27192 17176
rect 27051 17145 27063 17148
rect 27005 17139 27063 17145
rect 27186 17136 27192 17148
rect 27244 17176 27250 17188
rect 27244 17148 27876 17176
rect 27244 17136 27250 17148
rect 27848 17120 27876 17148
rect 12742 17068 12748 17120
rect 12800 17108 12806 17120
rect 13021 17111 13079 17117
rect 13021 17108 13033 17111
rect 12800 17080 13033 17108
rect 12800 17068 12806 17080
rect 13021 17077 13033 17080
rect 13067 17077 13079 17111
rect 13021 17071 13079 17077
rect 14677 17111 14735 17117
rect 14677 17077 14689 17111
rect 14723 17108 14735 17111
rect 14950 17108 14956 17120
rect 14723 17080 14956 17108
rect 14723 17077 14735 17080
rect 14677 17071 14735 17077
rect 14950 17068 14956 17080
rect 15008 17068 15014 17120
rect 19550 17108 19556 17120
rect 18740 17080 19556 17108
rect 6857 17043 6915 17049
rect 6857 17040 6869 17043
rect 5532 17012 5577 17040
rect 6320 17012 6869 17040
rect 5532 17000 5538 17012
rect 6857 17009 6869 17012
rect 6903 17040 6915 17043
rect 7406 17040 7412 17052
rect 6903 17012 7412 17040
rect 6903 17009 6915 17012
rect 6857 17003 6915 17009
rect 7406 17000 7412 17012
rect 7464 17000 7470 17052
rect 9062 17040 9068 17052
rect 9023 17012 9068 17040
rect 9062 17000 9068 17012
rect 9120 17000 9126 17052
rect 9154 17000 9160 17052
rect 9212 17040 9218 17052
rect 9709 17043 9767 17049
rect 9709 17040 9721 17043
rect 9212 17012 9721 17040
rect 9212 17000 9218 17012
rect 9709 17009 9721 17012
rect 9755 17040 9767 17043
rect 11270 17040 11276 17052
rect 9755 17012 11276 17040
rect 9755 17009 9767 17012
rect 9709 17003 9767 17009
rect 11270 17000 11276 17012
rect 11328 17000 11334 17052
rect 12926 17000 12932 17052
rect 12984 17040 12990 17052
rect 13205 17043 13263 17049
rect 13205 17040 13217 17043
rect 12984 17012 13217 17040
rect 12984 17000 12990 17012
rect 13205 17009 13217 17012
rect 13251 17009 13263 17043
rect 15962 17040 15968 17052
rect 15923 17012 15968 17040
rect 13205 17003 13263 17009
rect 15962 17000 15968 17012
rect 16020 17000 16026 17052
rect 16422 17040 16428 17052
rect 16383 17012 16428 17040
rect 16422 17000 16428 17012
rect 16480 17000 16486 17052
rect 17710 17000 17716 17052
rect 17768 17040 17774 17052
rect 18740 17049 18768 17080
rect 19550 17068 19556 17080
rect 19608 17108 19614 17120
rect 27830 17108 27836 17120
rect 19608 17080 20884 17108
rect 27743 17080 27836 17108
rect 19608 17068 19614 17080
rect 18725 17043 18783 17049
rect 18725 17040 18737 17043
rect 17768 17012 18737 17040
rect 17768 17000 17774 17012
rect 18725 17009 18737 17012
rect 18771 17009 18783 17043
rect 18725 17003 18783 17009
rect 18814 17000 18820 17052
rect 18872 17040 18878 17052
rect 19093 17043 19151 17049
rect 19093 17040 19105 17043
rect 18872 17012 19105 17040
rect 18872 17000 18878 17012
rect 19093 17009 19105 17012
rect 19139 17040 19151 17043
rect 20102 17040 20108 17052
rect 19139 17012 20108 17040
rect 19139 17009 19151 17012
rect 19093 17003 19151 17009
rect 20102 17000 20108 17012
rect 20160 17000 20166 17052
rect 20856 17049 20884 17080
rect 27830 17068 27836 17080
rect 27888 17068 27894 17120
rect 20841 17043 20899 17049
rect 20841 17009 20853 17043
rect 20887 17040 20899 17043
rect 20930 17040 20936 17052
rect 20887 17012 20936 17040
rect 20887 17009 20899 17012
rect 20841 17003 20899 17009
rect 20930 17000 20936 17012
rect 20988 17000 20994 17052
rect 21209 17043 21267 17049
rect 21209 17009 21221 17043
rect 21255 17040 21267 17043
rect 21390 17040 21396 17052
rect 21255 17012 21396 17040
rect 21255 17009 21267 17012
rect 21209 17003 21267 17009
rect 21390 17000 21396 17012
rect 21448 17000 21454 17052
rect 22954 17040 22960 17052
rect 22915 17012 22960 17040
rect 22954 17000 22960 17012
rect 23012 17000 23018 17052
rect 23322 17040 23328 17052
rect 23283 17012 23328 17040
rect 23322 17000 23328 17012
rect 23380 17000 23386 17052
rect 27738 17040 27744 17052
rect 27699 17012 27744 17040
rect 27738 17000 27744 17012
rect 27796 17000 27802 17052
rect 27925 17043 27983 17049
rect 27925 17009 27937 17043
rect 27971 17040 27983 17043
rect 28014 17040 28020 17052
rect 27971 17012 28020 17040
rect 27971 17009 27983 17012
rect 27925 17003 27983 17009
rect 28014 17000 28020 17012
rect 28072 17000 28078 17052
rect 1702 16972 1708 16984
rect 1663 16944 1708 16972
rect 1702 16932 1708 16944
rect 1760 16932 1766 16984
rect 3361 16975 3419 16981
rect 3361 16972 3373 16975
rect 2548 16944 3373 16972
rect 2548 16848 2576 16944
rect 3361 16941 3373 16944
rect 3407 16941 3419 16975
rect 3910 16972 3916 16984
rect 3871 16944 3916 16972
rect 3361 16935 3419 16941
rect 3376 16904 3404 16935
rect 3910 16932 3916 16944
rect 3968 16932 3974 16984
rect 4094 16932 4100 16984
rect 4152 16972 4158 16984
rect 4370 16972 4376 16984
rect 4152 16944 4376 16972
rect 4152 16932 4158 16944
rect 4370 16932 4376 16944
rect 4428 16932 4434 16984
rect 5750 16972 5756 16984
rect 5711 16944 5756 16972
rect 5750 16932 5756 16944
rect 5808 16932 5814 16984
rect 6762 16972 6768 16984
rect 6723 16944 6768 16972
rect 6762 16932 6768 16944
rect 6820 16932 6826 16984
rect 7130 16932 7136 16984
rect 7188 16972 7194 16984
rect 7317 16975 7375 16981
rect 7317 16972 7329 16975
rect 7188 16944 7329 16972
rect 7188 16932 7194 16944
rect 7317 16941 7329 16944
rect 7363 16972 7375 16975
rect 7590 16972 7596 16984
rect 7363 16944 7596 16972
rect 7363 16941 7375 16944
rect 7317 16935 7375 16941
rect 7590 16932 7596 16944
rect 7648 16932 7654 16984
rect 9798 16972 9804 16984
rect 9759 16944 9804 16972
rect 9798 16932 9804 16944
rect 9856 16932 9862 16984
rect 16514 16972 16520 16984
rect 16475 16944 16520 16972
rect 16514 16932 16520 16944
rect 16572 16932 16578 16984
rect 18538 16972 18544 16984
rect 18499 16944 18544 16972
rect 18538 16932 18544 16944
rect 18596 16932 18602 16984
rect 18998 16972 19004 16984
rect 18911 16944 19004 16972
rect 18998 16932 19004 16944
rect 19056 16972 19062 16984
rect 19918 16972 19924 16984
rect 19056 16944 19924 16972
rect 19056 16932 19062 16944
rect 19918 16932 19924 16944
rect 19976 16932 19982 16984
rect 20470 16932 20476 16984
rect 20528 16972 20534 16984
rect 20657 16975 20715 16981
rect 20657 16972 20669 16975
rect 20528 16944 20669 16972
rect 20528 16932 20534 16944
rect 20657 16941 20669 16944
rect 20703 16941 20715 16975
rect 20657 16935 20715 16941
rect 21117 16975 21175 16981
rect 21117 16941 21129 16975
rect 21163 16972 21175 16975
rect 21666 16972 21672 16984
rect 21163 16944 21672 16972
rect 21163 16941 21175 16944
rect 21117 16935 21175 16941
rect 4462 16904 4468 16916
rect 3376 16876 4468 16904
rect 4462 16864 4468 16876
rect 4520 16864 4526 16916
rect 9249 16907 9307 16913
rect 9249 16873 9261 16907
rect 9295 16904 9307 16907
rect 9522 16904 9528 16916
rect 9295 16876 9528 16904
rect 9295 16873 9307 16876
rect 9249 16867 9307 16873
rect 9522 16864 9528 16876
rect 9580 16864 9586 16916
rect 17802 16904 17808 16916
rect 14784 16876 17808 16904
rect 14784 16848 14812 16876
rect 17802 16864 17808 16876
rect 17860 16864 17866 16916
rect 20286 16864 20292 16916
rect 20344 16904 20350 16916
rect 21132 16904 21160 16935
rect 21666 16932 21672 16944
rect 21724 16932 21730 16984
rect 22494 16932 22500 16984
rect 22552 16972 22558 16984
rect 22865 16975 22923 16981
rect 22865 16972 22877 16975
rect 22552 16944 22877 16972
rect 22552 16932 22558 16944
rect 22865 16941 22877 16944
rect 22911 16941 22923 16975
rect 22865 16935 22923 16941
rect 23138 16932 23144 16984
rect 23196 16972 23202 16984
rect 23417 16975 23475 16981
rect 23417 16972 23429 16975
rect 23196 16944 23429 16972
rect 23196 16932 23202 16944
rect 23417 16941 23429 16944
rect 23463 16941 23475 16975
rect 23417 16935 23475 16941
rect 20344 16876 21160 16904
rect 22405 16907 22463 16913
rect 20344 16864 20350 16876
rect 22405 16873 22417 16907
rect 22451 16904 22463 16907
rect 23230 16904 23236 16916
rect 22451 16876 23236 16904
rect 22451 16873 22463 16876
rect 22405 16867 22463 16873
rect 23230 16864 23236 16876
rect 23288 16864 23294 16916
rect 1061 16839 1119 16845
rect 1061 16805 1073 16839
rect 1107 16836 1119 16839
rect 2530 16836 2536 16848
rect 1107 16808 2536 16836
rect 1107 16805 1119 16808
rect 1061 16799 1119 16805
rect 2530 16796 2536 16808
rect 2588 16796 2594 16848
rect 8513 16839 8571 16845
rect 8513 16805 8525 16839
rect 8559 16836 8571 16839
rect 9706 16836 9712 16848
rect 8559 16808 9712 16836
rect 8559 16805 8571 16808
rect 8513 16799 8571 16805
rect 9706 16796 9712 16808
rect 9764 16796 9770 16848
rect 14766 16836 14772 16848
rect 14727 16808 14772 16836
rect 14766 16796 14772 16808
rect 14824 16796 14830 16848
rect 17529 16839 17587 16845
rect 17529 16805 17541 16839
rect 17575 16836 17587 16839
rect 17710 16836 17716 16848
rect 17575 16808 17716 16836
rect 17575 16805 17587 16808
rect 17529 16799 17587 16805
rect 17710 16796 17716 16808
rect 17768 16796 17774 16848
rect 19366 16836 19372 16848
rect 19327 16808 19372 16836
rect 19366 16796 19372 16808
rect 19424 16796 19430 16848
rect 24058 16836 24064 16848
rect 24019 16808 24064 16836
rect 24058 16796 24064 16808
rect 24116 16796 24122 16848
rect 27922 16796 27928 16848
rect 27980 16836 27986 16848
rect 28109 16839 28167 16845
rect 28109 16836 28121 16839
rect 27980 16808 28121 16836
rect 27980 16796 27986 16808
rect 28109 16805 28121 16808
rect 28155 16805 28167 16839
rect 28109 16799 28167 16805
rect 400 16746 31680 16768
rect 400 16694 3510 16746
rect 3562 16694 3574 16746
rect 3626 16694 3638 16746
rect 3690 16694 3702 16746
rect 3754 16694 3766 16746
rect 3818 16694 31680 16746
rect 400 16672 31680 16694
rect 3910 16632 3916 16644
rect 3871 16604 3916 16632
rect 3910 16592 3916 16604
rect 3968 16592 3974 16644
rect 4094 16632 4100 16644
rect 4055 16604 4100 16632
rect 4094 16592 4100 16604
rect 4152 16592 4158 16644
rect 4278 16632 4284 16644
rect 4239 16604 4284 16632
rect 4278 16592 4284 16604
rect 4336 16592 4342 16644
rect 4462 16632 4468 16644
rect 4423 16604 4468 16632
rect 4462 16592 4468 16604
rect 4520 16592 4526 16644
rect 5198 16632 5204 16644
rect 5159 16604 5204 16632
rect 5198 16592 5204 16604
rect 5256 16592 5262 16644
rect 5382 16592 5388 16644
rect 5440 16632 5446 16644
rect 5569 16635 5627 16641
rect 5569 16632 5581 16635
rect 5440 16604 5581 16632
rect 5440 16592 5446 16604
rect 5569 16601 5581 16604
rect 5615 16601 5627 16635
rect 5750 16632 5756 16644
rect 5711 16604 5756 16632
rect 5569 16595 5627 16601
rect 5750 16592 5756 16604
rect 5808 16592 5814 16644
rect 7406 16632 7412 16644
rect 7367 16604 7412 16632
rect 7406 16592 7412 16604
rect 7464 16592 7470 16644
rect 7590 16632 7596 16644
rect 7551 16604 7596 16632
rect 7590 16592 7596 16604
rect 7648 16592 7654 16644
rect 14950 16592 14956 16644
rect 15008 16632 15014 16644
rect 15321 16635 15379 16641
rect 15321 16632 15333 16635
rect 15008 16604 15333 16632
rect 15008 16592 15014 16604
rect 15321 16601 15333 16604
rect 15367 16601 15379 16635
rect 15962 16632 15968 16644
rect 15923 16604 15968 16632
rect 15321 16595 15379 16601
rect 15962 16592 15968 16604
rect 16020 16592 16026 16644
rect 16425 16635 16483 16641
rect 16425 16601 16437 16635
rect 16471 16632 16483 16635
rect 16514 16632 16520 16644
rect 16471 16604 16520 16632
rect 16471 16601 16483 16604
rect 16425 16595 16483 16601
rect 16514 16592 16520 16604
rect 16572 16592 16578 16644
rect 18170 16592 18176 16644
rect 18228 16632 18234 16644
rect 18265 16635 18323 16641
rect 18265 16632 18277 16635
rect 18228 16604 18277 16632
rect 18228 16592 18234 16604
rect 18265 16601 18277 16604
rect 18311 16601 18323 16635
rect 20286 16632 20292 16644
rect 20247 16604 20292 16632
rect 18265 16595 18323 16601
rect 20286 16592 20292 16604
rect 20344 16592 20350 16644
rect 20473 16635 20531 16641
rect 20473 16601 20485 16635
rect 20519 16632 20531 16635
rect 20746 16632 20752 16644
rect 20519 16604 20752 16632
rect 20519 16601 20531 16604
rect 20473 16595 20531 16601
rect 20746 16592 20752 16604
rect 20804 16592 20810 16644
rect 20841 16635 20899 16641
rect 20841 16601 20853 16635
rect 20887 16632 20899 16635
rect 21390 16632 21396 16644
rect 20887 16604 21396 16632
rect 20887 16601 20899 16604
rect 20841 16595 20899 16601
rect 21390 16592 21396 16604
rect 21448 16592 21454 16644
rect 22494 16632 22500 16644
rect 22455 16604 22500 16632
rect 22494 16592 22500 16604
rect 22552 16592 22558 16644
rect 23230 16632 23236 16644
rect 23191 16604 23236 16632
rect 23230 16592 23236 16604
rect 23288 16592 23294 16644
rect 23693 16635 23751 16641
rect 23693 16601 23705 16635
rect 23739 16632 23751 16635
rect 24150 16632 24156 16644
rect 23739 16604 24156 16632
rect 23739 16601 23751 16604
rect 23693 16595 23751 16601
rect 24150 16592 24156 16604
rect 24208 16632 24214 16644
rect 24245 16635 24303 16641
rect 24245 16632 24257 16635
rect 24208 16604 24257 16632
rect 24208 16592 24214 16604
rect 24245 16601 24257 16604
rect 24291 16601 24303 16635
rect 26910 16632 26916 16644
rect 26871 16604 26916 16632
rect 24245 16595 24303 16601
rect 26910 16592 26916 16604
rect 26968 16592 26974 16644
rect 27830 16632 27836 16644
rect 27791 16604 27836 16632
rect 27830 16592 27836 16604
rect 27888 16592 27894 16644
rect 27922 16592 27928 16644
rect 27980 16632 27986 16644
rect 28201 16635 28259 16641
rect 28201 16632 28213 16635
rect 27980 16604 28213 16632
rect 27980 16592 27986 16604
rect 28201 16601 28213 16604
rect 28247 16601 28259 16635
rect 28201 16595 28259 16601
rect 3545 16567 3603 16573
rect 3545 16564 3557 16567
rect 3284 16536 3557 16564
rect 877 16499 935 16505
rect 877 16465 889 16499
rect 923 16496 935 16499
rect 2441 16499 2499 16505
rect 923 16468 1932 16496
rect 923 16465 935 16468
rect 877 16459 935 16465
rect 1904 16440 1932 16468
rect 2441 16465 2453 16499
rect 2487 16496 2499 16499
rect 2487 16468 3036 16496
rect 2487 16465 2499 16468
rect 2441 16459 2499 16465
rect 1613 16431 1671 16437
rect 1613 16397 1625 16431
rect 1659 16397 1671 16431
rect 1794 16428 1800 16440
rect 1755 16400 1800 16428
rect 1613 16391 1671 16397
rect 1153 16363 1211 16369
rect 1153 16329 1165 16363
rect 1199 16329 1211 16363
rect 1628 16360 1656 16391
rect 1794 16388 1800 16400
rect 1852 16388 1858 16440
rect 1886 16388 1892 16440
rect 1944 16428 1950 16440
rect 1981 16431 2039 16437
rect 1981 16428 1993 16431
rect 1944 16400 1993 16428
rect 1944 16388 1950 16400
rect 1981 16397 1993 16400
rect 2027 16397 2039 16431
rect 2530 16428 2536 16440
rect 2491 16400 2536 16428
rect 1981 16391 2039 16397
rect 2530 16388 2536 16400
rect 2588 16388 2594 16440
rect 1702 16360 1708 16372
rect 1615 16332 1708 16360
rect 1153 16323 1211 16329
rect 966 16292 972 16304
rect 927 16264 972 16292
rect 966 16252 972 16264
rect 1024 16292 1030 16304
rect 1168 16292 1196 16323
rect 1702 16320 1708 16332
rect 1760 16360 1766 16372
rect 3008 16369 3036 16468
rect 3284 16440 3312 16536
rect 3545 16533 3557 16536
rect 3591 16533 3603 16567
rect 5474 16564 5480 16576
rect 5435 16536 5480 16564
rect 3545 16527 3603 16533
rect 5474 16524 5480 16536
rect 5532 16524 5538 16576
rect 3361 16499 3419 16505
rect 3361 16465 3373 16499
rect 3407 16465 3419 16499
rect 3361 16459 3419 16465
rect 3177 16431 3235 16437
rect 3177 16397 3189 16431
rect 3223 16428 3235 16431
rect 3266 16428 3272 16440
rect 3223 16400 3272 16428
rect 3223 16397 3235 16400
rect 3177 16391 3235 16397
rect 3266 16388 3272 16400
rect 3324 16388 3330 16440
rect 3376 16428 3404 16459
rect 4370 16456 4376 16508
rect 4428 16496 4434 16508
rect 5768 16496 5796 16592
rect 11730 16524 11736 16576
rect 11788 16564 11794 16576
rect 12193 16567 12251 16573
rect 12193 16564 12205 16567
rect 11788 16536 12205 16564
rect 11788 16524 11794 16536
rect 12193 16533 12205 16536
rect 12239 16533 12251 16567
rect 12193 16527 12251 16533
rect 4428 16468 5796 16496
rect 4428 16456 4434 16468
rect 6854 16456 6860 16508
rect 6912 16496 6918 16508
rect 6912 16468 8188 16496
rect 6912 16456 6918 16468
rect 3729 16431 3787 16437
rect 3729 16428 3741 16431
rect 3376 16400 3741 16428
rect 3729 16397 3741 16400
rect 3775 16428 3787 16431
rect 4278 16428 4284 16440
rect 3775 16400 4284 16428
rect 3775 16397 3787 16400
rect 3729 16391 3787 16397
rect 4278 16388 4284 16400
rect 4336 16388 4342 16440
rect 7222 16428 7228 16440
rect 7135 16400 7228 16428
rect 7222 16388 7228 16400
rect 7280 16428 7286 16440
rect 7777 16431 7835 16437
rect 7777 16428 7789 16431
rect 7280 16400 7789 16428
rect 7280 16388 7286 16400
rect 7777 16397 7789 16400
rect 7823 16397 7835 16431
rect 8160 16428 8188 16468
rect 8234 16456 8240 16508
rect 8292 16496 8298 16508
rect 8329 16499 8387 16505
rect 8329 16496 8341 16499
rect 8292 16468 8341 16496
rect 8292 16456 8298 16468
rect 8329 16465 8341 16468
rect 8375 16496 8387 16499
rect 10445 16499 10503 16505
rect 10445 16496 10457 16499
rect 8375 16468 10457 16496
rect 8375 16465 8387 16468
rect 8329 16459 8387 16465
rect 10445 16465 10457 16468
rect 10491 16465 10503 16499
rect 13938 16496 13944 16508
rect 10445 16459 10503 16465
rect 11380 16468 13944 16496
rect 8418 16428 8424 16440
rect 8160 16400 8424 16428
rect 7777 16391 7835 16397
rect 8418 16388 8424 16400
rect 8476 16388 8482 16440
rect 9706 16388 9712 16440
rect 9764 16428 9770 16440
rect 11380 16428 11408 16468
rect 13938 16456 13944 16468
rect 13996 16456 14002 16508
rect 14493 16499 14551 16505
rect 14493 16465 14505 16499
rect 14539 16496 14551 16499
rect 14953 16499 15011 16505
rect 14953 16496 14965 16499
rect 14539 16468 14965 16496
rect 14539 16465 14551 16468
rect 14493 16459 14551 16465
rect 14953 16465 14965 16468
rect 14999 16496 15011 16499
rect 16149 16499 16207 16505
rect 16149 16496 16161 16499
rect 14999 16468 16161 16496
rect 14999 16465 15011 16468
rect 14953 16459 15011 16465
rect 16149 16465 16161 16468
rect 16195 16496 16207 16499
rect 16422 16496 16428 16508
rect 16195 16468 16428 16496
rect 16195 16465 16207 16468
rect 16149 16459 16207 16465
rect 16422 16456 16428 16468
rect 16480 16456 16486 16508
rect 16532 16496 16560 16592
rect 17526 16524 17532 16576
rect 17584 16564 17590 16576
rect 18081 16567 18139 16573
rect 18081 16564 18093 16567
rect 17584 16536 18093 16564
rect 17584 16524 17590 16536
rect 18081 16533 18093 16536
rect 18127 16564 18139 16567
rect 18998 16564 19004 16576
rect 18127 16536 19004 16564
rect 18127 16533 18139 16536
rect 18081 16527 18139 16533
rect 18998 16524 19004 16536
rect 19056 16524 19062 16576
rect 20930 16564 20936 16576
rect 20891 16536 20936 16564
rect 20930 16524 20936 16536
rect 20988 16524 20994 16576
rect 23506 16524 23512 16576
rect 23564 16564 23570 16576
rect 23785 16567 23843 16573
rect 23785 16564 23797 16567
rect 23564 16536 23797 16564
rect 23564 16524 23570 16536
rect 23785 16533 23797 16536
rect 23831 16564 23843 16567
rect 23831 16536 24012 16564
rect 23831 16533 23843 16536
rect 23785 16527 23843 16533
rect 19274 16496 19280 16508
rect 16532 16468 19280 16496
rect 19274 16456 19280 16468
rect 19332 16456 19338 16508
rect 22405 16499 22463 16505
rect 22405 16465 22417 16499
rect 22451 16496 22463 16499
rect 23322 16496 23328 16508
rect 22451 16468 23328 16496
rect 22451 16465 22463 16468
rect 22405 16459 22463 16465
rect 23322 16456 23328 16468
rect 23380 16496 23386 16508
rect 23417 16499 23475 16505
rect 23417 16496 23429 16499
rect 23380 16468 23429 16496
rect 23380 16456 23386 16468
rect 23417 16465 23429 16468
rect 23463 16496 23475 16499
rect 23984 16496 24012 16536
rect 24058 16524 24064 16576
rect 24116 16564 24122 16576
rect 24116 16536 25024 16564
rect 24116 16524 24122 16536
rect 24889 16499 24947 16505
rect 24889 16496 24901 16499
rect 23463 16468 23874 16496
rect 23984 16468 24901 16496
rect 23463 16465 23475 16468
rect 23417 16459 23475 16465
rect 11730 16428 11736 16440
rect 9764 16400 11408 16428
rect 11691 16400 11736 16428
rect 9764 16388 9770 16400
rect 11730 16388 11736 16400
rect 11788 16388 11794 16440
rect 12558 16388 12564 16440
rect 12616 16428 12622 16440
rect 14217 16431 14275 16437
rect 14217 16428 14229 16431
rect 12616 16400 14229 16428
rect 12616 16388 12622 16400
rect 14217 16397 14229 16400
rect 14263 16428 14275 16431
rect 14769 16431 14827 16437
rect 14769 16428 14781 16431
rect 14263 16400 14781 16428
rect 14263 16397 14275 16400
rect 14217 16391 14275 16397
rect 14769 16397 14781 16400
rect 14815 16397 14827 16431
rect 14769 16391 14827 16397
rect 17161 16431 17219 16437
rect 17161 16397 17173 16431
rect 17207 16428 17219 16431
rect 17434 16428 17440 16440
rect 17207 16400 17440 16428
rect 17207 16397 17219 16400
rect 17161 16391 17219 16397
rect 17434 16388 17440 16400
rect 17492 16388 17498 16440
rect 17710 16428 17716 16440
rect 17671 16400 17716 16428
rect 17710 16388 17716 16400
rect 17768 16388 17774 16440
rect 19366 16428 19372 16440
rect 19327 16400 19372 16428
rect 19366 16388 19372 16400
rect 19424 16388 19430 16440
rect 19737 16431 19795 16437
rect 19737 16397 19749 16431
rect 19783 16397 19795 16431
rect 19737 16391 19795 16397
rect 2717 16363 2775 16369
rect 2717 16360 2729 16363
rect 1760 16332 2729 16360
rect 1760 16320 1766 16332
rect 2717 16329 2729 16332
rect 2763 16329 2775 16363
rect 2717 16323 2775 16329
rect 2993 16363 3051 16369
rect 2993 16329 3005 16363
rect 3039 16360 3051 16363
rect 3358 16360 3364 16372
rect 3039 16332 3364 16360
rect 3039 16329 3051 16332
rect 2993 16323 3051 16329
rect 3358 16320 3364 16332
rect 3416 16320 3422 16372
rect 6673 16363 6731 16369
rect 6673 16329 6685 16363
rect 6719 16360 6731 16363
rect 7314 16360 7320 16372
rect 6719 16332 7320 16360
rect 6719 16329 6731 16332
rect 6673 16323 6731 16329
rect 7314 16320 7320 16332
rect 7372 16320 7378 16372
rect 7958 16320 7964 16372
rect 8016 16360 8022 16372
rect 8145 16363 8203 16369
rect 8145 16360 8157 16363
rect 8016 16332 8157 16360
rect 8016 16320 8022 16332
rect 8145 16329 8157 16332
rect 8191 16360 8203 16363
rect 8697 16363 8755 16369
rect 8697 16360 8709 16363
rect 8191 16332 8709 16360
rect 8191 16329 8203 16332
rect 8145 16323 8203 16329
rect 8697 16329 8709 16332
rect 8743 16329 8755 16363
rect 12098 16360 12104 16372
rect 12011 16332 12104 16360
rect 8697 16323 8755 16329
rect 12098 16320 12104 16332
rect 12156 16360 12162 16372
rect 12377 16363 12435 16369
rect 12377 16360 12389 16363
rect 12156 16332 12389 16360
rect 12156 16320 12162 16332
rect 12377 16329 12389 16332
rect 12423 16329 12435 16363
rect 12377 16323 12435 16329
rect 18725 16363 18783 16369
rect 18725 16329 18737 16363
rect 18771 16360 18783 16363
rect 19458 16360 19464 16372
rect 18771 16332 19464 16360
rect 18771 16329 18783 16332
rect 18725 16323 18783 16329
rect 19458 16320 19464 16332
rect 19516 16320 19522 16372
rect 6762 16292 6768 16304
rect 1024 16264 1196 16292
rect 6723 16264 6768 16292
rect 1024 16252 1030 16264
rect 6762 16252 6768 16264
rect 6820 16252 6826 16304
rect 10534 16252 10540 16304
rect 10592 16292 10598 16304
rect 14766 16292 14772 16304
rect 10592 16264 14772 16292
rect 10592 16252 10598 16264
rect 14766 16252 14772 16264
rect 14824 16292 14830 16304
rect 15137 16295 15195 16301
rect 15137 16292 15149 16295
rect 14824 16264 15149 16292
rect 14824 16252 14830 16264
rect 15137 16261 15149 16264
rect 15183 16261 15195 16295
rect 15137 16255 15195 16261
rect 18446 16252 18452 16304
rect 18504 16292 18510 16304
rect 18541 16295 18599 16301
rect 18541 16292 18553 16295
rect 18504 16264 18553 16292
rect 18504 16252 18510 16264
rect 18541 16261 18553 16264
rect 18587 16292 18599 16295
rect 19752 16292 19780 16391
rect 19826 16388 19832 16440
rect 19884 16428 19890 16440
rect 23138 16428 23144 16440
rect 19884 16400 19929 16428
rect 22696 16400 23144 16428
rect 19884 16388 19890 16400
rect 21574 16320 21580 16372
rect 21632 16360 21638 16372
rect 22696 16369 22724 16400
rect 23138 16388 23144 16400
rect 23196 16388 23202 16440
rect 23846 16428 23874 16468
rect 24889 16465 24901 16468
rect 24935 16465 24947 16499
rect 24889 16459 24947 16465
rect 24150 16428 24156 16440
rect 23846 16400 24156 16428
rect 24150 16388 24156 16400
rect 24208 16428 24214 16440
rect 24429 16431 24487 16437
rect 24429 16428 24441 16431
rect 24208 16400 24441 16428
rect 24208 16388 24214 16400
rect 24429 16397 24441 16400
rect 24475 16397 24487 16431
rect 24610 16428 24616 16440
rect 24571 16400 24616 16428
rect 24429 16391 24487 16397
rect 24610 16388 24616 16400
rect 24668 16388 24674 16440
rect 24996 16437 25024 16536
rect 25901 16499 25959 16505
rect 25901 16465 25913 16499
rect 25947 16496 25959 16499
rect 26174 16496 26180 16508
rect 25947 16468 26180 16496
rect 25947 16465 25959 16468
rect 25901 16459 25959 16465
rect 26174 16456 26180 16468
rect 26232 16456 26238 16508
rect 26928 16496 26956 16592
rect 27738 16564 27744 16576
rect 27699 16536 27744 16564
rect 27738 16524 27744 16536
rect 27796 16524 27802 16576
rect 26284 16468 26956 16496
rect 24981 16431 25039 16437
rect 24981 16397 24993 16431
rect 25027 16428 25039 16431
rect 25254 16428 25260 16440
rect 25027 16400 25260 16428
rect 25027 16397 25039 16400
rect 24981 16391 25039 16397
rect 25254 16388 25260 16400
rect 25312 16388 25318 16440
rect 25438 16388 25444 16440
rect 25496 16428 25502 16440
rect 26284 16437 26312 16468
rect 26269 16431 26327 16437
rect 26269 16428 26281 16431
rect 25496 16400 26281 16428
rect 25496 16388 25502 16400
rect 26269 16397 26281 16400
rect 26315 16397 26327 16431
rect 26269 16391 26327 16397
rect 26453 16431 26511 16437
rect 26453 16397 26465 16431
rect 26499 16397 26511 16431
rect 26453 16391 26511 16397
rect 29949 16431 30007 16437
rect 29949 16397 29961 16431
rect 29995 16428 30007 16431
rect 30038 16428 30044 16440
rect 29995 16400 30044 16428
rect 29995 16397 30007 16400
rect 29949 16391 30007 16397
rect 22681 16363 22739 16369
rect 22681 16360 22693 16363
rect 21632 16332 22693 16360
rect 21632 16320 21638 16332
rect 22681 16329 22693 16332
rect 22727 16329 22739 16363
rect 22681 16323 22739 16329
rect 22954 16320 22960 16372
rect 23012 16360 23018 16372
rect 23049 16363 23107 16369
rect 23049 16360 23061 16363
rect 23012 16332 23061 16360
rect 23012 16320 23018 16332
rect 23049 16329 23061 16332
rect 23095 16360 23107 16363
rect 25717 16363 25775 16369
rect 25717 16360 25729 16363
rect 23095 16332 25729 16360
rect 23095 16329 23107 16332
rect 23049 16323 23107 16329
rect 25717 16329 25729 16332
rect 25763 16360 25775 16363
rect 25763 16332 26036 16360
rect 25763 16329 25775 16332
rect 25717 16323 25775 16329
rect 18587 16264 19780 16292
rect 18587 16261 18599 16264
rect 18541 16255 18599 16261
rect 20470 16252 20476 16304
rect 20528 16292 20534 16304
rect 20565 16295 20623 16301
rect 20565 16292 20577 16295
rect 20528 16264 20577 16292
rect 20528 16252 20534 16264
rect 20565 16261 20577 16264
rect 20611 16261 20623 16295
rect 26008 16292 26036 16332
rect 26174 16320 26180 16372
rect 26232 16360 26238 16372
rect 26468 16360 26496 16391
rect 30038 16388 30044 16400
rect 30096 16428 30102 16440
rect 30317 16431 30375 16437
rect 30317 16428 30329 16431
rect 30096 16400 30329 16428
rect 30096 16388 30102 16400
rect 30317 16397 30329 16400
rect 30363 16397 30375 16431
rect 30317 16391 30375 16397
rect 26232 16332 26496 16360
rect 26232 16320 26238 16332
rect 26085 16295 26143 16301
rect 26085 16292 26097 16295
rect 26008 16264 26097 16292
rect 20565 16255 20623 16261
rect 26085 16261 26097 16264
rect 26131 16261 26143 16295
rect 28014 16292 28020 16304
rect 27975 16264 28020 16292
rect 26085 16255 26143 16261
rect 28014 16252 28020 16264
rect 28072 16252 28078 16304
rect 29946 16292 29952 16304
rect 29907 16264 29952 16292
rect 29946 16252 29952 16264
rect 30004 16292 30010 16304
rect 30133 16295 30191 16301
rect 30133 16292 30145 16295
rect 30004 16264 30145 16292
rect 30004 16252 30010 16264
rect 30133 16261 30145 16264
rect 30179 16261 30191 16295
rect 30133 16255 30191 16261
rect 400 16202 31680 16224
rect 400 16150 18870 16202
rect 18922 16150 18934 16202
rect 18986 16150 18998 16202
rect 19050 16150 19062 16202
rect 19114 16150 19126 16202
rect 19178 16150 31680 16202
rect 400 16128 31680 16150
rect 1702 16088 1708 16100
rect 1663 16060 1708 16088
rect 1702 16048 1708 16060
rect 1760 16048 1766 16100
rect 7314 16048 7320 16100
rect 7372 16088 7378 16100
rect 9249 16091 9307 16097
rect 9249 16088 9261 16091
rect 7372 16060 9261 16088
rect 7372 16048 7378 16060
rect 9249 16057 9261 16060
rect 9295 16088 9307 16091
rect 9798 16088 9804 16100
rect 9295 16060 9804 16088
rect 9295 16057 9307 16060
rect 9249 16051 9307 16057
rect 9798 16048 9804 16060
rect 9856 16048 9862 16100
rect 18357 16091 18415 16097
rect 18357 16057 18369 16091
rect 18403 16088 18415 16091
rect 18722 16088 18728 16100
rect 18403 16060 18728 16088
rect 18403 16057 18415 16060
rect 18357 16051 18415 16057
rect 18722 16048 18728 16060
rect 18780 16048 18786 16100
rect 19274 16088 19280 16100
rect 19235 16060 19280 16088
rect 19274 16048 19280 16060
rect 19332 16048 19338 16100
rect 22126 16048 22132 16100
rect 22184 16088 22190 16100
rect 22184 16060 24012 16088
rect 22184 16048 22190 16060
rect 1610 16020 1616 16032
rect 1571 15992 1616 16020
rect 1610 15980 1616 15992
rect 1668 15980 1674 16032
rect 6762 16020 6768 16032
rect 1996 15992 6768 16020
rect 1996 15964 2024 15992
rect 6762 15980 6768 15992
rect 6820 15980 6826 16032
rect 1150 15952 1156 15964
rect 1111 15924 1156 15952
rect 1150 15912 1156 15924
rect 1208 15912 1214 15964
rect 1978 15952 1984 15964
rect 1891 15924 1984 15952
rect 1978 15912 1984 15924
rect 2036 15912 2042 15964
rect 3266 15912 3272 15964
rect 3324 15952 3330 15964
rect 3361 15955 3419 15961
rect 3361 15952 3373 15955
rect 3324 15924 3373 15952
rect 3324 15912 3330 15924
rect 3361 15921 3373 15924
rect 3407 15921 3419 15955
rect 3361 15915 3419 15921
rect 3545 15955 3603 15961
rect 3545 15921 3557 15955
rect 3591 15952 3603 15955
rect 4002 15952 4008 15964
rect 3591 15924 4008 15952
rect 3591 15921 3603 15924
rect 3545 15915 3603 15921
rect 4002 15912 4008 15924
rect 4060 15912 4066 15964
rect 5750 15912 5756 15964
rect 5808 15952 5814 15964
rect 5937 15955 5995 15961
rect 5937 15952 5949 15955
rect 5808 15924 5949 15952
rect 5808 15912 5814 15924
rect 5937 15921 5949 15924
rect 5983 15921 5995 15955
rect 6302 15952 6308 15964
rect 6263 15924 6308 15952
rect 5937 15915 5995 15921
rect 1429 15887 1487 15893
rect 1429 15853 1441 15887
rect 1475 15884 1487 15887
rect 2254 15884 2260 15896
rect 1475 15856 2260 15884
rect 1475 15853 1487 15856
rect 1429 15847 1487 15853
rect 2254 15844 2260 15856
rect 2312 15844 2318 15896
rect 5842 15884 5848 15896
rect 5803 15856 5848 15884
rect 5842 15844 5848 15856
rect 5900 15844 5906 15896
rect 5952 15884 5980 15915
rect 6302 15912 6308 15924
rect 6360 15912 6366 15964
rect 6486 15952 6492 15964
rect 6399 15924 6492 15952
rect 6486 15912 6492 15924
rect 6544 15952 6550 15964
rect 7332 15952 7360 16048
rect 8234 16020 8240 16032
rect 7608 15992 8240 16020
rect 7608 15961 7636 15992
rect 8234 15980 8240 15992
rect 8292 15980 8298 16032
rect 8418 16020 8424 16032
rect 8379 15992 8424 16020
rect 8418 15980 8424 15992
rect 8476 16020 8482 16032
rect 8786 16020 8792 16032
rect 8476 15992 8792 16020
rect 8476 15980 8482 15992
rect 8786 15980 8792 15992
rect 8844 15980 8850 16032
rect 9065 16023 9123 16029
rect 9065 15989 9077 16023
rect 9111 16020 9123 16023
rect 9154 16020 9160 16032
rect 9111 15992 9160 16020
rect 9111 15989 9123 15992
rect 9065 15983 9123 15989
rect 9154 15980 9160 15992
rect 9212 15980 9218 16032
rect 12469 16023 12527 16029
rect 12469 15989 12481 16023
rect 12515 16020 12527 16023
rect 12558 16020 12564 16032
rect 12515 15992 12564 16020
rect 12515 15989 12527 15992
rect 12469 15983 12527 15989
rect 12558 15980 12564 15992
rect 12616 15980 12622 16032
rect 13754 15980 13760 16032
rect 13812 16020 13818 16032
rect 13812 15992 14214 16020
rect 13812 15980 13818 15992
rect 6544 15924 7360 15952
rect 7593 15955 7651 15961
rect 6544 15912 6550 15924
rect 7593 15921 7605 15955
rect 7639 15921 7651 15955
rect 7593 15915 7651 15921
rect 7682 15912 7688 15964
rect 7740 15952 7746 15964
rect 7777 15955 7835 15961
rect 7777 15952 7789 15955
rect 7740 15924 7789 15952
rect 7740 15912 7746 15924
rect 7777 15921 7789 15924
rect 7823 15921 7835 15955
rect 10718 15952 10724 15964
rect 7777 15915 7835 15921
rect 8252 15924 10724 15952
rect 6946 15884 6952 15896
rect 5952 15856 6952 15884
rect 6946 15844 6952 15856
rect 7004 15884 7010 15896
rect 7406 15884 7412 15896
rect 7004 15856 7412 15884
rect 7004 15844 7010 15856
rect 7406 15844 7412 15856
rect 7464 15884 7470 15896
rect 7869 15887 7927 15893
rect 7869 15884 7881 15887
rect 7464 15856 7881 15884
rect 7464 15844 7470 15856
rect 7869 15853 7881 15856
rect 7915 15853 7927 15887
rect 7869 15847 7927 15853
rect 7038 15776 7044 15828
rect 7096 15816 7102 15828
rect 8252 15816 8280 15924
rect 10718 15912 10724 15924
rect 10776 15912 10782 15964
rect 10994 15912 11000 15964
rect 11052 15952 11058 15964
rect 11917 15955 11975 15961
rect 11917 15952 11929 15955
rect 11052 15924 11929 15952
rect 11052 15912 11058 15924
rect 11917 15921 11929 15924
rect 11963 15921 11975 15955
rect 12098 15952 12104 15964
rect 12059 15924 12104 15952
rect 11917 15915 11975 15921
rect 12098 15912 12104 15924
rect 12156 15912 12162 15964
rect 14186 15952 14214 15992
rect 15226 15980 15232 16032
rect 15284 16020 15290 16032
rect 15284 15992 15732 16020
rect 15284 15980 15290 15992
rect 15505 15955 15563 15961
rect 15505 15952 15517 15955
rect 14186 15924 15517 15952
rect 15505 15921 15517 15924
rect 15551 15952 15563 15955
rect 15594 15952 15600 15964
rect 15551 15924 15600 15952
rect 15551 15921 15563 15924
rect 15505 15915 15563 15921
rect 15594 15912 15600 15924
rect 15652 15912 15658 15964
rect 15704 15961 15732 15992
rect 15962 15980 15968 16032
rect 16020 16020 16026 16032
rect 16057 16023 16115 16029
rect 16057 16020 16069 16023
rect 16020 15992 16069 16020
rect 16020 15980 16026 15992
rect 16057 15989 16069 15992
rect 16103 16020 16115 16023
rect 17434 16020 17440 16032
rect 16103 15992 17440 16020
rect 16103 15989 16115 15992
rect 16057 15983 16115 15989
rect 17434 15980 17440 15992
rect 17492 15980 17498 16032
rect 17710 15980 17716 16032
rect 17768 16020 17774 16032
rect 18449 16023 18507 16029
rect 18449 16020 18461 16023
rect 17768 15992 18461 16020
rect 17768 15980 17774 15992
rect 18449 15989 18461 15992
rect 18495 15989 18507 16023
rect 18449 15983 18507 15989
rect 22586 15980 22592 16032
rect 22644 15980 22650 16032
rect 23984 16029 24012 16060
rect 24058 16048 24064 16100
rect 24116 16088 24122 16100
rect 24245 16091 24303 16097
rect 24245 16088 24257 16091
rect 24116 16060 24257 16088
rect 24116 16048 24122 16060
rect 24245 16057 24257 16060
rect 24291 16057 24303 16091
rect 26726 16088 26732 16100
rect 26639 16060 26732 16088
rect 24245 16051 24303 16057
rect 26726 16048 26732 16060
rect 26784 16088 26790 16100
rect 27278 16088 27284 16100
rect 26784 16060 27284 16088
rect 26784 16048 26790 16060
rect 27278 16048 27284 16060
rect 27336 16048 27342 16100
rect 23969 16023 24027 16029
rect 23969 15989 23981 16023
rect 24015 16020 24027 16023
rect 25438 16020 25444 16032
rect 24015 15992 25444 16020
rect 24015 15989 24027 15992
rect 23969 15983 24027 15989
rect 25438 15980 25444 15992
rect 25496 15980 25502 16032
rect 27554 16020 27560 16032
rect 27515 15992 27560 16020
rect 27554 15980 27560 15992
rect 27612 15980 27618 16032
rect 15689 15955 15747 15961
rect 15689 15921 15701 15955
rect 15735 15921 15747 15955
rect 19458 15952 19464 15964
rect 19371 15924 19464 15952
rect 15689 15915 15747 15921
rect 19458 15912 19464 15924
rect 19516 15952 19522 15964
rect 22310 15952 22316 15964
rect 19516 15924 22316 15952
rect 19516 15912 19522 15924
rect 22310 15912 22316 15924
rect 22368 15912 22374 15964
rect 23874 15912 23880 15964
rect 23932 15952 23938 15964
rect 25806 15952 25812 15964
rect 23932 15924 25812 15952
rect 23932 15912 23938 15924
rect 25806 15912 25812 15924
rect 25864 15912 25870 15964
rect 28198 15952 28204 15964
rect 28159 15924 28204 15952
rect 28198 15912 28204 15924
rect 28256 15912 28262 15964
rect 28474 15912 28480 15964
rect 28532 15952 28538 15964
rect 28569 15955 28627 15961
rect 28569 15952 28581 15955
rect 28532 15924 28581 15952
rect 28532 15912 28538 15924
rect 28569 15921 28581 15924
rect 28615 15921 28627 15955
rect 28569 15915 28627 15921
rect 12282 15844 12288 15896
rect 12340 15884 12346 15896
rect 18081 15887 18139 15893
rect 18081 15884 18093 15887
rect 12340 15856 18093 15884
rect 12340 15844 12346 15856
rect 18081 15853 18093 15856
rect 18127 15884 18139 15887
rect 18538 15884 18544 15896
rect 18127 15856 18544 15884
rect 18127 15853 18139 15856
rect 18081 15847 18139 15853
rect 18538 15844 18544 15856
rect 18596 15844 18602 15896
rect 19093 15887 19151 15893
rect 19093 15853 19105 15887
rect 19139 15884 19151 15887
rect 19826 15884 19832 15896
rect 19139 15856 19832 15884
rect 19139 15853 19151 15856
rect 19093 15847 19151 15853
rect 19826 15844 19832 15856
rect 19884 15844 19890 15896
rect 21850 15884 21856 15896
rect 21811 15856 21856 15884
rect 21850 15844 21856 15856
rect 21908 15844 21914 15896
rect 22218 15884 22224 15896
rect 22179 15856 22224 15884
rect 22218 15844 22224 15856
rect 22276 15844 22282 15896
rect 28106 15884 28112 15896
rect 28067 15856 28112 15884
rect 28106 15844 28112 15856
rect 28164 15844 28170 15896
rect 28382 15844 28388 15896
rect 28440 15884 28446 15896
rect 28661 15887 28719 15893
rect 28661 15884 28673 15887
rect 28440 15856 28673 15884
rect 28440 15844 28446 15856
rect 28661 15853 28673 15856
rect 28707 15853 28719 15887
rect 28661 15847 28719 15853
rect 7096 15788 8280 15816
rect 7096 15776 7102 15788
rect 8326 15776 8332 15828
rect 8384 15816 8390 15828
rect 9062 15816 9068 15828
rect 8384 15788 9068 15816
rect 8384 15776 8390 15788
rect 9062 15776 9068 15788
rect 9120 15816 9126 15828
rect 9341 15819 9399 15825
rect 9341 15816 9353 15819
rect 9120 15788 9353 15816
rect 9120 15776 9126 15788
rect 9341 15785 9353 15788
rect 9387 15785 9399 15819
rect 24610 15816 24616 15828
rect 9341 15779 9399 15785
rect 24076 15788 24616 15816
rect 24076 15760 24104 15788
rect 24610 15776 24616 15788
rect 24668 15776 24674 15828
rect 3358 15708 3364 15760
rect 3416 15748 3422 15760
rect 3637 15751 3695 15757
rect 3637 15748 3649 15751
rect 3416 15720 3649 15748
rect 3416 15708 3422 15720
rect 3637 15717 3649 15720
rect 3683 15717 3695 15751
rect 4738 15748 4744 15760
rect 4699 15720 4744 15748
rect 3637 15711 3695 15717
rect 4738 15708 4744 15720
rect 4796 15708 4802 15760
rect 5382 15748 5388 15760
rect 5343 15720 5388 15748
rect 5382 15708 5388 15720
rect 5440 15708 5446 15760
rect 9522 15748 9528 15760
rect 9483 15720 9528 15748
rect 9522 15708 9528 15720
rect 9580 15708 9586 15760
rect 10994 15748 11000 15760
rect 10955 15720 11000 15748
rect 10994 15708 11000 15720
rect 11052 15708 11058 15760
rect 18906 15748 18912 15760
rect 18867 15720 18912 15748
rect 18906 15708 18912 15720
rect 18964 15708 18970 15760
rect 18998 15708 19004 15760
rect 19056 15748 19062 15760
rect 21850 15748 21856 15760
rect 19056 15720 21856 15748
rect 19056 15708 19062 15720
rect 21850 15708 21856 15720
rect 21908 15748 21914 15760
rect 22402 15748 22408 15760
rect 21908 15720 22408 15748
rect 21908 15708 21914 15720
rect 22402 15708 22408 15720
rect 22460 15708 22466 15760
rect 24058 15708 24064 15760
rect 24116 15748 24122 15760
rect 26542 15748 26548 15760
rect 24116 15720 24161 15748
rect 26503 15720 26548 15748
rect 24116 15708 24122 15720
rect 26542 15708 26548 15720
rect 26600 15708 26606 15760
rect 400 15658 31680 15680
rect 400 15606 3510 15658
rect 3562 15606 3574 15658
rect 3626 15606 3638 15658
rect 3690 15606 3702 15658
rect 3754 15606 3766 15658
rect 3818 15606 31680 15658
rect 400 15584 31680 15606
rect 1061 15547 1119 15553
rect 1061 15513 1073 15547
rect 1107 15544 1119 15547
rect 1150 15544 1156 15556
rect 1107 15516 1156 15544
rect 1107 15513 1119 15516
rect 1061 15507 1119 15513
rect 1150 15504 1156 15516
rect 1208 15504 1214 15556
rect 1978 15544 1984 15556
rect 1939 15516 1984 15544
rect 1978 15504 1984 15516
rect 2036 15504 2042 15556
rect 2901 15547 2959 15553
rect 2901 15513 2913 15547
rect 2947 15544 2959 15547
rect 3453 15547 3511 15553
rect 3453 15544 3465 15547
rect 2947 15516 3465 15544
rect 2947 15513 2959 15516
rect 2901 15507 2959 15513
rect 3453 15513 3465 15516
rect 3499 15544 3511 15547
rect 4462 15544 4468 15556
rect 3499 15516 4468 15544
rect 3499 15513 3511 15516
rect 3453 15507 3511 15513
rect 4462 15504 4468 15516
rect 4520 15504 4526 15556
rect 4738 15504 4744 15556
rect 4796 15544 4802 15556
rect 4925 15547 4983 15553
rect 4925 15544 4937 15547
rect 4796 15516 4937 15544
rect 4796 15504 4802 15516
rect 4925 15513 4937 15516
rect 4971 15513 4983 15547
rect 5750 15544 5756 15556
rect 5711 15516 5756 15544
rect 4925 15507 4983 15513
rect 5750 15504 5756 15516
rect 5808 15504 5814 15556
rect 6213 15547 6271 15553
rect 6213 15513 6225 15547
rect 6259 15544 6271 15547
rect 6486 15544 6492 15556
rect 6259 15516 6492 15544
rect 6259 15513 6271 15516
rect 6213 15507 6271 15513
rect 6486 15504 6492 15516
rect 6544 15504 6550 15556
rect 6946 15544 6952 15556
rect 6907 15516 6952 15544
rect 6946 15504 6952 15516
rect 7004 15504 7010 15556
rect 7958 15544 7964 15556
rect 7919 15516 7964 15544
rect 7958 15504 7964 15516
rect 8016 15504 8022 15556
rect 10718 15544 10724 15556
rect 10679 15516 10724 15544
rect 10718 15504 10724 15516
rect 10776 15504 10782 15556
rect 10994 15544 11000 15556
rect 10955 15516 11000 15544
rect 10994 15504 11000 15516
rect 11052 15544 11058 15556
rect 11457 15547 11515 15553
rect 11457 15544 11469 15547
rect 11052 15516 11469 15544
rect 11052 15504 11058 15516
rect 11457 15513 11469 15516
rect 11503 15513 11515 15547
rect 11457 15507 11515 15513
rect 3913 15479 3971 15485
rect 3913 15445 3925 15479
rect 3959 15476 3971 15479
rect 4002 15476 4008 15488
rect 3959 15448 4008 15476
rect 3959 15445 3971 15448
rect 3913 15439 3971 15445
rect 4002 15436 4008 15448
rect 4060 15436 4066 15488
rect 4094 15436 4100 15488
rect 4152 15476 4158 15488
rect 4152 15448 4197 15476
rect 4152 15436 4158 15448
rect 4830 15436 4836 15488
rect 4888 15476 4894 15488
rect 5842 15476 5848 15488
rect 4888 15448 5848 15476
rect 4888 15436 4894 15448
rect 5842 15436 5848 15448
rect 5900 15436 5906 15488
rect 6857 15479 6915 15485
rect 6857 15445 6869 15479
rect 6903 15476 6915 15479
rect 9522 15476 9528 15488
rect 6903 15448 9528 15476
rect 6903 15445 6915 15448
rect 6857 15439 6915 15445
rect 2254 15340 2260 15352
rect 2167 15312 2260 15340
rect 2254 15300 2260 15312
rect 2312 15340 2318 15352
rect 3361 15343 3419 15349
rect 3361 15340 3373 15343
rect 2312 15312 3373 15340
rect 2312 15300 2318 15312
rect 3361 15309 3373 15312
rect 3407 15340 3419 15343
rect 4112 15340 4140 15436
rect 4278 15368 4284 15420
rect 4336 15408 4342 15420
rect 4465 15411 4523 15417
rect 4465 15408 4477 15411
rect 4336 15380 4477 15408
rect 4336 15368 4342 15380
rect 4465 15377 4477 15380
rect 4511 15408 4523 15411
rect 7225 15411 7283 15417
rect 4511 15380 4692 15408
rect 4511 15377 4523 15380
rect 4465 15371 4523 15377
rect 4664 15349 4692 15380
rect 7225 15377 7237 15411
rect 7271 15408 7283 15411
rect 7774 15408 7780 15420
rect 7271 15380 7780 15408
rect 7271 15377 7283 15380
rect 7225 15371 7283 15377
rect 7774 15368 7780 15380
rect 7832 15408 7838 15420
rect 8234 15408 8240 15420
rect 7832 15380 8240 15408
rect 7832 15368 7838 15380
rect 8234 15368 8240 15380
rect 8292 15368 8298 15420
rect 3407 15312 4140 15340
rect 4649 15343 4707 15349
rect 3407 15309 3419 15312
rect 3361 15303 3419 15309
rect 4649 15309 4661 15343
rect 4695 15309 4707 15343
rect 4649 15303 4707 15309
rect 4833 15343 4891 15349
rect 4833 15309 4845 15343
rect 4879 15340 4891 15343
rect 8326 15340 8332 15352
rect 4879 15312 5336 15340
rect 8287 15312 8332 15340
rect 4879 15309 4891 15312
rect 4833 15303 4891 15309
rect 3085 15275 3143 15281
rect 3085 15241 3097 15275
rect 3131 15272 3143 15275
rect 3177 15275 3235 15281
rect 3177 15272 3189 15275
rect 3131 15244 3189 15272
rect 3131 15241 3143 15244
rect 3085 15235 3143 15241
rect 3177 15241 3189 15244
rect 3223 15272 3235 15275
rect 3266 15272 3272 15284
rect 3223 15244 3272 15272
rect 3223 15241 3235 15244
rect 3177 15235 3235 15241
rect 3266 15232 3272 15244
rect 3324 15272 3330 15284
rect 4189 15275 4247 15281
rect 4189 15272 4201 15275
rect 3324 15244 4201 15272
rect 3324 15232 3330 15244
rect 4189 15241 4201 15244
rect 4235 15241 4247 15275
rect 4189 15235 4247 15241
rect 5308 15216 5336 15312
rect 8326 15300 8332 15312
rect 8384 15300 8390 15352
rect 8712 15349 8740 15448
rect 9522 15436 9528 15448
rect 9580 15436 9586 15488
rect 8697 15343 8755 15349
rect 8697 15309 8709 15343
rect 8743 15309 8755 15343
rect 8697 15303 8755 15309
rect 8789 15343 8847 15349
rect 8789 15309 8801 15343
rect 8835 15309 8847 15343
rect 11472 15340 11500 15507
rect 12098 15504 12104 15556
rect 12156 15544 12162 15556
rect 12561 15547 12619 15553
rect 12561 15544 12573 15547
rect 12156 15516 12573 15544
rect 12156 15504 12162 15516
rect 12561 15513 12573 15516
rect 12607 15513 12619 15547
rect 12561 15507 12619 15513
rect 14861 15547 14919 15553
rect 14861 15513 14873 15547
rect 14907 15544 14919 15547
rect 14950 15544 14956 15556
rect 14907 15516 14956 15544
rect 14907 15513 14919 15516
rect 14861 15507 14919 15513
rect 14950 15504 14956 15516
rect 15008 15504 15014 15556
rect 15962 15544 15968 15556
rect 15923 15516 15968 15544
rect 15962 15504 15968 15516
rect 16020 15504 16026 15556
rect 22126 15544 22132 15556
rect 22087 15516 22132 15544
rect 22126 15504 22132 15516
rect 22184 15544 22190 15556
rect 22310 15544 22316 15556
rect 22184 15516 22316 15544
rect 22184 15504 22190 15516
rect 22310 15504 22316 15516
rect 22368 15504 22374 15556
rect 22402 15504 22408 15556
rect 22460 15544 22466 15556
rect 23969 15547 24027 15553
rect 22460 15516 22505 15544
rect 22460 15504 22466 15516
rect 23969 15513 23981 15547
rect 24015 15544 24027 15547
rect 24242 15544 24248 15556
rect 24015 15516 24248 15544
rect 24015 15513 24027 15516
rect 23969 15507 24027 15513
rect 24242 15504 24248 15516
rect 24300 15544 24306 15556
rect 24521 15547 24579 15553
rect 24521 15544 24533 15547
rect 24300 15516 24533 15544
rect 24300 15504 24306 15516
rect 24521 15513 24533 15516
rect 24567 15513 24579 15547
rect 24521 15507 24579 15513
rect 26545 15547 26603 15553
rect 26545 15513 26557 15547
rect 26591 15544 26603 15547
rect 26726 15544 26732 15556
rect 26591 15516 26732 15544
rect 26591 15513 26603 15516
rect 26545 15507 26603 15513
rect 26726 15504 26732 15516
rect 26784 15504 26790 15556
rect 27186 15544 27192 15556
rect 26836 15516 27192 15544
rect 11730 15436 11736 15488
rect 11788 15476 11794 15488
rect 11914 15476 11920 15488
rect 11788 15448 11920 15476
rect 11788 15436 11794 15448
rect 11914 15436 11920 15448
rect 11972 15476 11978 15488
rect 12377 15479 12435 15485
rect 12377 15476 12389 15479
rect 11972 15448 12389 15476
rect 11972 15436 11978 15448
rect 12377 15445 12389 15448
rect 12423 15445 12435 15479
rect 12377 15439 12435 15445
rect 23598 15436 23604 15488
rect 23656 15476 23662 15488
rect 24153 15479 24211 15485
rect 24153 15476 24165 15479
rect 23656 15448 24165 15476
rect 23656 15436 23662 15448
rect 24153 15445 24165 15448
rect 24199 15476 24211 15479
rect 24199 15448 25484 15476
rect 24199 15445 24211 15448
rect 24153 15439 24211 15445
rect 12745 15411 12803 15417
rect 12745 15408 12757 15411
rect 11748 15380 12757 15408
rect 11748 15349 11776 15380
rect 12745 15377 12757 15380
rect 12791 15377 12803 15411
rect 12745 15371 12803 15377
rect 17802 15368 17808 15420
rect 17860 15408 17866 15420
rect 18538 15408 18544 15420
rect 17860 15380 18544 15408
rect 17860 15368 17866 15380
rect 18538 15368 18544 15380
rect 18596 15408 18602 15420
rect 18817 15411 18875 15417
rect 18817 15408 18829 15411
rect 18596 15380 18829 15408
rect 18596 15368 18602 15380
rect 18817 15377 18829 15380
rect 18863 15408 18875 15411
rect 18998 15408 19004 15420
rect 18863 15380 19004 15408
rect 18863 15377 18875 15380
rect 18817 15371 18875 15377
rect 18998 15368 19004 15380
rect 19056 15368 19062 15420
rect 20562 15408 20568 15420
rect 20523 15380 20568 15408
rect 20562 15368 20568 15380
rect 20620 15368 20626 15420
rect 23785 15411 23843 15417
rect 23785 15377 23797 15411
rect 23831 15408 23843 15411
rect 25456 15408 25484 15448
rect 26082 15436 26088 15488
rect 26140 15476 26146 15488
rect 26177 15479 26235 15485
rect 26177 15476 26189 15479
rect 26140 15448 26189 15476
rect 26140 15436 26146 15448
rect 26177 15445 26189 15448
rect 26223 15476 26235 15479
rect 26836 15476 26864 15516
rect 27186 15504 27192 15516
rect 27244 15504 27250 15556
rect 28017 15547 28075 15553
rect 28017 15513 28029 15547
rect 28063 15544 28075 15547
rect 28106 15544 28112 15556
rect 28063 15516 28112 15544
rect 28063 15513 28075 15516
rect 28017 15507 28075 15513
rect 28106 15504 28112 15516
rect 28164 15504 28170 15556
rect 28842 15544 28848 15556
rect 28803 15516 28848 15544
rect 28842 15504 28848 15516
rect 28900 15504 28906 15556
rect 26223 15448 26864 15476
rect 26223 15445 26235 15448
rect 26177 15439 26235 15445
rect 26910 15436 26916 15488
rect 26968 15476 26974 15488
rect 28198 15476 28204 15488
rect 26968 15448 28204 15476
rect 26968 15436 26974 15448
rect 28198 15436 28204 15448
rect 28256 15476 28262 15488
rect 28293 15479 28351 15485
rect 28293 15476 28305 15479
rect 28256 15448 28305 15476
rect 28256 15436 28262 15448
rect 28293 15445 28305 15448
rect 28339 15445 28351 15479
rect 28293 15439 28351 15445
rect 25530 15408 25536 15420
rect 23831 15380 24932 15408
rect 23831 15377 23843 15380
rect 23785 15371 23843 15377
rect 24904 15352 24932 15380
rect 25456 15380 25536 15408
rect 11733 15343 11791 15349
rect 11733 15340 11745 15343
rect 11472 15312 11745 15340
rect 8789 15303 8847 15309
rect 11733 15309 11745 15312
rect 11779 15309 11791 15343
rect 11914 15340 11920 15352
rect 11875 15312 11920 15340
rect 11733 15303 11791 15309
rect 6394 15232 6400 15284
rect 6452 15272 6458 15284
rect 7317 15275 7375 15281
rect 7317 15272 7329 15275
rect 6452 15244 7329 15272
rect 6452 15232 6458 15244
rect 7317 15241 7329 15244
rect 7363 15272 7375 15275
rect 7501 15275 7559 15281
rect 7501 15272 7513 15275
rect 7363 15244 7513 15272
rect 7363 15241 7375 15244
rect 7317 15235 7375 15241
rect 7501 15241 7513 15244
rect 7547 15272 7559 15275
rect 7682 15272 7688 15284
rect 7547 15244 7688 15272
rect 7547 15241 7559 15244
rect 7501 15235 7559 15241
rect 7682 15232 7688 15244
rect 7740 15272 7746 15284
rect 8804 15272 8832 15303
rect 11914 15300 11920 15312
rect 11972 15300 11978 15352
rect 18906 15300 18912 15352
rect 18964 15340 18970 15352
rect 19185 15343 19243 15349
rect 19185 15340 19197 15343
rect 18964 15312 19197 15340
rect 18964 15300 18970 15312
rect 19185 15309 19197 15312
rect 19231 15309 19243 15343
rect 19185 15303 19243 15309
rect 24150 15300 24156 15352
rect 24208 15340 24214 15352
rect 24705 15343 24763 15349
rect 24705 15340 24717 15343
rect 24208 15312 24717 15340
rect 24208 15300 24214 15312
rect 24705 15309 24717 15312
rect 24751 15309 24763 15343
rect 24886 15340 24892 15352
rect 24847 15312 24892 15340
rect 24705 15303 24763 15309
rect 24886 15300 24892 15312
rect 24944 15300 24950 15352
rect 25254 15340 25260 15352
rect 25215 15312 25260 15340
rect 25254 15300 25260 15312
rect 25312 15300 25318 15352
rect 25456 15349 25484 15380
rect 25530 15368 25536 15380
rect 25588 15368 25594 15420
rect 26542 15368 26548 15420
rect 26600 15408 26606 15420
rect 27554 15408 27560 15420
rect 26600 15380 27560 15408
rect 26600 15368 26606 15380
rect 27554 15368 27560 15380
rect 27612 15368 27618 15420
rect 27830 15368 27836 15420
rect 27888 15408 27894 15420
rect 28569 15411 28627 15417
rect 28569 15408 28581 15411
rect 27888 15380 28581 15408
rect 27888 15368 27894 15380
rect 28569 15377 28581 15380
rect 28615 15408 28627 15411
rect 29213 15411 29271 15417
rect 29213 15408 29225 15411
rect 28615 15380 29225 15408
rect 28615 15377 28627 15380
rect 28569 15371 28627 15377
rect 29213 15377 29225 15380
rect 29259 15377 29271 15411
rect 29213 15371 29271 15377
rect 25441 15343 25499 15349
rect 25441 15309 25453 15343
rect 25487 15309 25499 15343
rect 25441 15303 25499 15309
rect 25993 15343 26051 15349
rect 25993 15309 26005 15343
rect 26039 15340 26051 15343
rect 27094 15340 27100 15352
rect 26039 15312 27100 15340
rect 26039 15309 26051 15312
rect 25993 15303 26051 15309
rect 27094 15300 27100 15312
rect 27152 15300 27158 15352
rect 27186 15300 27192 15352
rect 27244 15340 27250 15352
rect 27465 15343 27523 15349
rect 27244 15312 27289 15340
rect 27244 15300 27250 15312
rect 27465 15309 27477 15343
rect 27511 15340 27523 15343
rect 27741 15343 27799 15349
rect 27741 15340 27753 15343
rect 27511 15312 27753 15340
rect 27511 15309 27523 15312
rect 27465 15303 27523 15309
rect 27741 15309 27753 15312
rect 27787 15340 27799 15343
rect 28474 15340 28480 15352
rect 27787 15312 28480 15340
rect 27787 15309 27799 15312
rect 27741 15303 27799 15309
rect 7740 15244 8832 15272
rect 11365 15275 11423 15281
rect 7740 15232 7746 15244
rect 11365 15241 11377 15275
rect 11411 15272 11423 15275
rect 12285 15275 12343 15281
rect 12285 15272 12297 15275
rect 11411 15244 12297 15272
rect 11411 15241 11423 15244
rect 11365 15235 11423 15241
rect 12285 15241 12297 15244
rect 12331 15272 12343 15275
rect 13110 15272 13116 15284
rect 12331 15244 13116 15272
rect 12331 15241 12343 15244
rect 12285 15235 12343 15241
rect 13110 15232 13116 15244
rect 13168 15232 13174 15284
rect 14125 15275 14183 15281
rect 14125 15241 14137 15275
rect 14171 15241 14183 15275
rect 14125 15235 14183 15241
rect 14493 15275 14551 15281
rect 14493 15241 14505 15275
rect 14539 15272 14551 15275
rect 14677 15275 14735 15281
rect 14677 15272 14689 15275
rect 14539 15244 14689 15272
rect 14539 15241 14551 15244
rect 14493 15235 14551 15241
rect 14677 15241 14689 15244
rect 14723 15272 14735 15275
rect 14858 15272 14864 15284
rect 14723 15244 14864 15272
rect 14723 15241 14735 15244
rect 14677 15235 14735 15241
rect 5290 15204 5296 15216
rect 5251 15176 5296 15204
rect 5290 15164 5296 15176
rect 5348 15204 5354 15216
rect 5477 15207 5535 15213
rect 5477 15204 5489 15207
rect 5348 15176 5489 15204
rect 5348 15164 5354 15176
rect 5477 15173 5489 15176
rect 5523 15173 5535 15207
rect 14140 15204 14168 15235
rect 14858 15232 14864 15244
rect 14916 15232 14922 15284
rect 18446 15272 18452 15284
rect 18407 15244 18452 15272
rect 18446 15232 18452 15244
rect 18504 15232 18510 15284
rect 21853 15275 21911 15281
rect 21853 15272 21865 15275
rect 20212 15244 21865 15272
rect 20304 15216 20332 15244
rect 21853 15241 21865 15244
rect 21899 15272 21911 15275
rect 22586 15272 22592 15284
rect 21899 15244 22592 15272
rect 21899 15241 21911 15244
rect 21853 15235 21911 15241
rect 22586 15232 22592 15244
rect 22644 15232 22650 15284
rect 14950 15204 14956 15216
rect 14140 15176 14956 15204
rect 5477 15167 5535 15173
rect 14950 15164 14956 15176
rect 15008 15164 15014 15216
rect 15226 15164 15232 15216
rect 15284 15204 15290 15216
rect 15505 15207 15563 15213
rect 15505 15204 15517 15207
rect 15284 15176 15517 15204
rect 15284 15164 15290 15176
rect 15505 15173 15517 15176
rect 15551 15173 15563 15207
rect 15686 15204 15692 15216
rect 15647 15176 15692 15204
rect 15505 15167 15563 15173
rect 15686 15164 15692 15176
rect 15744 15164 15750 15216
rect 18262 15164 18268 15216
rect 18320 15204 18326 15216
rect 18725 15207 18783 15213
rect 18725 15204 18737 15207
rect 18320 15176 18737 15204
rect 18320 15164 18326 15176
rect 18725 15173 18737 15176
rect 18771 15204 18783 15207
rect 20286 15204 20292 15216
rect 18771 15176 20292 15204
rect 18771 15173 18783 15176
rect 18725 15167 18783 15173
rect 20286 15164 20292 15176
rect 20344 15164 20350 15216
rect 22218 15204 22224 15216
rect 22179 15176 22224 15204
rect 22218 15164 22224 15176
rect 22276 15164 22282 15216
rect 24702 15164 24708 15216
rect 24760 15204 24766 15216
rect 25272 15204 25300 15300
rect 24760 15176 25300 15204
rect 24760 15164 24766 15176
rect 26174 15164 26180 15216
rect 26232 15204 26238 15216
rect 26269 15207 26327 15213
rect 26269 15204 26281 15207
rect 26232 15176 26281 15204
rect 26232 15164 26238 15176
rect 26269 15173 26281 15176
rect 26315 15204 26327 15207
rect 27480 15204 27508 15303
rect 28474 15300 28480 15312
rect 28532 15300 28538 15352
rect 28658 15300 28664 15352
rect 28716 15340 28722 15352
rect 29397 15343 29455 15349
rect 29397 15340 29409 15343
rect 28716 15312 29409 15340
rect 28716 15300 28722 15312
rect 29397 15309 29409 15312
rect 29443 15309 29455 15343
rect 29397 15303 29455 15309
rect 27646 15232 27652 15284
rect 27704 15272 27710 15284
rect 28109 15275 28167 15281
rect 28109 15272 28121 15275
rect 27704 15244 28121 15272
rect 27704 15232 27710 15244
rect 28109 15241 28121 15244
rect 28155 15272 28167 15275
rect 28382 15272 28388 15284
rect 28155 15244 28388 15272
rect 28155 15241 28167 15244
rect 28109 15235 28167 15241
rect 28382 15232 28388 15244
rect 28440 15232 28446 15284
rect 26315 15176 27508 15204
rect 26315 15173 26327 15176
rect 26269 15167 26327 15173
rect 400 15114 31680 15136
rect 400 15062 18870 15114
rect 18922 15062 18934 15114
rect 18986 15062 18998 15114
rect 19050 15062 19062 15114
rect 19114 15062 19126 15114
rect 19178 15062 31680 15114
rect 400 15040 31680 15062
rect 785 15003 843 15009
rect 785 14969 797 15003
rect 831 15000 843 15003
rect 1978 15000 1984 15012
rect 831 14972 1984 15000
rect 831 14969 843 14972
rect 785 14963 843 14969
rect 1978 14960 1984 14972
rect 2036 14960 2042 15012
rect 3358 15000 3364 15012
rect 3319 14972 3364 15000
rect 3358 14960 3364 14972
rect 3416 14960 3422 15012
rect 5382 14960 5388 15012
rect 5440 15000 5446 15012
rect 5569 15003 5627 15009
rect 5569 15000 5581 15003
rect 5440 14972 5581 15000
rect 5440 14960 5446 14972
rect 5569 14969 5581 14972
rect 5615 14969 5627 15003
rect 6486 15000 6492 15012
rect 5569 14963 5627 14969
rect 6320 14972 6492 15000
rect 6320 14941 6348 14972
rect 6486 14960 6492 14972
rect 6544 14960 6550 15012
rect 7774 15000 7780 15012
rect 7735 14972 7780 15000
rect 7774 14960 7780 14972
rect 7832 14960 7838 15012
rect 7958 15000 7964 15012
rect 7919 14972 7964 15000
rect 7958 14960 7964 14972
rect 8016 14960 8022 15012
rect 8145 15003 8203 15009
rect 8145 14969 8157 15003
rect 8191 15000 8203 15003
rect 8326 15000 8332 15012
rect 8191 14972 8332 15000
rect 8191 14969 8203 14972
rect 8145 14963 8203 14969
rect 8326 14960 8332 14972
rect 8384 14960 8390 15012
rect 12101 15003 12159 15009
rect 12101 14969 12113 15003
rect 12147 15000 12159 15003
rect 12558 15000 12564 15012
rect 12147 14972 12564 15000
rect 12147 14969 12159 14972
rect 12101 14963 12159 14969
rect 12558 14960 12564 14972
rect 12616 14960 12622 15012
rect 18630 14960 18636 15012
rect 18688 15000 18694 15012
rect 19277 15003 19335 15009
rect 19277 15000 19289 15003
rect 18688 14972 19289 15000
rect 18688 14960 18694 14972
rect 19277 14969 19289 14972
rect 19323 15000 19335 15003
rect 20102 15000 20108 15012
rect 19323 14972 20108 15000
rect 19323 14969 19335 14972
rect 19277 14963 19335 14969
rect 20102 14960 20108 14972
rect 20160 14960 20166 15012
rect 27094 14960 27100 15012
rect 27152 15000 27158 15012
rect 28569 15003 28627 15009
rect 28569 15000 28581 15003
rect 27152 14972 28581 15000
rect 27152 14960 27158 14972
rect 28569 14969 28581 14972
rect 28615 15000 28627 15003
rect 28842 15000 28848 15012
rect 28615 14972 28848 15000
rect 28615 14969 28627 14972
rect 28569 14963 28627 14969
rect 28842 14960 28848 14972
rect 28900 14960 28906 15012
rect 6305 14935 6363 14941
rect 6305 14901 6317 14935
rect 6351 14901 6363 14935
rect 6305 14895 6363 14901
rect 10718 14892 10724 14944
rect 10776 14932 10782 14944
rect 11178 14932 11184 14944
rect 10776 14904 11184 14932
rect 10776 14892 10782 14904
rect 11178 14892 11184 14904
rect 11236 14932 11242 14944
rect 11365 14935 11423 14941
rect 11365 14932 11377 14935
rect 11236 14904 11377 14932
rect 11236 14892 11242 14904
rect 11365 14901 11377 14904
rect 11411 14901 11423 14935
rect 14674 14932 14680 14944
rect 14587 14904 14680 14932
rect 11365 14895 11423 14901
rect 14674 14892 14680 14904
rect 14732 14932 14738 14944
rect 14950 14932 14956 14944
rect 14732 14904 14956 14932
rect 14732 14892 14738 14904
rect 14950 14892 14956 14904
rect 15008 14892 15014 14944
rect 18354 14892 18360 14944
rect 18412 14932 18418 14944
rect 18538 14932 18544 14944
rect 18412 14904 18544 14932
rect 18412 14892 18418 14904
rect 18538 14892 18544 14904
rect 18596 14932 18602 14944
rect 18817 14935 18875 14941
rect 18817 14932 18829 14935
rect 18596 14904 18829 14932
rect 18596 14892 18602 14904
rect 18817 14901 18829 14904
rect 18863 14901 18875 14935
rect 18817 14895 18875 14901
rect 25990 14892 25996 14944
rect 26048 14932 26054 14944
rect 27738 14932 27744 14944
rect 26048 14904 27508 14932
rect 27699 14904 27744 14932
rect 26048 14892 26054 14904
rect 4462 14864 4468 14876
rect 4423 14836 4468 14864
rect 4462 14824 4468 14836
rect 4520 14864 4526 14876
rect 4554 14864 4560 14876
rect 4520 14836 4560 14864
rect 4520 14824 4526 14836
rect 4554 14824 4560 14836
rect 4612 14824 4618 14876
rect 4738 14864 4744 14876
rect 4699 14836 4744 14864
rect 4738 14824 4744 14836
rect 4796 14824 4802 14876
rect 4830 14824 4836 14876
rect 4888 14864 4894 14876
rect 4888 14836 4933 14864
rect 4888 14824 4894 14836
rect 6394 14824 6400 14876
rect 6452 14864 6458 14876
rect 6489 14867 6547 14873
rect 6489 14864 6501 14867
rect 6452 14836 6501 14864
rect 6452 14824 6458 14836
rect 6489 14833 6501 14836
rect 6535 14833 6547 14867
rect 6489 14827 6547 14833
rect 11549 14867 11607 14873
rect 11549 14833 11561 14867
rect 11595 14864 11607 14867
rect 11730 14864 11736 14876
rect 11595 14836 11736 14864
rect 11595 14833 11607 14836
rect 11549 14827 11607 14833
rect 11730 14824 11736 14836
rect 11788 14824 11794 14876
rect 23414 14864 23420 14876
rect 23375 14836 23420 14864
rect 23414 14824 23420 14836
rect 23472 14824 23478 14876
rect 26266 14824 26272 14876
rect 26324 14864 26330 14876
rect 26361 14867 26419 14873
rect 26361 14864 26373 14867
rect 26324 14836 26373 14864
rect 26324 14824 26330 14836
rect 26361 14833 26373 14836
rect 26407 14864 26419 14867
rect 26450 14864 26456 14876
rect 26407 14836 26456 14864
rect 26407 14833 26419 14836
rect 26361 14827 26419 14833
rect 26450 14824 26456 14836
rect 26508 14824 26514 14876
rect 27002 14864 27008 14876
rect 26963 14836 27008 14864
rect 27002 14824 27008 14836
rect 27060 14824 27066 14876
rect 27097 14867 27155 14873
rect 27097 14833 27109 14867
rect 27143 14864 27155 14867
rect 27186 14864 27192 14876
rect 27143 14836 27192 14864
rect 27143 14833 27155 14836
rect 27097 14827 27155 14833
rect 27186 14824 27192 14836
rect 27244 14824 27250 14876
rect 27480 14873 27508 14904
rect 27738 14892 27744 14904
rect 27796 14892 27802 14944
rect 27373 14867 27431 14873
rect 27373 14833 27385 14867
rect 27419 14833 27431 14867
rect 27373 14827 27431 14833
rect 27465 14867 27523 14873
rect 27465 14833 27477 14867
rect 27511 14833 27523 14867
rect 27465 14827 27523 14833
rect 4002 14796 4008 14808
rect 3963 14768 4008 14796
rect 4002 14756 4008 14768
rect 4060 14756 4066 14808
rect 4094 14756 4100 14808
rect 4152 14796 4158 14808
rect 5109 14799 5167 14805
rect 5109 14796 5121 14799
rect 4152 14768 5121 14796
rect 4152 14756 4158 14768
rect 5109 14765 5121 14768
rect 5155 14765 5167 14799
rect 5382 14796 5388 14808
rect 5343 14768 5388 14796
rect 5109 14759 5167 14765
rect 969 14663 1027 14669
rect 969 14629 981 14663
rect 1015 14660 1027 14663
rect 1426 14660 1432 14672
rect 1015 14632 1432 14660
rect 1015 14629 1027 14632
rect 969 14623 1027 14629
rect 1426 14620 1432 14632
rect 1484 14620 1490 14672
rect 5124 14660 5152 14759
rect 5382 14756 5388 14768
rect 5440 14756 5446 14808
rect 11086 14756 11092 14808
rect 11144 14796 11150 14808
rect 11917 14799 11975 14805
rect 11917 14796 11929 14799
rect 11144 14768 11929 14796
rect 11144 14756 11150 14768
rect 11917 14765 11929 14768
rect 11963 14796 11975 14799
rect 14490 14796 14496 14808
rect 11963 14768 14496 14796
rect 11963 14765 11975 14768
rect 11917 14759 11975 14765
rect 14490 14756 14496 14768
rect 14548 14756 14554 14808
rect 23693 14799 23751 14805
rect 23693 14765 23705 14799
rect 23739 14796 23751 14799
rect 24242 14796 24248 14808
rect 23739 14768 24248 14796
rect 23739 14765 23751 14768
rect 23693 14759 23751 14765
rect 24242 14756 24248 14768
rect 24300 14796 24306 14808
rect 26174 14796 26180 14808
rect 24300 14768 26180 14796
rect 24300 14756 24306 14768
rect 26174 14756 26180 14768
rect 26232 14756 26238 14808
rect 10718 14688 10724 14740
rect 10776 14728 10782 14740
rect 10776 14700 14214 14728
rect 10776 14688 10782 14700
rect 6581 14663 6639 14669
rect 6581 14660 6593 14663
rect 5124 14632 6593 14660
rect 6581 14629 6593 14632
rect 6627 14660 6639 14663
rect 6670 14660 6676 14672
rect 6627 14632 6676 14660
rect 6627 14629 6639 14632
rect 6581 14623 6639 14629
rect 6670 14620 6676 14632
rect 6728 14620 6734 14672
rect 14186 14660 14214 14700
rect 26266 14688 26272 14740
rect 26324 14728 26330 14740
rect 27388 14728 27416 14827
rect 26324 14700 27416 14728
rect 26324 14688 26330 14700
rect 14950 14660 14956 14672
rect 14186 14632 14956 14660
rect 14950 14620 14956 14632
rect 15008 14620 15014 14672
rect 19182 14660 19188 14672
rect 19143 14632 19188 14660
rect 19182 14620 19188 14632
rect 19240 14620 19246 14672
rect 24150 14620 24156 14672
rect 24208 14660 24214 14672
rect 24245 14663 24303 14669
rect 24245 14660 24257 14663
rect 24208 14632 24257 14660
rect 24208 14620 24214 14632
rect 24245 14629 24257 14632
rect 24291 14629 24303 14663
rect 24245 14623 24303 14629
rect 400 14570 31680 14592
rect 400 14518 3510 14570
rect 3562 14518 3574 14570
rect 3626 14518 3638 14570
rect 3690 14518 3702 14570
rect 3754 14518 3766 14570
rect 3818 14518 31680 14570
rect 400 14496 31680 14518
rect 4002 14456 4008 14468
rect 3963 14428 4008 14456
rect 4002 14416 4008 14428
rect 4060 14416 4066 14468
rect 4465 14459 4523 14465
rect 4465 14425 4477 14459
rect 4511 14456 4523 14459
rect 4738 14456 4744 14468
rect 4511 14428 4744 14456
rect 4511 14425 4523 14428
rect 4465 14419 4523 14425
rect 4738 14416 4744 14428
rect 4796 14416 4802 14468
rect 6486 14456 6492 14468
rect 6447 14428 6492 14456
rect 6486 14416 6492 14428
rect 6544 14416 6550 14468
rect 6670 14456 6676 14468
rect 6631 14428 6676 14456
rect 6670 14416 6676 14428
rect 6728 14416 6734 14468
rect 11086 14456 11092 14468
rect 11047 14428 11092 14456
rect 11086 14416 11092 14428
rect 11144 14416 11150 14468
rect 11178 14416 11184 14468
rect 11236 14456 11242 14468
rect 11457 14459 11515 14465
rect 11236 14428 11281 14456
rect 11236 14416 11242 14428
rect 11457 14425 11469 14459
rect 11503 14456 11515 14459
rect 11730 14456 11736 14468
rect 11503 14428 11736 14456
rect 11503 14425 11515 14428
rect 11457 14419 11515 14425
rect 11730 14416 11736 14428
rect 11788 14416 11794 14468
rect 12098 14416 12104 14468
rect 12156 14456 12162 14468
rect 12377 14459 12435 14465
rect 12377 14456 12389 14459
rect 12156 14428 12389 14456
rect 12156 14416 12162 14428
rect 12377 14425 12389 14428
rect 12423 14425 12435 14459
rect 12377 14419 12435 14425
rect 14950 14416 14956 14468
rect 15008 14456 15014 14468
rect 15321 14459 15379 14465
rect 15321 14456 15333 14459
rect 15008 14428 15333 14456
rect 15008 14416 15014 14428
rect 15321 14425 15333 14428
rect 15367 14425 15379 14459
rect 15321 14419 15379 14425
rect 15594 14416 15600 14468
rect 15652 14456 15658 14468
rect 16698 14456 16704 14468
rect 15652 14428 16704 14456
rect 15652 14416 15658 14428
rect 16698 14416 16704 14428
rect 16756 14456 16762 14468
rect 17526 14456 17532 14468
rect 16756 14428 17532 14456
rect 16756 14416 16762 14428
rect 17526 14416 17532 14428
rect 17584 14416 17590 14468
rect 18722 14456 18728 14468
rect 18683 14428 18728 14456
rect 18722 14416 18728 14428
rect 18780 14456 18786 14468
rect 19369 14459 19427 14465
rect 19369 14456 19381 14459
rect 18780 14428 19381 14456
rect 18780 14416 18786 14428
rect 19369 14425 19381 14428
rect 19415 14425 19427 14459
rect 26082 14456 26088 14468
rect 26043 14428 26088 14456
rect 19369 14419 19427 14425
rect 26082 14416 26088 14428
rect 26140 14416 26146 14468
rect 26910 14456 26916 14468
rect 26871 14428 26916 14456
rect 26910 14416 26916 14428
rect 26968 14416 26974 14468
rect 27557 14459 27615 14465
rect 27557 14425 27569 14459
rect 27603 14456 27615 14459
rect 28658 14456 28664 14468
rect 27603 14428 28664 14456
rect 27603 14425 27615 14428
rect 27557 14419 27615 14425
rect 3729 14391 3787 14397
rect 3729 14357 3741 14391
rect 3775 14388 3787 14391
rect 4925 14391 4983 14397
rect 4925 14388 4937 14391
rect 3775 14360 4937 14388
rect 3775 14357 3787 14360
rect 3729 14351 3787 14357
rect 4925 14357 4937 14360
rect 4971 14388 4983 14391
rect 5382 14388 5388 14400
rect 4971 14360 5388 14388
rect 4971 14357 4983 14360
rect 4925 14351 4983 14357
rect 5382 14348 5388 14360
rect 5440 14388 5446 14400
rect 5477 14391 5535 14397
rect 5477 14388 5489 14391
rect 5440 14360 5489 14388
rect 5440 14348 5446 14360
rect 5477 14357 5489 14360
rect 5523 14357 5535 14391
rect 15410 14388 15416 14400
rect 5477 14351 5535 14357
rect 14232 14360 15416 14388
rect 1978 14280 1984 14332
rect 2036 14320 2042 14332
rect 2717 14323 2775 14329
rect 2717 14320 2729 14323
rect 2036 14292 2729 14320
rect 2036 14280 2042 14292
rect 2717 14289 2729 14292
rect 2763 14289 2775 14323
rect 2717 14283 2775 14289
rect 3913 14323 3971 14329
rect 3913 14289 3925 14323
rect 3959 14320 3971 14323
rect 4094 14320 4100 14332
rect 3959 14292 4100 14320
rect 3959 14289 3971 14292
rect 3913 14283 3971 14289
rect 4094 14280 4100 14292
rect 4152 14280 4158 14332
rect 4281 14323 4339 14329
rect 4281 14289 4293 14323
rect 4327 14320 4339 14323
rect 4830 14320 4836 14332
rect 4327 14292 4836 14320
rect 4327 14289 4339 14292
rect 4281 14283 4339 14289
rect 4830 14280 4836 14292
rect 4888 14280 4894 14332
rect 5842 14280 5848 14332
rect 5900 14320 5906 14332
rect 12561 14323 12619 14329
rect 12561 14320 12573 14323
rect 5900 14292 7636 14320
rect 5900 14280 5906 14292
rect 690 14252 696 14264
rect 651 14224 696 14252
rect 690 14212 696 14224
rect 748 14212 754 14264
rect 4554 14212 4560 14264
rect 4612 14252 4618 14264
rect 5109 14255 5167 14261
rect 4612 14224 4657 14252
rect 4612 14212 4618 14224
rect 5109 14221 5121 14255
rect 5155 14252 5167 14255
rect 5385 14255 5443 14261
rect 5385 14252 5397 14255
rect 5155 14224 5397 14252
rect 5155 14221 5167 14224
rect 5109 14215 5167 14221
rect 5385 14221 5397 14224
rect 5431 14252 5443 14255
rect 5474 14252 5480 14264
rect 5431 14224 5480 14252
rect 5431 14221 5443 14224
rect 5385 14215 5443 14221
rect 5474 14212 5480 14224
rect 5532 14212 5538 14264
rect 7608 14261 7636 14292
rect 11748 14292 12573 14320
rect 7593 14255 7651 14261
rect 7593 14221 7605 14255
rect 7639 14252 7651 14255
rect 8329 14255 8387 14261
rect 8329 14252 8341 14255
rect 7639 14224 8341 14252
rect 7639 14221 7651 14224
rect 7593 14215 7651 14221
rect 8329 14221 8341 14224
rect 8375 14221 8387 14255
rect 8329 14215 8387 14221
rect 11178 14212 11184 14264
rect 11236 14252 11242 14264
rect 11748 14261 11776 14292
rect 12561 14289 12573 14292
rect 12607 14289 12619 14323
rect 12561 14283 12619 14289
rect 11733 14255 11791 14261
rect 11733 14252 11745 14255
rect 11236 14224 11745 14252
rect 11236 14212 11242 14224
rect 11733 14221 11745 14224
rect 11779 14221 11791 14255
rect 11733 14215 11791 14221
rect 11917 14255 11975 14261
rect 11917 14221 11929 14255
rect 11963 14252 11975 14255
rect 12098 14252 12104 14264
rect 11963 14224 12104 14252
rect 11963 14221 11975 14224
rect 11917 14215 11975 14221
rect 12098 14212 12104 14224
rect 12156 14212 12162 14264
rect 966 14184 972 14196
rect 927 14156 972 14184
rect 966 14144 972 14156
rect 1024 14144 1030 14196
rect 1702 14144 1708 14196
rect 1760 14144 1766 14196
rect 7869 14187 7927 14193
rect 7869 14153 7881 14187
rect 7915 14184 7927 14187
rect 8234 14184 8240 14196
rect 7915 14156 8240 14184
rect 7915 14153 7927 14156
rect 7869 14147 7927 14153
rect 8234 14144 8240 14156
rect 8292 14144 8298 14196
rect 14232 14184 14260 14360
rect 15410 14348 15416 14360
rect 15468 14388 15474 14400
rect 16054 14388 16060 14400
rect 15468 14360 16060 14388
rect 15468 14348 15474 14360
rect 16054 14348 16060 14360
rect 16112 14388 16118 14400
rect 16517 14391 16575 14397
rect 16517 14388 16529 14391
rect 16112 14360 16529 14388
rect 16112 14348 16118 14360
rect 16517 14357 16529 14360
rect 16563 14357 16575 14391
rect 16517 14351 16575 14357
rect 18924 14360 20332 14388
rect 15781 14323 15839 14329
rect 14416 14292 15272 14320
rect 12024 14156 14260 14184
rect 14309 14187 14367 14193
rect 3910 14076 3916 14128
rect 3968 14116 3974 14128
rect 4278 14116 4284 14128
rect 3968 14088 4284 14116
rect 3968 14076 3974 14088
rect 4278 14076 4284 14088
rect 4336 14076 4342 14128
rect 5290 14076 5296 14128
rect 5348 14116 5354 14128
rect 6305 14119 6363 14125
rect 6305 14116 6317 14119
rect 5348 14088 6317 14116
rect 5348 14076 5354 14088
rect 6305 14085 6317 14088
rect 6351 14116 6363 14119
rect 6394 14116 6400 14128
rect 6351 14088 6400 14116
rect 6351 14085 6363 14088
rect 6305 14079 6363 14085
rect 6394 14076 6400 14088
rect 6452 14076 6458 14128
rect 11822 14076 11828 14128
rect 11880 14116 11886 14128
rect 12024 14125 12052 14156
rect 14309 14153 14321 14187
rect 14355 14184 14367 14187
rect 14416 14184 14444 14292
rect 14493 14255 14551 14261
rect 14493 14221 14505 14255
rect 14539 14252 14551 14255
rect 14539 14224 14720 14252
rect 14539 14221 14551 14224
rect 14493 14215 14551 14221
rect 14355 14156 14444 14184
rect 14355 14153 14367 14156
rect 14309 14147 14367 14153
rect 12009 14119 12067 14125
rect 12009 14116 12021 14119
rect 11880 14088 12021 14116
rect 11880 14076 11886 14088
rect 12009 14085 12021 14088
rect 12055 14085 12067 14119
rect 12009 14079 12067 14085
rect 14214 14076 14220 14128
rect 14272 14116 14278 14128
rect 14585 14119 14643 14125
rect 14585 14116 14597 14119
rect 14272 14088 14597 14116
rect 14272 14076 14278 14088
rect 14585 14085 14597 14088
rect 14631 14085 14643 14119
rect 14692 14116 14720 14224
rect 15042 14116 15048 14128
rect 14692 14088 15048 14116
rect 14585 14079 14643 14085
rect 15042 14076 15048 14088
rect 15100 14076 15106 14128
rect 15244 14125 15272 14292
rect 15781 14289 15793 14323
rect 15827 14320 15839 14323
rect 16425 14323 16483 14329
rect 16425 14320 16437 14323
rect 15827 14292 16437 14320
rect 15827 14289 15839 14292
rect 15781 14283 15839 14289
rect 16425 14289 16437 14292
rect 16471 14320 16483 14323
rect 18081 14323 18139 14329
rect 16471 14292 17848 14320
rect 16471 14289 16483 14292
rect 16425 14283 16483 14289
rect 16054 14212 16060 14264
rect 16112 14252 16118 14264
rect 17820 14261 17848 14292
rect 18081 14289 18093 14323
rect 18127 14320 18139 14323
rect 18538 14320 18544 14332
rect 18127 14292 18544 14320
rect 18127 14289 18139 14292
rect 18081 14283 18139 14289
rect 18538 14280 18544 14292
rect 18596 14280 18602 14332
rect 17805 14255 17863 14261
rect 16112 14224 16157 14252
rect 16112 14212 16118 14224
rect 17805 14221 17817 14255
rect 17851 14252 17863 14255
rect 18357 14255 18415 14261
rect 18357 14252 18369 14255
rect 17851 14224 18369 14252
rect 17851 14221 17863 14224
rect 17805 14215 17863 14221
rect 18357 14221 18369 14224
rect 18403 14221 18415 14255
rect 18357 14215 18415 14221
rect 15594 14144 15600 14196
rect 15652 14184 15658 14196
rect 15870 14184 15876 14196
rect 15652 14156 15876 14184
rect 15652 14144 15658 14156
rect 15870 14144 15876 14156
rect 15928 14144 15934 14196
rect 15229 14119 15287 14125
rect 15229 14085 15241 14119
rect 15275 14116 15287 14119
rect 15962 14116 15968 14128
rect 15275 14088 15968 14116
rect 15275 14085 15287 14088
rect 15229 14079 15287 14085
rect 15962 14076 15968 14088
rect 16020 14076 16026 14128
rect 17894 14076 17900 14128
rect 17952 14116 17958 14128
rect 18446 14116 18452 14128
rect 17952 14088 18452 14116
rect 17952 14076 17958 14088
rect 18446 14076 18452 14088
rect 18504 14116 18510 14128
rect 18924 14125 18952 14360
rect 19182 14280 19188 14332
rect 19240 14320 19246 14332
rect 19553 14323 19611 14329
rect 19553 14320 19565 14323
rect 19240 14292 19565 14320
rect 19240 14280 19246 14292
rect 19553 14289 19565 14292
rect 19599 14320 19611 14323
rect 20010 14320 20016 14332
rect 19599 14292 20016 14320
rect 19599 14289 19611 14292
rect 19553 14283 19611 14289
rect 20010 14280 20016 14292
rect 20068 14280 20074 14332
rect 19458 14212 19464 14264
rect 19516 14252 19522 14264
rect 19737 14255 19795 14261
rect 19737 14252 19749 14255
rect 19516 14224 19749 14252
rect 19516 14212 19522 14224
rect 19737 14221 19749 14224
rect 19783 14221 19795 14255
rect 20102 14252 20108 14264
rect 20063 14224 20108 14252
rect 19737 14215 19795 14221
rect 20102 14212 20108 14224
rect 20160 14212 20166 14264
rect 20304 14261 20332 14360
rect 26818 14348 26824 14400
rect 26876 14388 26882 14400
rect 27572 14388 27600 14419
rect 28658 14416 28664 14428
rect 28716 14416 28722 14468
rect 26876 14360 27600 14388
rect 26876 14348 26882 14360
rect 25254 14280 25260 14332
rect 25312 14320 25318 14332
rect 26637 14323 26695 14329
rect 26637 14320 26649 14323
rect 25312 14292 26649 14320
rect 25312 14280 25318 14292
rect 26637 14289 26649 14292
rect 26683 14320 26695 14323
rect 27281 14323 27339 14329
rect 27281 14320 27293 14323
rect 26683 14292 27293 14320
rect 26683 14289 26695 14292
rect 26637 14283 26695 14289
rect 27281 14289 27293 14292
rect 27327 14289 27339 14323
rect 27281 14283 27339 14289
rect 20289 14255 20347 14261
rect 20289 14221 20301 14255
rect 20335 14252 20347 14255
rect 20562 14252 20568 14264
rect 20335 14224 20568 14252
rect 20335 14221 20347 14224
rect 20289 14215 20347 14221
rect 20562 14212 20568 14224
rect 20620 14212 20626 14264
rect 23233 14255 23291 14261
rect 23233 14221 23245 14255
rect 23279 14252 23291 14255
rect 26729 14255 26787 14261
rect 23279 14224 24104 14252
rect 23279 14221 23291 14224
rect 23233 14215 23291 14221
rect 22402 14144 22408 14196
rect 22460 14184 22466 14196
rect 24076 14193 24104 14224
rect 26729 14221 26741 14255
rect 26775 14252 26787 14255
rect 26818 14252 26824 14264
rect 26775 14224 26824 14252
rect 26775 14221 26787 14224
rect 26729 14215 26787 14221
rect 26818 14212 26824 14224
rect 26876 14212 26882 14264
rect 23049 14187 23107 14193
rect 23049 14184 23061 14187
rect 22460 14156 23061 14184
rect 22460 14144 22466 14156
rect 23049 14153 23061 14156
rect 23095 14184 23107 14187
rect 23509 14187 23567 14193
rect 23509 14184 23521 14187
rect 23095 14156 23521 14184
rect 23095 14153 23107 14156
rect 23049 14147 23107 14153
rect 23509 14153 23521 14156
rect 23555 14153 23567 14187
rect 24061 14187 24119 14193
rect 24061 14184 24073 14187
rect 24039 14156 24073 14184
rect 23509 14147 23567 14153
rect 24061 14153 24073 14156
rect 24107 14184 24119 14187
rect 24702 14184 24708 14196
rect 24107 14156 24708 14184
rect 24107 14153 24119 14156
rect 24061 14147 24119 14153
rect 24702 14144 24708 14156
rect 24760 14144 24766 14196
rect 25901 14187 25959 14193
rect 25901 14153 25913 14187
rect 25947 14184 25959 14187
rect 27002 14184 27008 14196
rect 25947 14156 27008 14184
rect 25947 14153 25959 14156
rect 25901 14147 25959 14153
rect 27002 14144 27008 14156
rect 27060 14144 27066 14196
rect 18909 14119 18967 14125
rect 18909 14116 18921 14119
rect 18504 14088 18921 14116
rect 18504 14076 18510 14088
rect 18909 14085 18921 14088
rect 18955 14085 18967 14119
rect 18909 14079 18967 14085
rect 23414 14076 23420 14128
rect 23472 14116 23478 14128
rect 23785 14119 23843 14125
rect 23785 14116 23797 14119
rect 23472 14088 23797 14116
rect 23472 14076 23478 14088
rect 23785 14085 23797 14088
rect 23831 14085 23843 14119
rect 24242 14116 24248 14128
rect 24203 14088 24248 14116
rect 23785 14079 23843 14085
rect 24242 14076 24248 14088
rect 24300 14076 24306 14128
rect 25990 14076 25996 14128
rect 26048 14116 26054 14128
rect 26177 14119 26235 14125
rect 26177 14116 26189 14119
rect 26048 14088 26189 14116
rect 26048 14076 26054 14088
rect 26177 14085 26189 14088
rect 26223 14085 26235 14119
rect 26177 14079 26235 14085
rect 26266 14076 26272 14128
rect 26324 14116 26330 14128
rect 26361 14119 26419 14125
rect 26361 14116 26373 14119
rect 26324 14088 26373 14116
rect 26324 14076 26330 14088
rect 26361 14085 26373 14088
rect 26407 14085 26419 14119
rect 26361 14079 26419 14085
rect 28842 14076 28848 14128
rect 28900 14116 28906 14128
rect 29394 14116 29400 14128
rect 28900 14088 29400 14116
rect 28900 14076 28906 14088
rect 29394 14076 29400 14088
rect 29452 14076 29458 14128
rect 400 14026 31680 14048
rect 400 13974 18870 14026
rect 18922 13974 18934 14026
rect 18986 13974 18998 14026
rect 19050 13974 19062 14026
rect 19114 13974 19126 14026
rect 19178 13974 31680 14026
rect 400 13952 31680 13974
rect 785 13915 843 13921
rect 785 13881 797 13915
rect 831 13912 843 13915
rect 966 13912 972 13924
rect 831 13884 972 13912
rect 831 13881 843 13884
rect 785 13875 843 13881
rect 966 13872 972 13884
rect 1024 13872 1030 13924
rect 2622 13872 2628 13924
rect 2680 13912 2686 13924
rect 14674 13912 14680 13924
rect 2680 13884 14214 13912
rect 14635 13884 14680 13912
rect 2680 13872 2686 13884
rect 4094 13804 4100 13856
rect 4152 13804 4158 13856
rect 11822 13844 11828 13856
rect 11783 13816 11828 13844
rect 11822 13804 11828 13816
rect 11880 13804 11886 13856
rect 14186 13844 14214 13884
rect 14674 13872 14680 13884
rect 14732 13872 14738 13924
rect 18262 13912 18268 13924
rect 16072 13884 18268 13912
rect 16072 13856 16100 13884
rect 18262 13872 18268 13884
rect 18320 13872 18326 13924
rect 19737 13915 19795 13921
rect 19737 13881 19749 13915
rect 19783 13912 19795 13915
rect 20102 13912 20108 13924
rect 19783 13884 20108 13912
rect 19783 13881 19795 13884
rect 19737 13875 19795 13881
rect 20102 13872 20108 13884
rect 20160 13912 20166 13924
rect 21022 13912 21028 13924
rect 20160 13884 21028 13912
rect 20160 13872 20166 13884
rect 21022 13872 21028 13884
rect 21080 13872 21086 13924
rect 21666 13912 21672 13924
rect 21579 13884 21672 13912
rect 21666 13872 21672 13884
rect 21724 13912 21730 13924
rect 22218 13912 22224 13924
rect 21724 13884 22224 13912
rect 21724 13872 21730 13884
rect 22218 13872 22224 13884
rect 22276 13872 22282 13924
rect 24794 13912 24800 13924
rect 24755 13884 24800 13912
rect 24794 13872 24800 13884
rect 24852 13872 24858 13924
rect 26358 13872 26364 13924
rect 26416 13912 26422 13924
rect 26453 13915 26511 13921
rect 26453 13912 26465 13915
rect 26416 13884 26465 13912
rect 26416 13872 26422 13884
rect 26453 13881 26465 13884
rect 26499 13881 26511 13915
rect 26453 13875 26511 13881
rect 26729 13915 26787 13921
rect 26729 13881 26741 13915
rect 26775 13912 26787 13915
rect 26910 13912 26916 13924
rect 26775 13884 26916 13912
rect 26775 13881 26787 13884
rect 26729 13875 26787 13881
rect 26910 13872 26916 13884
rect 26968 13872 26974 13924
rect 15134 13844 15140 13856
rect 14186 13816 15140 13844
rect 15134 13804 15140 13816
rect 15192 13804 15198 13856
rect 15229 13847 15287 13853
rect 15229 13813 15241 13847
rect 15275 13844 15287 13847
rect 15318 13844 15324 13856
rect 15275 13816 15324 13844
rect 15275 13813 15287 13816
rect 15229 13807 15287 13813
rect 15318 13804 15324 13816
rect 15376 13844 15382 13856
rect 15597 13847 15655 13853
rect 15597 13844 15609 13847
rect 15376 13816 15609 13844
rect 15376 13804 15382 13816
rect 15597 13813 15609 13816
rect 15643 13813 15655 13847
rect 15597 13807 15655 13813
rect 16054 13804 16060 13856
rect 16112 13804 16118 13856
rect 19185 13847 19243 13853
rect 19185 13813 19197 13847
rect 19231 13844 19243 13847
rect 19366 13844 19372 13856
rect 19231 13816 19372 13844
rect 19231 13813 19243 13816
rect 19185 13807 19243 13813
rect 19366 13804 19372 13816
rect 19424 13804 19430 13856
rect 29118 13804 29124 13856
rect 29176 13804 29182 13856
rect 12834 13776 12840 13788
rect 12795 13748 12840 13776
rect 12834 13736 12840 13748
rect 12892 13736 12898 13788
rect 13021 13779 13079 13785
rect 13021 13745 13033 13779
rect 13067 13776 13079 13779
rect 13110 13776 13116 13788
rect 13067 13748 13116 13776
rect 13067 13745 13079 13748
rect 13021 13739 13079 13745
rect 13110 13736 13116 13748
rect 13168 13776 13174 13788
rect 15042 13776 15048 13788
rect 13168 13748 15048 13776
rect 13168 13736 13174 13748
rect 15042 13736 15048 13748
rect 15100 13736 15106 13788
rect 18630 13776 18636 13788
rect 18591 13748 18636 13776
rect 18630 13736 18636 13748
rect 18688 13736 18694 13788
rect 18722 13736 18728 13788
rect 18780 13776 18786 13788
rect 18780 13748 18825 13776
rect 18780 13736 18786 13748
rect 20010 13736 20016 13788
rect 20068 13776 20074 13788
rect 22037 13779 22095 13785
rect 22037 13776 22049 13779
rect 20068 13748 22049 13776
rect 20068 13736 20074 13748
rect 22037 13745 22049 13748
rect 22083 13776 22095 13779
rect 22126 13776 22132 13788
rect 22083 13748 22132 13776
rect 22083 13745 22095 13748
rect 22037 13739 22095 13745
rect 22126 13736 22132 13748
rect 22184 13736 22190 13788
rect 22402 13776 22408 13788
rect 22363 13748 22408 13776
rect 22402 13736 22408 13748
rect 22460 13736 22466 13788
rect 23414 13776 23420 13788
rect 23375 13748 23420 13776
rect 23414 13736 23420 13748
rect 23472 13736 23478 13788
rect 25806 13776 25812 13788
rect 25767 13748 25812 13776
rect 25806 13736 25812 13748
rect 25864 13736 25870 13788
rect 25898 13736 25904 13788
rect 25956 13776 25962 13788
rect 25956 13748 26001 13776
rect 25956 13736 25962 13748
rect 3358 13708 3364 13720
rect 3319 13680 3364 13708
rect 3358 13668 3364 13680
rect 3416 13668 3422 13720
rect 3637 13711 3695 13717
rect 3637 13677 3649 13711
rect 3683 13708 3695 13711
rect 4002 13708 4008 13720
rect 3683 13680 4008 13708
rect 3683 13677 3695 13680
rect 3637 13671 3695 13677
rect 4002 13668 4008 13680
rect 4060 13668 4066 13720
rect 5382 13708 5388 13720
rect 5343 13680 5388 13708
rect 5382 13668 5388 13680
rect 5440 13668 5446 13720
rect 14398 13668 14404 13720
rect 14456 13708 14462 13720
rect 14858 13708 14864 13720
rect 14456 13680 14864 13708
rect 14456 13668 14462 13680
rect 14858 13668 14864 13680
rect 14916 13708 14922 13720
rect 15321 13711 15379 13717
rect 15321 13708 15333 13711
rect 14916 13680 15333 13708
rect 14916 13668 14922 13680
rect 15321 13677 15333 13680
rect 15367 13708 15379 13711
rect 16330 13708 16336 13720
rect 15367 13680 16336 13708
rect 15367 13677 15379 13680
rect 15321 13671 15379 13677
rect 16330 13668 16336 13680
rect 16388 13668 16394 13720
rect 17342 13708 17348 13720
rect 17303 13680 17348 13708
rect 17342 13668 17348 13680
rect 17400 13668 17406 13720
rect 21850 13708 21856 13720
rect 21811 13680 21856 13708
rect 21850 13668 21856 13680
rect 21908 13668 21914 13720
rect 22310 13708 22316 13720
rect 22271 13680 22316 13708
rect 22310 13668 22316 13680
rect 22368 13668 22374 13720
rect 23693 13711 23751 13717
rect 23693 13677 23705 13711
rect 23739 13708 23751 13711
rect 24150 13708 24156 13720
rect 23739 13680 24156 13708
rect 23739 13677 23751 13680
rect 23693 13671 23751 13677
rect 24150 13668 24156 13680
rect 24208 13668 24214 13720
rect 28382 13708 28388 13720
rect 28343 13680 28388 13708
rect 28382 13668 28388 13680
rect 28440 13668 28446 13720
rect 28750 13708 28756 13720
rect 28711 13680 28756 13708
rect 28750 13668 28756 13680
rect 28808 13668 28814 13720
rect 29026 13668 29032 13720
rect 29084 13708 29090 13720
rect 30133 13711 30191 13717
rect 30133 13708 30145 13711
rect 29084 13680 30145 13708
rect 29084 13668 29090 13680
rect 30133 13677 30145 13680
rect 30179 13677 30191 13711
rect 30133 13671 30191 13677
rect 12374 13600 12380 13652
rect 12432 13640 12438 13652
rect 12432 13612 13156 13640
rect 12432 13600 12438 13612
rect 690 13532 696 13584
rect 748 13572 754 13584
rect 966 13572 972 13584
rect 748 13544 972 13572
rect 748 13532 754 13544
rect 966 13532 972 13544
rect 1024 13532 1030 13584
rect 12009 13575 12067 13581
rect 12009 13541 12021 13575
rect 12055 13572 12067 13575
rect 12742 13572 12748 13584
rect 12055 13544 12748 13572
rect 12055 13541 12067 13544
rect 12009 13535 12067 13541
rect 12742 13532 12748 13544
rect 12800 13532 12806 13584
rect 13128 13581 13156 13612
rect 24702 13600 24708 13652
rect 24760 13640 24766 13652
rect 24760 13612 26128 13640
rect 24760 13600 24766 13612
rect 13113 13575 13171 13581
rect 13113 13541 13125 13575
rect 13159 13572 13171 13575
rect 13386 13572 13392 13584
rect 13159 13544 13392 13572
rect 13159 13541 13171 13544
rect 13113 13535 13171 13541
rect 13386 13532 13392 13544
rect 13444 13532 13450 13584
rect 18446 13572 18452 13584
rect 18359 13544 18452 13572
rect 18446 13532 18452 13544
rect 18504 13572 18510 13584
rect 19277 13575 19335 13581
rect 19277 13572 19289 13575
rect 18504 13544 19289 13572
rect 18504 13532 18510 13544
rect 19277 13541 19289 13544
rect 19323 13572 19335 13575
rect 19550 13572 19556 13584
rect 19323 13544 19556 13572
rect 19323 13541 19335 13544
rect 19277 13535 19335 13541
rect 19550 13532 19556 13544
rect 19608 13572 19614 13584
rect 19734 13572 19740 13584
rect 19608 13544 19740 13572
rect 19608 13532 19614 13544
rect 19734 13532 19740 13544
rect 19792 13532 19798 13584
rect 24613 13575 24671 13581
rect 24613 13541 24625 13575
rect 24659 13572 24671 13575
rect 25530 13572 25536 13584
rect 24659 13544 25536 13572
rect 24659 13541 24671 13544
rect 24613 13535 24671 13541
rect 25530 13532 25536 13544
rect 25588 13532 25594 13584
rect 26100 13581 26128 13612
rect 26085 13575 26143 13581
rect 26085 13541 26097 13575
rect 26131 13572 26143 13575
rect 26174 13572 26180 13584
rect 26131 13544 26180 13572
rect 26131 13541 26143 13544
rect 26085 13535 26143 13541
rect 26174 13532 26180 13544
rect 26232 13532 26238 13584
rect 400 13482 31680 13504
rect 400 13430 3510 13482
rect 3562 13430 3574 13482
rect 3626 13430 3638 13482
rect 3690 13430 3702 13482
rect 3754 13430 3766 13482
rect 3818 13430 31680 13482
rect 400 13408 31680 13430
rect 3637 13371 3695 13377
rect 3637 13337 3649 13371
rect 3683 13368 3695 13371
rect 4002 13368 4008 13380
rect 3683 13340 4008 13368
rect 3683 13337 3695 13340
rect 3637 13331 3695 13337
rect 4002 13328 4008 13340
rect 4060 13328 4066 13380
rect 13110 13368 13116 13380
rect 13071 13340 13116 13368
rect 13110 13328 13116 13340
rect 13168 13328 13174 13380
rect 13386 13368 13392 13380
rect 13347 13340 13392 13368
rect 13386 13328 13392 13340
rect 13444 13328 13450 13380
rect 14677 13371 14735 13377
rect 14677 13337 14689 13371
rect 14723 13368 14735 13371
rect 15318 13368 15324 13380
rect 14723 13340 15324 13368
rect 14723 13337 14735 13340
rect 14677 13331 14735 13337
rect 15318 13328 15324 13340
rect 15376 13368 15382 13380
rect 15413 13371 15471 13377
rect 15413 13368 15425 13371
rect 15376 13340 15425 13368
rect 15376 13328 15382 13340
rect 15413 13337 15425 13340
rect 15459 13337 15471 13371
rect 15413 13331 15471 13337
rect 16330 13328 16336 13380
rect 16388 13368 16394 13380
rect 16517 13371 16575 13377
rect 16517 13368 16529 13371
rect 16388 13340 16529 13368
rect 16388 13328 16394 13340
rect 16517 13337 16529 13340
rect 16563 13337 16575 13371
rect 18446 13368 18452 13380
rect 18407 13340 18452 13368
rect 16517 13331 16575 13337
rect 18446 13328 18452 13340
rect 18504 13328 18510 13380
rect 18630 13368 18636 13380
rect 18591 13340 18636 13368
rect 18630 13328 18636 13340
rect 18688 13328 18694 13380
rect 19093 13371 19151 13377
rect 19093 13337 19105 13371
rect 19139 13368 19151 13371
rect 19366 13368 19372 13380
rect 19139 13340 19372 13368
rect 19139 13337 19151 13340
rect 19093 13331 19151 13337
rect 19366 13328 19372 13340
rect 19424 13328 19430 13380
rect 20102 13368 20108 13380
rect 20063 13340 20108 13368
rect 20102 13328 20108 13340
rect 20160 13328 20166 13380
rect 21666 13368 21672 13380
rect 21627 13340 21672 13368
rect 21666 13328 21672 13340
rect 21724 13328 21730 13380
rect 22126 13368 22132 13380
rect 22087 13340 22132 13368
rect 22126 13328 22132 13340
rect 22184 13328 22190 13380
rect 23414 13328 23420 13380
rect 23472 13368 23478 13380
rect 23509 13371 23567 13377
rect 23509 13368 23521 13371
rect 23472 13340 23521 13368
rect 23472 13328 23478 13340
rect 23509 13337 23521 13340
rect 23555 13337 23567 13371
rect 24242 13368 24248 13380
rect 24203 13340 24248 13368
rect 23509 13331 23567 13337
rect 24242 13328 24248 13340
rect 24300 13328 24306 13380
rect 24794 13368 24800 13380
rect 24755 13340 24800 13368
rect 24794 13328 24800 13340
rect 24852 13328 24858 13380
rect 25806 13368 25812 13380
rect 25767 13340 25812 13368
rect 25806 13328 25812 13340
rect 25864 13328 25870 13380
rect 26174 13368 26180 13380
rect 26135 13340 26180 13368
rect 26174 13328 26180 13340
rect 26232 13328 26238 13380
rect 28750 13328 28756 13380
rect 28808 13368 28814 13380
rect 28937 13371 28995 13377
rect 28937 13368 28949 13371
rect 28808 13340 28949 13368
rect 28808 13328 28814 13340
rect 28937 13337 28949 13340
rect 28983 13368 28995 13371
rect 29302 13368 29308 13380
rect 28983 13340 29308 13368
rect 28983 13337 28995 13340
rect 28937 13331 28995 13337
rect 29302 13328 29308 13340
rect 29360 13328 29366 13380
rect 3358 13260 3364 13312
rect 3416 13300 3422 13312
rect 3910 13300 3916 13312
rect 3416 13272 3916 13300
rect 3416 13260 3422 13272
rect 3910 13260 3916 13272
rect 3968 13260 3974 13312
rect 12282 13260 12288 13312
rect 12340 13300 12346 13312
rect 12340 13272 12512 13300
rect 12340 13260 12346 13272
rect 3453 13235 3511 13241
rect 3453 13201 3465 13235
rect 3499 13232 3511 13235
rect 5382 13232 5388 13244
rect 3499 13204 5388 13232
rect 3499 13201 3511 13204
rect 3453 13195 3511 13201
rect 5382 13192 5388 13204
rect 5440 13192 5446 13244
rect 12484 13241 12512 13272
rect 12834 13260 12840 13312
rect 12892 13300 12898 13312
rect 13205 13303 13263 13309
rect 13205 13300 13217 13303
rect 12892 13272 13217 13300
rect 12892 13260 12898 13272
rect 13205 13269 13217 13272
rect 13251 13269 13263 13303
rect 13205 13263 13263 13269
rect 14953 13303 15011 13309
rect 14953 13269 14965 13303
rect 14999 13300 15011 13303
rect 16054 13300 16060 13312
rect 14999 13272 16060 13300
rect 14999 13269 15011 13272
rect 14953 13263 15011 13269
rect 11181 13235 11239 13241
rect 11181 13201 11193 13235
rect 11227 13232 11239 13235
rect 12469 13235 12527 13241
rect 11227 13204 12420 13232
rect 11227 13201 11239 13204
rect 11181 13195 11239 13201
rect 12392 13176 12420 13204
rect 12469 13201 12481 13235
rect 12515 13201 12527 13235
rect 12469 13195 12527 13201
rect 3910 13124 3916 13176
rect 3968 13164 3974 13176
rect 8786 13164 8792 13176
rect 3968 13136 8792 13164
rect 3968 13124 3974 13136
rect 8786 13124 8792 13136
rect 8844 13124 8850 13176
rect 12374 13164 12380 13176
rect 12287 13136 12380 13164
rect 12374 13124 12380 13136
rect 12432 13124 12438 13176
rect 12742 13164 12748 13176
rect 12703 13136 12748 13164
rect 12742 13124 12748 13136
rect 12800 13124 12806 13176
rect 12834 13124 12840 13176
rect 12892 13164 12898 13176
rect 12892 13136 12937 13164
rect 12892 13124 12898 13136
rect 3821 13099 3879 13105
rect 3821 13065 3833 13099
rect 3867 13096 3879 13099
rect 4094 13096 4100 13108
rect 3867 13068 4100 13096
rect 3867 13065 3879 13068
rect 3821 13059 3879 13065
rect 4094 13056 4100 13068
rect 4152 13056 4158 13108
rect 10810 13056 10816 13108
rect 10868 13096 10874 13108
rect 11365 13099 11423 13105
rect 11365 13096 11377 13099
rect 10868 13068 11377 13096
rect 10868 13056 10874 13068
rect 11365 13065 11377 13068
rect 11411 13096 11423 13099
rect 11733 13099 11791 13105
rect 11733 13096 11745 13099
rect 11411 13068 11745 13096
rect 11411 13065 11423 13068
rect 11365 13059 11423 13065
rect 11733 13065 11745 13068
rect 11779 13065 11791 13099
rect 13220 13096 13248 13263
rect 16054 13260 16060 13272
rect 16112 13260 16118 13312
rect 16422 13260 16428 13312
rect 16480 13300 16486 13312
rect 18722 13300 18728 13312
rect 16480 13272 18728 13300
rect 16480 13260 16486 13272
rect 18722 13260 18728 13272
rect 18780 13300 18786 13312
rect 18817 13303 18875 13309
rect 18817 13300 18829 13303
rect 18780 13272 18829 13300
rect 18780 13260 18786 13272
rect 18817 13269 18829 13272
rect 18863 13269 18875 13303
rect 18817 13263 18875 13269
rect 19277 13303 19335 13309
rect 19277 13269 19289 13303
rect 19323 13300 19335 13303
rect 21485 13303 21543 13309
rect 19323 13272 19872 13300
rect 19323 13269 19335 13272
rect 19277 13263 19335 13269
rect 19384 13244 19412 13272
rect 14861 13235 14919 13241
rect 14861 13201 14873 13235
rect 14907 13232 14919 13235
rect 16606 13232 16612 13244
rect 14907 13204 16612 13232
rect 14907 13201 14919 13204
rect 14861 13195 14919 13201
rect 13849 13167 13907 13173
rect 13849 13133 13861 13167
rect 13895 13164 13907 13167
rect 14214 13164 14220 13176
rect 13895 13136 14220 13164
rect 13895 13133 13907 13136
rect 13849 13127 13907 13133
rect 14214 13124 14220 13136
rect 14272 13164 14278 13176
rect 15597 13167 15655 13173
rect 15597 13164 15609 13167
rect 14272 13136 14317 13164
rect 14876 13136 15609 13164
rect 14272 13124 14278 13136
rect 14306 13096 14312 13108
rect 13220 13068 14312 13096
rect 11733 13059 11791 13065
rect 14306 13056 14312 13068
rect 14364 13096 14370 13108
rect 14674 13096 14680 13108
rect 14364 13068 14680 13096
rect 14364 13056 14370 13068
rect 14674 13056 14680 13068
rect 14732 13056 14738 13108
rect 14876 13040 14904 13136
rect 15597 13133 15609 13136
rect 15643 13133 15655 13167
rect 15778 13164 15784 13176
rect 15739 13136 15784 13164
rect 15597 13127 15655 13133
rect 15778 13124 15784 13136
rect 15836 13124 15842 13176
rect 16146 13164 16152 13176
rect 16107 13136 16152 13164
rect 16146 13124 16152 13136
rect 16204 13124 16210 13176
rect 16348 13173 16376 13204
rect 16606 13192 16612 13204
rect 16664 13232 16670 13244
rect 17250 13232 17256 13244
rect 16664 13204 17256 13232
rect 16664 13192 16670 13204
rect 17250 13192 17256 13204
rect 17308 13192 17314 13244
rect 19366 13192 19372 13244
rect 19424 13192 19430 13244
rect 16333 13167 16391 13173
rect 16333 13133 16345 13167
rect 16379 13133 16391 13167
rect 17526 13164 17532 13176
rect 17487 13136 17532 13164
rect 16333 13127 16391 13133
rect 17526 13124 17532 13136
rect 17584 13164 17590 13176
rect 17989 13167 18047 13173
rect 17989 13164 18001 13167
rect 17584 13136 18001 13164
rect 17584 13124 17590 13136
rect 17989 13133 18001 13136
rect 18035 13133 18047 13167
rect 19734 13164 19740 13176
rect 19695 13136 19740 13164
rect 17989 13127 18047 13133
rect 19734 13124 19740 13136
rect 19792 13124 19798 13176
rect 19844 13164 19872 13272
rect 21485 13269 21497 13303
rect 21531 13300 21543 13303
rect 22310 13300 22316 13312
rect 21531 13272 22316 13300
rect 21531 13269 21543 13272
rect 21485 13263 21543 13269
rect 22310 13260 22316 13272
rect 22368 13260 22374 13312
rect 23141 13235 23199 13241
rect 23141 13232 23153 13235
rect 22512 13204 23153 13232
rect 19921 13167 19979 13173
rect 19921 13164 19933 13167
rect 19844 13136 19933 13164
rect 19921 13133 19933 13136
rect 19967 13133 19979 13167
rect 19921 13127 19979 13133
rect 20746 13124 20752 13176
rect 20804 13164 20810 13176
rect 21850 13164 21856 13176
rect 20804 13136 21856 13164
rect 20804 13124 20810 13136
rect 21850 13124 21856 13136
rect 21908 13164 21914 13176
rect 22512 13173 22540 13204
rect 23141 13201 23153 13204
rect 23187 13201 23199 13235
rect 24260 13232 24288 13328
rect 25824 13300 25852 13328
rect 26542 13300 26548 13312
rect 25824 13272 26548 13300
rect 26542 13260 26548 13272
rect 26600 13260 26606 13312
rect 24260 13204 25208 13232
rect 23141 13195 23199 13201
rect 21945 13167 22003 13173
rect 21945 13164 21957 13167
rect 21908 13136 21957 13164
rect 21908 13124 21914 13136
rect 21945 13133 21957 13136
rect 21991 13164 22003 13167
rect 22497 13167 22555 13173
rect 22497 13164 22509 13167
rect 21991 13136 22509 13164
rect 21991 13133 22003 13136
rect 21945 13127 22003 13133
rect 22497 13133 22509 13136
rect 22543 13133 22555 13167
rect 22497 13127 22555 13133
rect 22773 13167 22831 13173
rect 22773 13133 22785 13167
rect 22819 13164 22831 13167
rect 22957 13167 23015 13173
rect 22957 13164 22969 13167
rect 22819 13136 22969 13164
rect 22819 13133 22831 13136
rect 22773 13127 22831 13133
rect 22957 13133 22969 13136
rect 23003 13164 23015 13167
rect 23693 13167 23751 13173
rect 23693 13164 23705 13167
rect 23003 13136 23705 13164
rect 23003 13133 23015 13136
rect 22957 13127 23015 13133
rect 23693 13133 23705 13136
rect 23739 13164 23751 13167
rect 24150 13164 24156 13176
rect 23739 13136 24156 13164
rect 23739 13133 23751 13136
rect 23693 13127 23751 13133
rect 24150 13124 24156 13136
rect 24208 13124 24214 13176
rect 25180 13173 25208 13204
rect 24981 13167 25039 13173
rect 24981 13133 24993 13167
rect 25027 13133 25039 13167
rect 24981 13127 25039 13133
rect 25165 13167 25223 13173
rect 25165 13133 25177 13167
rect 25211 13133 25223 13167
rect 25530 13164 25536 13176
rect 25491 13136 25536 13164
rect 25165 13127 25223 13133
rect 15042 13056 15048 13108
rect 15100 13096 15106 13108
rect 17345 13099 17403 13105
rect 17345 13096 17357 13099
rect 15100 13068 17357 13096
rect 15100 13056 15106 13068
rect 17345 13065 17357 13068
rect 17391 13096 17403 13099
rect 18173 13099 18231 13105
rect 18173 13096 18185 13099
rect 17391 13068 18185 13096
rect 17391 13065 17403 13068
rect 17345 13059 17403 13065
rect 18173 13065 18185 13068
rect 18219 13065 18231 13099
rect 19829 13099 19887 13105
rect 19829 13096 19841 13099
rect 18173 13059 18231 13065
rect 19476 13068 19841 13096
rect 19476 13040 19504 13068
rect 19829 13065 19841 13068
rect 19875 13065 19887 13099
rect 22402 13096 22408 13108
rect 19829 13059 19887 13065
rect 21776 13068 22408 13096
rect 9246 12988 9252 13040
rect 9304 13028 9310 13040
rect 9890 13028 9896 13040
rect 9304 13000 9896 13028
rect 9304 12988 9310 13000
rect 9890 12988 9896 13000
rect 9948 12988 9954 13040
rect 11454 13028 11460 13040
rect 11415 13000 11460 13028
rect 11454 12988 11460 13000
rect 11512 12988 11518 13040
rect 13665 13031 13723 13037
rect 13665 12997 13677 13031
rect 13711 13028 13723 13031
rect 14030 13028 14036 13040
rect 13711 13000 14036 13028
rect 13711 12997 13723 13000
rect 13665 12991 13723 12997
rect 14030 12988 14036 13000
rect 14088 12988 14094 13040
rect 14493 13031 14551 13037
rect 14493 12997 14505 13031
rect 14539 13028 14551 13031
rect 14858 13028 14864 13040
rect 14539 13000 14864 13028
rect 14539 12997 14551 13000
rect 14493 12991 14551 12997
rect 14858 12988 14864 13000
rect 14916 12988 14922 13040
rect 17161 13031 17219 13037
rect 17161 12997 17173 13031
rect 17207 13028 17219 13031
rect 17618 13028 17624 13040
rect 17207 13000 17624 13028
rect 17207 12997 17219 13000
rect 17161 12991 17219 12997
rect 17618 12988 17624 13000
rect 17676 12988 17682 13040
rect 19458 13028 19464 13040
rect 19419 13000 19464 13028
rect 19458 12988 19464 13000
rect 19516 12988 19522 13040
rect 19734 12988 19740 13040
rect 19792 13028 19798 13040
rect 20473 13031 20531 13037
rect 20473 13028 20485 13031
rect 19792 13000 20485 13028
rect 19792 12988 19798 13000
rect 20473 12997 20485 13000
rect 20519 12997 20531 13031
rect 20473 12991 20531 12997
rect 21666 12988 21672 13040
rect 21724 13028 21730 13040
rect 21776 13037 21804 13068
rect 22402 13056 22408 13068
rect 22460 13056 22466 13108
rect 24996 13096 25024 13127
rect 25530 13124 25536 13136
rect 25588 13124 25594 13176
rect 25717 13167 25775 13173
rect 25717 13133 25729 13167
rect 25763 13133 25775 13167
rect 25717 13127 25775 13133
rect 23984 13068 25024 13096
rect 25732 13096 25760 13127
rect 25806 13124 25812 13176
rect 25864 13164 25870 13176
rect 27370 13164 27376 13176
rect 25864 13136 27376 13164
rect 25864 13124 25870 13136
rect 27370 13124 27376 13136
rect 27428 13124 27434 13176
rect 25898 13096 25904 13108
rect 25732 13068 25904 13096
rect 23984 13040 24012 13068
rect 21761 13031 21819 13037
rect 21761 13028 21773 13031
rect 21724 13000 21773 13028
rect 21724 12988 21730 13000
rect 21761 12997 21773 13000
rect 21807 12997 21819 13031
rect 23966 13028 23972 13040
rect 23927 13000 23972 13028
rect 21761 12991 21819 12997
rect 23966 12988 23972 13000
rect 24024 12988 24030 13040
rect 24429 13031 24487 13037
rect 24429 12997 24441 13031
rect 24475 13028 24487 13031
rect 25732 13028 25760 13068
rect 25898 13056 25904 13068
rect 25956 13096 25962 13108
rect 25956 13068 26128 13096
rect 25956 13056 25962 13068
rect 26100 13037 26128 13068
rect 28382 13056 28388 13108
rect 28440 13096 28446 13108
rect 29121 13099 29179 13105
rect 29121 13096 29133 13099
rect 28440 13068 29133 13096
rect 28440 13056 28446 13068
rect 29121 13065 29133 13068
rect 29167 13065 29179 13099
rect 29121 13059 29179 13065
rect 24475 13000 25760 13028
rect 26085 13031 26143 13037
rect 24475 12997 24487 13000
rect 24429 12991 24487 12997
rect 26085 12997 26097 13031
rect 26131 13028 26143 13031
rect 26726 13028 26732 13040
rect 26131 13000 26732 13028
rect 26131 12997 26143 13000
rect 26085 12991 26143 12997
rect 26726 12988 26732 13000
rect 26784 12988 26790 13040
rect 28566 13028 28572 13040
rect 28527 13000 28572 13028
rect 28566 12988 28572 13000
rect 28624 12988 28630 13040
rect 28845 13031 28903 13037
rect 28845 12997 28857 13031
rect 28891 13028 28903 13031
rect 29026 13028 29032 13040
rect 28891 13000 29032 13028
rect 28891 12997 28903 13000
rect 28845 12991 28903 12997
rect 29026 12988 29032 13000
rect 29084 12988 29090 13040
rect 400 12938 31680 12960
rect 400 12886 18870 12938
rect 18922 12886 18934 12938
rect 18986 12886 18998 12938
rect 19050 12886 19062 12938
rect 19114 12886 19126 12938
rect 19178 12886 31680 12938
rect 400 12864 31680 12886
rect 14950 12824 14956 12836
rect 4526 12796 14956 12824
rect 1150 12688 1156 12700
rect 1111 12660 1156 12688
rect 1150 12648 1156 12660
rect 1208 12648 1214 12700
rect 3361 12691 3419 12697
rect 3361 12657 3373 12691
rect 3407 12688 3419 12691
rect 4526 12688 4554 12796
rect 14950 12784 14956 12796
rect 15008 12784 15014 12836
rect 15873 12827 15931 12833
rect 15873 12793 15885 12827
rect 15919 12824 15931 12827
rect 16146 12824 16152 12836
rect 15919 12796 16152 12824
rect 15919 12793 15931 12796
rect 15873 12787 15931 12793
rect 16146 12784 16152 12796
rect 16204 12784 16210 12836
rect 26913 12827 26971 12833
rect 26913 12793 26925 12827
rect 26959 12824 26971 12827
rect 27002 12824 27008 12836
rect 26959 12796 27008 12824
rect 26959 12793 26971 12796
rect 26913 12787 26971 12793
rect 27002 12784 27008 12796
rect 27060 12784 27066 12836
rect 28658 12784 28664 12836
rect 28716 12824 28722 12836
rect 28716 12796 29164 12824
rect 28716 12784 28722 12796
rect 29136 12768 29164 12796
rect 8050 12756 8056 12768
rect 4646 12688 4652 12700
rect 3407 12660 4652 12688
rect 3407 12657 3419 12660
rect 3361 12651 3419 12657
rect 4646 12648 4652 12660
rect 4704 12648 4710 12700
rect 7332 12688 7360 12756
rect 8011 12728 8056 12756
rect 8050 12716 8056 12728
rect 8108 12716 8114 12768
rect 11454 12716 11460 12768
rect 11512 12756 11518 12768
rect 11917 12759 11975 12765
rect 11917 12756 11929 12759
rect 11512 12728 11929 12756
rect 11512 12716 11518 12728
rect 11917 12725 11929 12728
rect 11963 12725 11975 12759
rect 11917 12719 11975 12725
rect 12101 12759 12159 12765
rect 12101 12725 12113 12759
rect 12147 12756 12159 12759
rect 12282 12756 12288 12768
rect 12147 12728 12288 12756
rect 12147 12725 12159 12728
rect 12101 12719 12159 12725
rect 7406 12688 7412 12700
rect 7319 12660 7412 12688
rect 7406 12648 7412 12660
rect 7464 12688 7470 12700
rect 7958 12688 7964 12700
rect 7464 12660 7964 12688
rect 7464 12648 7470 12660
rect 7958 12648 7964 12660
rect 8016 12648 8022 12700
rect 11270 12648 11276 12700
rect 11328 12648 11334 12700
rect 11932 12688 11960 12719
rect 12282 12716 12288 12728
rect 12340 12716 12346 12768
rect 12374 12716 12380 12768
rect 12432 12756 12438 12768
rect 12745 12759 12803 12765
rect 12745 12756 12757 12759
rect 12432 12728 12757 12756
rect 12432 12716 12438 12728
rect 12745 12725 12757 12728
rect 12791 12725 12803 12759
rect 15597 12759 15655 12765
rect 15597 12756 15609 12759
rect 12745 12719 12803 12725
rect 14600 12728 15609 12756
rect 12466 12688 12472 12700
rect 11932 12660 12472 12688
rect 12466 12648 12472 12660
rect 12524 12688 12530 12700
rect 12834 12688 12840 12700
rect 12524 12660 12840 12688
rect 12524 12648 12530 12660
rect 12834 12648 12840 12660
rect 12892 12688 12898 12700
rect 12929 12691 12987 12697
rect 12929 12688 12941 12691
rect 12892 12660 12941 12688
rect 12892 12648 12898 12660
rect 12929 12657 12941 12660
rect 12975 12657 12987 12691
rect 12929 12651 12987 12657
rect 14214 12648 14220 12700
rect 14272 12688 14278 12700
rect 14600 12697 14628 12728
rect 15597 12725 15609 12728
rect 15643 12756 15655 12759
rect 15778 12756 15784 12768
rect 15643 12728 15784 12756
rect 15643 12725 15655 12728
rect 15597 12719 15655 12725
rect 15778 12716 15784 12728
rect 15836 12716 15842 12768
rect 17342 12756 17348 12768
rect 17268 12728 17348 12756
rect 14585 12691 14643 12697
rect 14585 12688 14597 12691
rect 14272 12660 14597 12688
rect 14272 12648 14278 12660
rect 14585 12657 14597 12660
rect 14631 12657 14643 12691
rect 14766 12688 14772 12700
rect 14727 12660 14772 12688
rect 14585 12651 14643 12657
rect 14766 12648 14772 12660
rect 14824 12648 14830 12700
rect 14861 12691 14919 12697
rect 14861 12657 14873 12691
rect 14907 12688 14919 12691
rect 14950 12688 14956 12700
rect 14907 12660 14956 12688
rect 14907 12657 14919 12660
rect 14861 12651 14919 12657
rect 14950 12648 14956 12660
rect 15008 12648 15014 12700
rect 15226 12648 15232 12700
rect 15284 12688 15290 12700
rect 15321 12691 15379 12697
rect 15321 12688 15333 12691
rect 15284 12660 15333 12688
rect 15284 12648 15290 12660
rect 15321 12657 15333 12660
rect 15367 12688 15379 12691
rect 16330 12688 16336 12700
rect 15367 12660 16336 12688
rect 15367 12657 15379 12660
rect 15321 12651 15379 12657
rect 16330 12648 16336 12660
rect 16388 12688 16394 12700
rect 17268 12697 17296 12728
rect 17342 12716 17348 12728
rect 17400 12716 17406 12768
rect 18538 12716 18544 12768
rect 18596 12756 18602 12768
rect 18725 12759 18783 12765
rect 18725 12756 18737 12759
rect 18596 12728 18737 12756
rect 18596 12716 18602 12728
rect 18725 12725 18737 12728
rect 18771 12756 18783 12759
rect 18771 12728 21804 12756
rect 18771 12725 18783 12728
rect 18725 12719 18783 12725
rect 16885 12691 16943 12697
rect 16885 12688 16897 12691
rect 16388 12660 16897 12688
rect 16388 12648 16394 12660
rect 16885 12657 16897 12660
rect 16931 12657 16943 12691
rect 16885 12651 16943 12657
rect 17253 12691 17311 12697
rect 17253 12657 17265 12691
rect 17299 12657 17311 12691
rect 17253 12651 17311 12657
rect 18814 12648 18820 12700
rect 18872 12688 18878 12700
rect 21776 12697 21804 12728
rect 29118 12716 29124 12768
rect 29176 12716 29182 12768
rect 18909 12691 18967 12697
rect 18909 12688 18921 12691
rect 18872 12660 18921 12688
rect 18872 12648 18878 12660
rect 18909 12657 18921 12660
rect 18955 12657 18967 12691
rect 18909 12651 18967 12657
rect 21761 12691 21819 12697
rect 21761 12657 21773 12691
rect 21807 12688 21819 12691
rect 21942 12688 21948 12700
rect 21807 12660 21948 12688
rect 21807 12657 21819 12660
rect 21761 12651 21819 12657
rect 21942 12648 21948 12660
rect 22000 12688 22006 12700
rect 23414 12688 23420 12700
rect 22000 12660 23420 12688
rect 22000 12648 22006 12660
rect 23414 12648 23420 12660
rect 23472 12648 23478 12700
rect 24334 12688 24340 12700
rect 24295 12660 24340 12688
rect 24334 12648 24340 12660
rect 24392 12648 24398 12700
rect 24702 12688 24708 12700
rect 24663 12660 24708 12688
rect 24702 12648 24708 12660
rect 24760 12648 24766 12700
rect 24889 12691 24947 12697
rect 24889 12657 24901 12691
rect 24935 12688 24947 12691
rect 25254 12688 25260 12700
rect 24935 12660 25260 12688
rect 24935 12657 24947 12660
rect 24889 12651 24947 12657
rect 1429 12623 1487 12629
rect 1429 12589 1441 12623
rect 1475 12620 1487 12623
rect 1702 12620 1708 12632
rect 1475 12592 1708 12620
rect 1475 12589 1487 12592
rect 1429 12583 1487 12589
rect 1702 12580 1708 12592
rect 1760 12580 1766 12632
rect 3266 12580 3272 12632
rect 3324 12620 3330 12632
rect 3545 12623 3603 12629
rect 3545 12620 3557 12623
rect 3324 12592 3557 12620
rect 3324 12580 3330 12592
rect 3545 12589 3557 12592
rect 3591 12589 3603 12623
rect 4830 12620 4836 12632
rect 4791 12592 4836 12620
rect 3545 12583 3603 12589
rect 4830 12580 4836 12592
rect 4888 12620 4894 12632
rect 5842 12620 5848 12632
rect 4888 12592 5848 12620
rect 4888 12580 4894 12592
rect 5842 12580 5848 12592
rect 5900 12580 5906 12632
rect 5937 12623 5995 12629
rect 5937 12589 5949 12623
rect 5983 12620 5995 12623
rect 6118 12620 6124 12632
rect 5983 12592 6124 12620
rect 5983 12589 5995 12592
rect 5937 12583 5995 12589
rect 6118 12580 6124 12592
rect 6176 12580 6182 12632
rect 6302 12620 6308 12632
rect 6263 12592 6308 12620
rect 6302 12580 6308 12592
rect 6360 12580 6366 12632
rect 9890 12620 9896 12632
rect 9851 12592 9896 12620
rect 9890 12580 9896 12592
rect 9948 12580 9954 12632
rect 10169 12623 10227 12629
rect 10169 12589 10181 12623
rect 10215 12620 10227 12623
rect 10810 12620 10816 12632
rect 10215 12592 10816 12620
rect 10215 12589 10227 12592
rect 10169 12583 10227 12589
rect 10810 12580 10816 12592
rect 10868 12580 10874 12632
rect 13294 12620 13300 12632
rect 13255 12592 13300 12620
rect 13294 12580 13300 12592
rect 13352 12580 13358 12632
rect 15505 12623 15563 12629
rect 15505 12589 15517 12623
rect 15551 12620 15563 12623
rect 16606 12620 16612 12632
rect 15551 12592 16612 12620
rect 15551 12589 15563 12592
rect 15505 12583 15563 12589
rect 16606 12580 16612 12592
rect 16664 12580 16670 12632
rect 16974 12620 16980 12632
rect 16935 12592 16980 12620
rect 16974 12580 16980 12592
rect 17032 12580 17038 12632
rect 17342 12620 17348 12632
rect 17303 12592 17348 12620
rect 17342 12580 17348 12592
rect 17400 12580 17406 12632
rect 18170 12580 18176 12632
rect 18228 12620 18234 12632
rect 19550 12620 19556 12632
rect 18228 12592 19556 12620
rect 18228 12580 18234 12592
rect 19550 12580 19556 12592
rect 19608 12580 19614 12632
rect 24150 12620 24156 12632
rect 24111 12592 24156 12620
rect 24150 12580 24156 12592
rect 24208 12580 24214 12632
rect 23138 12512 23144 12564
rect 23196 12552 23202 12564
rect 24904 12552 24932 12651
rect 25254 12648 25260 12660
rect 25312 12648 25318 12700
rect 27097 12691 27155 12697
rect 27097 12657 27109 12691
rect 27143 12688 27155 12691
rect 27370 12688 27376 12700
rect 27143 12660 27376 12688
rect 27143 12657 27155 12660
rect 27097 12651 27155 12657
rect 27370 12648 27376 12660
rect 27428 12648 27434 12700
rect 26358 12580 26364 12632
rect 26416 12620 26422 12632
rect 28382 12620 28388 12632
rect 26416 12592 28388 12620
rect 26416 12580 26422 12592
rect 28382 12580 28388 12592
rect 28440 12580 28446 12632
rect 28750 12620 28756 12632
rect 28711 12592 28756 12620
rect 28750 12580 28756 12592
rect 28808 12580 28814 12632
rect 30130 12620 30136 12632
rect 30091 12592 30136 12620
rect 30130 12580 30136 12592
rect 30188 12580 30194 12632
rect 23196 12524 24932 12552
rect 23196 12512 23202 12524
rect 8237 12487 8295 12493
rect 8237 12453 8249 12487
rect 8283 12484 8295 12487
rect 8510 12484 8516 12496
rect 8283 12456 8516 12484
rect 8283 12453 8295 12456
rect 8237 12447 8295 12453
rect 8510 12444 8516 12456
rect 8568 12444 8574 12496
rect 16333 12487 16391 12493
rect 16333 12453 16345 12487
rect 16379 12484 16391 12487
rect 16422 12484 16428 12496
rect 16379 12456 16428 12484
rect 16379 12453 16391 12456
rect 16333 12447 16391 12453
rect 16422 12444 16428 12456
rect 16480 12444 16486 12496
rect 18446 12444 18452 12496
rect 18504 12484 18510 12496
rect 19001 12487 19059 12493
rect 19001 12484 19013 12487
rect 18504 12456 19013 12484
rect 18504 12444 18510 12456
rect 19001 12453 19013 12456
rect 19047 12484 19059 12487
rect 19458 12484 19464 12496
rect 19047 12456 19464 12484
rect 19047 12453 19059 12456
rect 19001 12447 19059 12453
rect 19458 12444 19464 12456
rect 19516 12444 19522 12496
rect 20562 12444 20568 12496
rect 20620 12484 20626 12496
rect 20657 12487 20715 12493
rect 20657 12484 20669 12487
rect 20620 12456 20669 12484
rect 20620 12444 20626 12456
rect 20657 12453 20669 12456
rect 20703 12453 20715 12487
rect 21758 12484 21764 12496
rect 21719 12456 21764 12484
rect 20657 12447 20715 12453
rect 21758 12444 21764 12456
rect 21816 12444 21822 12496
rect 23601 12487 23659 12493
rect 23601 12453 23613 12487
rect 23647 12484 23659 12487
rect 23874 12484 23880 12496
rect 23647 12456 23880 12484
rect 23647 12453 23659 12456
rect 23601 12447 23659 12453
rect 23874 12444 23880 12456
rect 23932 12484 23938 12496
rect 23969 12487 24027 12493
rect 23969 12484 23981 12487
rect 23932 12456 23981 12484
rect 23932 12444 23938 12456
rect 23969 12453 23981 12456
rect 24015 12453 24027 12487
rect 23969 12447 24027 12453
rect 400 12394 31680 12416
rect 400 12342 3510 12394
rect 3562 12342 3574 12394
rect 3626 12342 3638 12394
rect 3690 12342 3702 12394
rect 3754 12342 3766 12394
rect 3818 12342 31680 12394
rect 400 12320 31680 12342
rect 1702 12280 1708 12292
rect 1663 12252 1708 12280
rect 1702 12240 1708 12252
rect 1760 12240 1766 12292
rect 3637 12283 3695 12289
rect 3637 12280 3649 12283
rect 3008 12252 3649 12280
rect 1242 12144 1248 12156
rect 1203 12116 1248 12144
rect 1242 12104 1248 12116
rect 1300 12144 1306 12156
rect 3008 12153 3036 12252
rect 3637 12249 3649 12252
rect 3683 12280 3695 12283
rect 4094 12280 4100 12292
rect 3683 12252 4100 12280
rect 3683 12249 3695 12252
rect 3637 12243 3695 12249
rect 4094 12240 4100 12252
rect 4152 12240 4158 12292
rect 4646 12280 4652 12292
rect 4526 12252 4652 12280
rect 3453 12215 3511 12221
rect 3453 12181 3465 12215
rect 3499 12212 3511 12215
rect 4526 12212 4554 12252
rect 4646 12240 4652 12252
rect 4704 12240 4710 12292
rect 6302 12240 6308 12292
rect 6360 12280 6366 12292
rect 6397 12283 6455 12289
rect 6397 12280 6409 12283
rect 6360 12252 6409 12280
rect 6360 12240 6366 12252
rect 6397 12249 6409 12252
rect 6443 12249 6455 12283
rect 10534 12280 10540 12292
rect 6397 12243 6455 12249
rect 8160 12252 10540 12280
rect 3499 12184 4554 12212
rect 3499 12181 3511 12184
rect 3453 12175 3511 12181
rect 8160 12156 8188 12252
rect 10534 12240 10540 12252
rect 10592 12240 10598 12292
rect 10810 12280 10816 12292
rect 10771 12252 10816 12280
rect 10810 12240 10816 12252
rect 10868 12240 10874 12292
rect 12374 12240 12380 12292
rect 12432 12280 12438 12292
rect 12929 12283 12987 12289
rect 12929 12280 12941 12283
rect 12432 12252 12941 12280
rect 12432 12240 12438 12252
rect 12929 12249 12941 12252
rect 12975 12280 12987 12283
rect 13113 12283 13171 12289
rect 13113 12280 13125 12283
rect 12975 12252 13125 12280
rect 12975 12249 12987 12252
rect 12929 12243 12987 12249
rect 13113 12249 13125 12252
rect 13159 12249 13171 12283
rect 13294 12280 13300 12292
rect 13255 12252 13300 12280
rect 13113 12243 13171 12249
rect 13294 12240 13300 12252
rect 13352 12280 13358 12292
rect 14766 12280 14772 12292
rect 13352 12252 14772 12280
rect 13352 12240 13358 12252
rect 14766 12240 14772 12252
rect 14824 12240 14830 12292
rect 15226 12280 15232 12292
rect 15187 12252 15232 12280
rect 15226 12240 15232 12252
rect 15284 12240 15290 12292
rect 15597 12283 15655 12289
rect 15597 12249 15609 12283
rect 15643 12280 15655 12283
rect 16146 12280 16152 12292
rect 15643 12252 16152 12280
rect 15643 12249 15655 12252
rect 15597 12243 15655 12249
rect 16146 12240 16152 12252
rect 16204 12240 16210 12292
rect 16606 12280 16612 12292
rect 16567 12252 16612 12280
rect 16606 12240 16612 12252
rect 16664 12240 16670 12292
rect 16974 12240 16980 12292
rect 17032 12280 17038 12292
rect 17069 12283 17127 12289
rect 17069 12280 17081 12283
rect 17032 12252 17081 12280
rect 17032 12240 17038 12252
rect 17069 12249 17081 12252
rect 17115 12249 17127 12283
rect 18446 12280 18452 12292
rect 18407 12252 18452 12280
rect 17069 12243 17127 12249
rect 18446 12240 18452 12252
rect 18504 12240 18510 12292
rect 18722 12240 18728 12292
rect 18780 12280 18786 12292
rect 19185 12283 19243 12289
rect 19185 12280 19197 12283
rect 18780 12252 19197 12280
rect 18780 12240 18786 12252
rect 19185 12249 19197 12252
rect 19231 12249 19243 12283
rect 21942 12280 21948 12292
rect 21903 12252 21948 12280
rect 19185 12243 19243 12249
rect 21942 12240 21948 12252
rect 22000 12240 22006 12292
rect 23049 12283 23107 12289
rect 23049 12249 23061 12283
rect 23095 12280 23107 12283
rect 24702 12280 24708 12292
rect 23095 12252 24708 12280
rect 23095 12249 23107 12252
rect 23049 12243 23107 12249
rect 24702 12240 24708 12252
rect 24760 12240 24766 12292
rect 27002 12240 27008 12292
rect 27060 12280 27066 12292
rect 27557 12283 27615 12289
rect 27557 12280 27569 12283
rect 27060 12252 27569 12280
rect 27060 12240 27066 12252
rect 27557 12249 27569 12252
rect 27603 12249 27615 12283
rect 27557 12243 27615 12249
rect 27833 12283 27891 12289
rect 27833 12249 27845 12283
rect 27879 12280 27891 12283
rect 28750 12280 28756 12292
rect 27879 12252 28756 12280
rect 27879 12249 27891 12252
rect 27833 12243 27891 12249
rect 28750 12240 28756 12252
rect 28808 12280 28814 12292
rect 28845 12283 28903 12289
rect 28845 12280 28857 12283
rect 28808 12252 28857 12280
rect 28808 12240 28814 12252
rect 28845 12249 28857 12252
rect 28891 12249 28903 12283
rect 28845 12243 28903 12249
rect 10629 12215 10687 12221
rect 10629 12181 10641 12215
rect 10675 12212 10687 12215
rect 11454 12212 11460 12224
rect 10675 12184 11460 12212
rect 10675 12181 10687 12184
rect 10629 12175 10687 12181
rect 11454 12172 11460 12184
rect 11512 12212 11518 12224
rect 12745 12215 12803 12221
rect 12745 12212 12757 12215
rect 11512 12184 12757 12212
rect 11512 12172 11518 12184
rect 12745 12181 12757 12184
rect 12791 12181 12803 12215
rect 12745 12175 12803 12181
rect 14214 12172 14220 12224
rect 14272 12212 14278 12224
rect 14585 12215 14643 12221
rect 14585 12212 14597 12215
rect 14272 12184 14597 12212
rect 14272 12172 14278 12184
rect 14585 12181 14597 12184
rect 14631 12181 14643 12215
rect 18538 12212 18544 12224
rect 18499 12184 18544 12212
rect 14585 12175 14643 12181
rect 18538 12172 18544 12184
rect 18596 12172 18602 12224
rect 21022 12172 21028 12224
rect 21080 12212 21086 12224
rect 23138 12212 23144 12224
rect 21080 12184 23144 12212
rect 21080 12172 21086 12184
rect 23138 12172 23144 12184
rect 23196 12172 23202 12224
rect 28382 12172 28388 12224
rect 28440 12212 28446 12224
rect 29857 12215 29915 12221
rect 29857 12212 29869 12215
rect 28440 12184 29869 12212
rect 28440 12172 28446 12184
rect 29857 12181 29869 12184
rect 29903 12181 29915 12215
rect 29857 12175 29915 12181
rect 1521 12147 1579 12153
rect 1521 12144 1533 12147
rect 1300 12116 1533 12144
rect 1300 12104 1306 12116
rect 1521 12113 1533 12116
rect 1567 12113 1579 12147
rect 1521 12107 1579 12113
rect 2993 12147 3051 12153
rect 2993 12113 3005 12147
rect 3039 12113 3051 12147
rect 2993 12107 3051 12113
rect 5106 12104 5112 12156
rect 5164 12144 5170 12156
rect 5569 12147 5627 12153
rect 5569 12144 5581 12147
rect 5164 12116 5581 12144
rect 5164 12104 5170 12116
rect 5569 12113 5581 12116
rect 5615 12144 5627 12147
rect 5753 12147 5811 12153
rect 5753 12144 5765 12147
rect 5615 12116 5765 12144
rect 5615 12113 5627 12116
rect 5569 12107 5627 12113
rect 5753 12113 5765 12116
rect 5799 12144 5811 12147
rect 8142 12144 8148 12156
rect 5799 12116 7360 12144
rect 8055 12116 8148 12144
rect 5799 12113 5811 12116
rect 5753 12107 5811 12113
rect 2717 12079 2775 12085
rect 2717 12076 2729 12079
rect 2548 12048 2729 12076
rect 1150 11900 1156 11952
rect 1208 11940 1214 11952
rect 1981 11943 2039 11949
rect 1981 11940 1993 11943
rect 1208 11912 1993 11940
rect 1208 11900 1214 11912
rect 1981 11909 1993 11912
rect 2027 11940 2039 11943
rect 2438 11940 2444 11952
rect 2027 11912 2444 11940
rect 2027 11909 2039 11912
rect 1981 11903 2039 11909
rect 2438 11900 2444 11912
rect 2496 11940 2502 11952
rect 2548 11949 2576 12048
rect 2717 12045 2729 12048
rect 2763 12076 2775 12079
rect 3266 12076 3272 12088
rect 2763 12048 3272 12076
rect 2763 12045 2775 12048
rect 2717 12039 2775 12045
rect 3266 12036 3272 12048
rect 3324 12076 3330 12088
rect 3729 12079 3787 12085
rect 3729 12076 3741 12079
rect 3324 12048 3741 12076
rect 3324 12036 3330 12048
rect 3729 12045 3741 12048
rect 3775 12045 3787 12079
rect 3729 12039 3787 12045
rect 5201 12079 5259 12085
rect 5201 12045 5213 12079
rect 5247 12076 5259 12079
rect 6118 12076 6124 12088
rect 5247 12048 6124 12076
rect 5247 12045 5259 12048
rect 5201 12039 5259 12045
rect 6118 12036 6124 12048
rect 6176 12036 6182 12088
rect 6578 12076 6584 12088
rect 6539 12048 6584 12076
rect 6578 12036 6584 12048
rect 6636 12036 6642 12088
rect 6762 12076 6768 12088
rect 6723 12048 6768 12076
rect 6762 12036 6768 12048
rect 6820 12036 6826 12088
rect 7332 12085 7360 12116
rect 8142 12104 8148 12116
rect 8200 12104 8206 12156
rect 8510 12144 8516 12156
rect 8471 12116 8516 12144
rect 8510 12104 8516 12116
rect 8568 12104 8574 12156
rect 9798 12104 9804 12156
rect 9856 12144 9862 12156
rect 9893 12147 9951 12153
rect 9893 12144 9905 12147
rect 9856 12116 9905 12144
rect 9856 12104 9862 12116
rect 9893 12113 9905 12116
rect 9939 12113 9951 12147
rect 9893 12107 9951 12113
rect 10445 12147 10503 12153
rect 10445 12113 10457 12147
rect 10491 12144 10503 12147
rect 11270 12144 11276 12156
rect 10491 12116 11276 12144
rect 10491 12113 10503 12116
rect 10445 12107 10503 12113
rect 7133 12079 7191 12085
rect 7133 12045 7145 12079
rect 7179 12045 7191 12079
rect 7133 12039 7191 12045
rect 7317 12079 7375 12085
rect 7317 12045 7329 12079
rect 7363 12076 7375 12079
rect 8050 12076 8056 12088
rect 7363 12048 8056 12076
rect 7363 12045 7375 12048
rect 7317 12039 7375 12045
rect 5385 12011 5443 12017
rect 5385 11977 5397 12011
rect 5431 12008 5443 12011
rect 7148 12008 7176 12039
rect 8050 12036 8056 12048
rect 8108 12036 8114 12088
rect 10460 12076 10488 12107
rect 11270 12104 11276 12116
rect 11328 12104 11334 12156
rect 14030 12104 14036 12156
rect 14088 12144 14094 12156
rect 15689 12147 15747 12153
rect 15689 12144 15701 12147
rect 14088 12116 15701 12144
rect 14088 12104 14094 12116
rect 15689 12113 15701 12116
rect 15735 12144 15747 12147
rect 16885 12147 16943 12153
rect 16885 12144 16897 12147
rect 15735 12116 16897 12144
rect 15735 12113 15747 12116
rect 15689 12107 15747 12113
rect 12374 12076 12380 12088
rect 9540 12048 10488 12076
rect 12335 12048 12380 12076
rect 7866 12008 7872 12020
rect 5431 11980 7872 12008
rect 5431 11977 5443 11980
rect 5385 11971 5443 11977
rect 7866 11968 7872 11980
rect 7924 11968 7930 12020
rect 2533 11943 2591 11949
rect 2533 11940 2545 11943
rect 2496 11912 2545 11940
rect 2496 11900 2502 11912
rect 2533 11909 2545 11912
rect 2579 11909 2591 11943
rect 4830 11940 4836 11952
rect 4791 11912 4836 11940
rect 2533 11903 2591 11909
rect 4830 11900 4836 11912
rect 4888 11900 4894 11952
rect 5934 11940 5940 11952
rect 5895 11912 5940 11940
rect 5934 11900 5940 11912
rect 5992 11900 5998 11952
rect 7682 11900 7688 11952
rect 7740 11940 7746 11952
rect 7777 11943 7835 11949
rect 7777 11940 7789 11943
rect 7740 11912 7789 11940
rect 7740 11900 7746 11912
rect 7777 11909 7789 11912
rect 7823 11909 7835 11943
rect 7777 11903 7835 11909
rect 7958 11900 7964 11952
rect 8016 11940 8022 11952
rect 8053 11943 8111 11949
rect 8053 11940 8065 11943
rect 8016 11912 8065 11940
rect 8016 11900 8022 11912
rect 8053 11909 8065 11912
rect 8099 11940 8111 11943
rect 8786 11940 8792 11952
rect 8099 11912 8792 11940
rect 8099 11909 8111 11912
rect 8053 11903 8111 11909
rect 8786 11900 8792 11912
rect 8844 11940 8850 11952
rect 9540 11940 9568 12048
rect 12374 12036 12380 12048
rect 12432 12036 12438 12088
rect 15980 12085 16008 12116
rect 16885 12113 16897 12116
rect 16931 12144 16943 12147
rect 17342 12144 17348 12156
rect 16931 12116 17348 12144
rect 16931 12113 16943 12116
rect 16885 12107 16943 12113
rect 17342 12104 17348 12116
rect 17400 12104 17406 12156
rect 17618 12104 17624 12156
rect 17676 12144 17682 12156
rect 19737 12147 19795 12153
rect 19737 12144 19749 12147
rect 17676 12116 19749 12144
rect 17676 12104 17682 12116
rect 15873 12079 15931 12085
rect 15873 12045 15885 12079
rect 15919 12045 15931 12079
rect 15873 12039 15931 12045
rect 15965 12079 16023 12085
rect 15965 12045 15977 12079
rect 16011 12045 16023 12079
rect 15965 12039 16023 12045
rect 14030 11968 14036 12020
rect 14088 12008 14094 12020
rect 15888 12008 15916 12039
rect 17434 12036 17440 12088
rect 17492 12076 17498 12088
rect 18725 12079 18783 12085
rect 18725 12076 18737 12079
rect 17492 12048 18737 12076
rect 17492 12036 17498 12048
rect 18725 12045 18737 12048
rect 18771 12076 18783 12079
rect 18814 12076 18820 12088
rect 18771 12048 18820 12076
rect 18771 12045 18783 12048
rect 18725 12039 18783 12045
rect 18814 12036 18820 12048
rect 18872 12036 18878 12088
rect 18924 12085 18952 12116
rect 19737 12113 19749 12116
rect 19783 12113 19795 12147
rect 19737 12107 19795 12113
rect 20565 12147 20623 12153
rect 20565 12113 20577 12147
rect 20611 12144 20623 12147
rect 20611 12116 21896 12144
rect 20611 12113 20623 12116
rect 20565 12107 20623 12113
rect 21868 12088 21896 12116
rect 23230 12104 23236 12156
rect 23288 12144 23294 12156
rect 24242 12144 24248 12156
rect 23288 12116 24248 12144
rect 23288 12104 23294 12116
rect 24242 12104 24248 12116
rect 24300 12104 24306 12156
rect 25254 12144 25260 12156
rect 25215 12116 25260 12144
rect 25254 12104 25260 12116
rect 25312 12104 25318 12156
rect 26818 12104 26824 12156
rect 26876 12144 26882 12156
rect 27005 12147 27063 12153
rect 27005 12144 27017 12147
rect 26876 12116 27017 12144
rect 26876 12104 26882 12116
rect 27005 12113 27017 12116
rect 27051 12113 27063 12147
rect 27005 12107 27063 12113
rect 28017 12147 28075 12153
rect 28017 12113 28029 12147
rect 28063 12144 28075 12147
rect 28201 12147 28259 12153
rect 28201 12144 28213 12147
rect 28063 12116 28213 12144
rect 28063 12113 28075 12116
rect 28017 12107 28075 12113
rect 28201 12113 28213 12116
rect 28247 12144 28259 12147
rect 28934 12144 28940 12156
rect 28247 12116 28940 12144
rect 28247 12113 28259 12116
rect 28201 12107 28259 12113
rect 28934 12104 28940 12116
rect 28992 12144 28998 12156
rect 28992 12116 29808 12144
rect 28992 12104 28998 12116
rect 18909 12079 18967 12085
rect 18909 12045 18921 12079
rect 18955 12045 18967 12079
rect 18909 12039 18967 12045
rect 19093 12079 19151 12085
rect 19093 12045 19105 12079
rect 19139 12076 19151 12079
rect 19139 12048 19504 12076
rect 19139 12045 19151 12048
rect 19093 12039 19151 12045
rect 16701 12011 16759 12017
rect 16701 12008 16713 12011
rect 14088 11980 16713 12008
rect 14088 11968 14094 11980
rect 16701 11977 16713 11980
rect 16747 12008 16759 12011
rect 17802 12008 17808 12020
rect 16747 11980 17808 12008
rect 16747 11977 16759 11980
rect 16701 11971 16759 11977
rect 17802 11968 17808 11980
rect 17860 11968 17866 12020
rect 19476 11952 19504 12048
rect 20746 12036 20752 12088
rect 20804 12076 20810 12088
rect 21117 12079 21175 12085
rect 21117 12076 21129 12079
rect 20804 12048 21129 12076
rect 20804 12036 20810 12048
rect 21117 12045 21129 12048
rect 21163 12045 21175 12079
rect 21298 12076 21304 12088
rect 21259 12048 21304 12076
rect 21117 12039 21175 12045
rect 21298 12036 21304 12048
rect 21356 12036 21362 12088
rect 21666 12076 21672 12088
rect 21579 12048 21672 12076
rect 21666 12036 21672 12048
rect 21724 12036 21730 12088
rect 21850 12076 21856 12088
rect 21763 12048 21856 12076
rect 21850 12036 21856 12048
rect 21908 12076 21914 12088
rect 23046 12076 23052 12088
rect 21908 12048 23052 12076
rect 21908 12036 21914 12048
rect 23046 12036 23052 12048
rect 23104 12036 23110 12088
rect 23506 12076 23512 12088
rect 23467 12048 23512 12076
rect 23506 12036 23512 12048
rect 23564 12036 23570 12088
rect 23874 12036 23880 12088
rect 23932 12076 23938 12088
rect 26453 12079 26511 12085
rect 23932 12048 23977 12076
rect 23932 12036 23938 12048
rect 26453 12045 26465 12079
rect 26499 12076 26511 12079
rect 26836 12076 26864 12104
rect 27278 12076 27284 12088
rect 26499 12048 26864 12076
rect 26928 12048 27284 12076
rect 26499 12045 26511 12048
rect 26453 12039 26511 12045
rect 20381 12011 20439 12017
rect 20381 11977 20393 12011
rect 20427 12008 20439 12011
rect 20654 12008 20660 12020
rect 20427 11980 20660 12008
rect 20427 11977 20439 11980
rect 20381 11971 20439 11977
rect 20654 11968 20660 11980
rect 20712 11968 20718 12020
rect 8844 11912 9568 11940
rect 12101 11943 12159 11949
rect 8844 11900 8850 11912
rect 12101 11909 12113 11943
rect 12147 11940 12159 11943
rect 12285 11943 12343 11949
rect 12285 11940 12297 11943
rect 12147 11912 12297 11940
rect 12147 11909 12159 11912
rect 12101 11903 12159 11909
rect 12285 11909 12297 11912
rect 12331 11940 12343 11943
rect 12558 11940 12564 11952
rect 12331 11912 12564 11940
rect 12331 11909 12343 11912
rect 12285 11903 12343 11909
rect 12558 11900 12564 11912
rect 12616 11900 12622 11952
rect 14950 11940 14956 11952
rect 14911 11912 14956 11940
rect 14950 11900 14956 11912
rect 15008 11900 15014 11952
rect 19458 11900 19464 11952
rect 19516 11940 19522 11952
rect 19553 11943 19611 11949
rect 19553 11940 19565 11943
rect 19516 11912 19565 11940
rect 19516 11900 19522 11912
rect 19553 11909 19565 11912
rect 19599 11909 19611 11943
rect 20102 11940 20108 11952
rect 20063 11912 20108 11940
rect 19553 11903 19611 11909
rect 20102 11900 20108 11912
rect 20160 11900 20166 11952
rect 20562 11900 20568 11952
rect 20620 11940 20626 11952
rect 21684 11940 21712 12036
rect 21758 11968 21764 12020
rect 21816 12008 21822 12020
rect 22221 12011 22279 12017
rect 22221 12008 22233 12011
rect 21816 11980 22233 12008
rect 21816 11968 21822 11980
rect 22221 11977 22233 11980
rect 22267 12008 22279 12011
rect 22267 11980 23460 12008
rect 22267 11977 22279 11980
rect 22221 11971 22279 11977
rect 20620 11912 21712 11940
rect 20620 11900 20626 11912
rect 23230 11900 23236 11952
rect 23288 11940 23294 11952
rect 23325 11943 23383 11949
rect 23325 11940 23337 11943
rect 23288 11912 23337 11940
rect 23288 11900 23294 11912
rect 23325 11909 23337 11912
rect 23371 11909 23383 11943
rect 23432 11940 23460 11980
rect 24242 11968 24248 12020
rect 24300 11968 24306 12020
rect 26468 11940 26496 12039
rect 26726 12008 26732 12020
rect 26639 11980 26732 12008
rect 26726 11968 26732 11980
rect 26784 12008 26790 12020
rect 26928 12008 26956 12048
rect 27278 12036 27284 12048
rect 27336 12036 27342 12088
rect 29029 12079 29087 12085
rect 29029 12045 29041 12079
rect 29075 12045 29087 12079
rect 29210 12076 29216 12088
rect 29171 12048 29216 12076
rect 29029 12039 29087 12045
rect 26784 11980 26956 12008
rect 26784 11968 26790 11980
rect 27186 11968 27192 12020
rect 27244 12008 27250 12020
rect 28293 12011 28351 12017
rect 28293 12008 28305 12011
rect 27244 11980 28305 12008
rect 27244 11968 27250 11980
rect 28293 11977 28305 11980
rect 28339 12008 28351 12011
rect 28566 12008 28572 12020
rect 28339 11980 28572 12008
rect 28339 11977 28351 11980
rect 28293 11971 28351 11977
rect 28566 11968 28572 11980
rect 28624 11968 28630 12020
rect 29044 12008 29072 12039
rect 29210 12036 29216 12048
rect 29268 12036 29274 12088
rect 29578 12076 29584 12088
rect 29539 12048 29584 12076
rect 29578 12036 29584 12048
rect 29636 12036 29642 12088
rect 29780 12085 29808 12116
rect 29765 12079 29823 12085
rect 29765 12045 29777 12079
rect 29811 12076 29823 12079
rect 30130 12076 30136 12088
rect 29811 12048 30136 12076
rect 29811 12045 29823 12048
rect 29765 12039 29823 12045
rect 30130 12036 30136 12048
rect 30188 12036 30194 12088
rect 29118 12008 29124 12020
rect 29044 11980 29124 12008
rect 29118 11968 29124 11980
rect 29176 11968 29182 12020
rect 27370 11940 27376 11952
rect 23432 11912 26496 11940
rect 27331 11912 27376 11940
rect 23325 11903 23383 11909
rect 27370 11900 27376 11912
rect 27428 11900 27434 11952
rect 400 11850 31680 11872
rect 400 11798 18870 11850
rect 18922 11798 18934 11850
rect 18986 11798 18998 11850
rect 19050 11798 19062 11850
rect 19114 11798 19126 11850
rect 19178 11798 31680 11850
rect 400 11776 31680 11798
rect 6029 11739 6087 11745
rect 6029 11705 6041 11739
rect 6075 11736 6087 11739
rect 6302 11736 6308 11748
rect 6075 11708 6308 11736
rect 6075 11705 6087 11708
rect 6029 11699 6087 11705
rect 6302 11696 6308 11708
rect 6360 11696 6366 11748
rect 8142 11736 8148 11748
rect 8103 11708 8148 11736
rect 8142 11696 8148 11708
rect 8200 11696 8206 11748
rect 9890 11696 9896 11748
rect 9948 11736 9954 11748
rect 10261 11739 10319 11745
rect 10261 11736 10273 11739
rect 9948 11708 10273 11736
rect 9948 11696 9954 11708
rect 10261 11705 10273 11708
rect 10307 11705 10319 11739
rect 16330 11736 16336 11748
rect 16291 11708 16336 11736
rect 10261 11699 10319 11705
rect 8510 11628 8516 11680
rect 8568 11668 8574 11680
rect 8973 11671 9031 11677
rect 8973 11668 8985 11671
rect 8568 11640 8985 11668
rect 8568 11628 8574 11640
rect 8973 11637 8985 11640
rect 9019 11668 9031 11671
rect 9154 11668 9160 11680
rect 9019 11640 9160 11668
rect 9019 11637 9031 11640
rect 8973 11631 9031 11637
rect 9154 11628 9160 11640
rect 9212 11628 9218 11680
rect 10276 11668 10304 11699
rect 16330 11696 16336 11708
rect 16388 11696 16394 11748
rect 16422 11696 16428 11748
rect 16480 11736 16486 11748
rect 16480 11708 16525 11736
rect 16480 11696 16486 11708
rect 16974 11696 16980 11748
rect 17032 11736 17038 11748
rect 17526 11736 17532 11748
rect 17032 11708 17532 11736
rect 17032 11696 17038 11708
rect 17526 11696 17532 11708
rect 17584 11736 17590 11748
rect 17713 11739 17771 11745
rect 17713 11736 17725 11739
rect 17584 11708 17725 11736
rect 17584 11696 17590 11708
rect 17713 11705 17725 11708
rect 17759 11705 17771 11739
rect 17713 11699 17771 11705
rect 18722 11696 18728 11748
rect 18780 11736 18786 11748
rect 18909 11739 18967 11745
rect 18909 11736 18921 11739
rect 18780 11708 18921 11736
rect 18780 11696 18786 11708
rect 18909 11705 18921 11708
rect 18955 11705 18967 11739
rect 18909 11699 18967 11705
rect 20102 11696 20108 11748
rect 20160 11736 20166 11748
rect 21298 11736 21304 11748
rect 20160 11708 21304 11736
rect 20160 11696 20166 11708
rect 21298 11696 21304 11708
rect 21356 11696 21362 11748
rect 23046 11736 23052 11748
rect 23007 11708 23052 11736
rect 23046 11696 23052 11708
rect 23104 11696 23110 11748
rect 23138 11696 23144 11748
rect 23196 11736 23202 11748
rect 23693 11739 23751 11745
rect 23693 11736 23705 11739
rect 23196 11708 23705 11736
rect 23196 11696 23202 11708
rect 23693 11705 23705 11708
rect 23739 11705 23751 11739
rect 23693 11699 23751 11705
rect 23874 11696 23880 11748
rect 23932 11736 23938 11748
rect 24150 11736 24156 11748
rect 23932 11708 23977 11736
rect 24111 11708 24156 11736
rect 23932 11696 23938 11708
rect 24150 11696 24156 11708
rect 24208 11696 24214 11748
rect 28661 11739 28719 11745
rect 26376 11708 27876 11736
rect 14398 11668 14404 11680
rect 10276 11640 14404 11668
rect 14398 11628 14404 11640
rect 14456 11668 14462 11680
rect 19274 11668 19280 11680
rect 14456 11640 19280 11668
rect 14456 11628 14462 11640
rect 19274 11628 19280 11640
rect 19332 11628 19338 11680
rect 21666 11628 21672 11680
rect 21724 11628 21730 11680
rect 24058 11628 24064 11680
rect 24116 11668 24122 11680
rect 26376 11668 26404 11708
rect 24116 11640 26404 11668
rect 24116 11628 24122 11640
rect 27186 11628 27192 11680
rect 27244 11628 27250 11680
rect 27848 11668 27876 11708
rect 28661 11705 28673 11739
rect 28707 11736 28719 11739
rect 28750 11736 28756 11748
rect 28707 11708 28756 11736
rect 28707 11705 28719 11708
rect 28661 11699 28719 11705
rect 28750 11696 28756 11708
rect 28808 11696 28814 11748
rect 28845 11671 28903 11677
rect 28845 11668 28857 11671
rect 27848 11640 28857 11668
rect 28845 11637 28857 11640
rect 28891 11668 28903 11671
rect 29118 11668 29124 11680
rect 28891 11640 29124 11668
rect 28891 11637 28903 11640
rect 28845 11631 28903 11637
rect 29118 11628 29124 11640
rect 29176 11628 29182 11680
rect 29302 11668 29308 11680
rect 29263 11640 29308 11668
rect 29302 11628 29308 11640
rect 29360 11628 29366 11680
rect 1245 11603 1303 11609
rect 1245 11569 1257 11603
rect 1291 11600 1303 11603
rect 1334 11600 1340 11612
rect 1291 11572 1340 11600
rect 1291 11569 1303 11572
rect 1245 11563 1303 11569
rect 1334 11560 1340 11572
rect 1392 11560 1398 11612
rect 9062 11560 9068 11612
rect 9120 11600 9126 11612
rect 9617 11603 9675 11609
rect 9617 11600 9629 11603
rect 9120 11572 9629 11600
rect 9120 11560 9126 11572
rect 9617 11569 9629 11572
rect 9663 11569 9675 11603
rect 9982 11600 9988 11612
rect 9943 11572 9988 11600
rect 9617 11563 9675 11569
rect 9982 11560 9988 11572
rect 10040 11560 10046 11612
rect 12558 11600 12564 11612
rect 12519 11572 12564 11600
rect 12558 11560 12564 11572
rect 12616 11560 12622 11612
rect 17618 11600 17624 11612
rect 17579 11572 17624 11600
rect 17618 11560 17624 11572
rect 17676 11560 17682 11612
rect 20654 11560 20660 11612
rect 20712 11600 20718 11612
rect 21298 11600 21304 11612
rect 20712 11572 21304 11600
rect 20712 11560 20718 11572
rect 21298 11560 21304 11572
rect 21356 11560 21362 11612
rect 29854 11600 29860 11612
rect 29366 11572 29860 11600
rect 6762 11532 6768 11544
rect 6675 11504 6768 11532
rect 6762 11492 6768 11504
rect 6820 11532 6826 11544
rect 9522 11532 9528 11544
rect 6820 11504 9528 11532
rect 6820 11492 6826 11504
rect 9522 11492 9528 11504
rect 9580 11492 9586 11544
rect 9706 11532 9712 11544
rect 9667 11504 9712 11532
rect 9706 11492 9712 11504
rect 9764 11492 9770 11544
rect 9893 11535 9951 11541
rect 9893 11501 9905 11535
rect 9939 11501 9951 11535
rect 9893 11495 9951 11501
rect 6578 11464 6584 11476
rect 6491 11436 6584 11464
rect 6578 11424 6584 11436
rect 6636 11464 6642 11476
rect 7590 11464 7596 11476
rect 6636 11436 7596 11464
rect 6636 11424 6642 11436
rect 7590 11424 7596 11436
rect 7648 11424 7654 11476
rect 8878 11424 8884 11476
rect 8936 11464 8942 11476
rect 9798 11464 9804 11476
rect 8936 11436 9804 11464
rect 8936 11424 8942 11436
rect 9798 11424 9804 11436
rect 9856 11464 9862 11476
rect 9908 11464 9936 11495
rect 12374 11492 12380 11544
rect 12432 11532 12438 11544
rect 12469 11535 12527 11541
rect 12469 11532 12481 11535
rect 12432 11504 12481 11532
rect 12432 11492 12438 11504
rect 12469 11501 12481 11504
rect 12515 11532 12527 11535
rect 14030 11532 14036 11544
rect 12515 11504 14036 11532
rect 12515 11501 12527 11504
rect 12469 11495 12527 11501
rect 14030 11492 14036 11504
rect 14088 11492 14094 11544
rect 18354 11492 18360 11544
rect 18412 11532 18418 11544
rect 20933 11535 20991 11541
rect 20933 11532 20945 11535
rect 18412 11504 20945 11532
rect 18412 11492 18418 11504
rect 20933 11501 20945 11504
rect 20979 11532 20991 11535
rect 21482 11532 21488 11544
rect 20979 11504 21488 11532
rect 20979 11501 20991 11504
rect 20933 11495 20991 11501
rect 21482 11492 21488 11504
rect 21540 11532 21546 11544
rect 22494 11532 22500 11544
rect 21540 11504 22500 11532
rect 21540 11492 21546 11504
rect 22494 11492 22500 11504
rect 22552 11532 22558 11544
rect 23506 11532 23512 11544
rect 22552 11504 23512 11532
rect 22552 11492 22558 11504
rect 23506 11492 23512 11504
rect 23564 11492 23570 11544
rect 26358 11532 26364 11544
rect 26319 11504 26364 11532
rect 26358 11492 26364 11504
rect 26416 11492 26422 11544
rect 26726 11532 26732 11544
rect 26687 11504 26732 11532
rect 26726 11492 26732 11504
rect 26784 11492 26790 11544
rect 28106 11532 28112 11544
rect 28067 11504 28112 11532
rect 28106 11492 28112 11504
rect 28164 11492 28170 11544
rect 28198 11492 28204 11544
rect 28256 11532 28262 11544
rect 28937 11535 28995 11541
rect 28937 11532 28949 11535
rect 28256 11504 28949 11532
rect 28256 11492 28262 11504
rect 28937 11501 28949 11504
rect 28983 11532 28995 11535
rect 29210 11532 29216 11544
rect 28983 11504 29216 11532
rect 28983 11501 28995 11504
rect 28937 11495 28995 11501
rect 29210 11492 29216 11504
rect 29268 11532 29274 11544
rect 29366 11532 29394 11572
rect 29854 11560 29860 11572
rect 29912 11600 29918 11612
rect 29949 11603 30007 11609
rect 29949 11600 29961 11603
rect 29912 11572 29961 11600
rect 29912 11560 29918 11572
rect 29949 11569 29961 11572
rect 29995 11569 30007 11603
rect 30317 11603 30375 11609
rect 30317 11600 30329 11603
rect 29949 11563 30007 11569
rect 30056 11572 30329 11600
rect 29268 11504 29394 11532
rect 29268 11492 29274 11504
rect 29670 11492 29676 11544
rect 29728 11532 29734 11544
rect 29765 11535 29823 11541
rect 29765 11532 29777 11535
rect 29728 11504 29777 11532
rect 29728 11492 29734 11504
rect 29765 11501 29777 11504
rect 29811 11501 29823 11535
rect 29765 11495 29823 11501
rect 30056 11476 30084 11572
rect 30317 11569 30329 11572
rect 30363 11569 30375 11603
rect 30317 11563 30375 11569
rect 30222 11532 30228 11544
rect 30183 11504 30228 11532
rect 30222 11492 30228 11504
rect 30280 11492 30286 11544
rect 12650 11464 12656 11476
rect 9856 11436 12656 11464
rect 9856 11424 9862 11436
rect 12650 11424 12656 11436
rect 12708 11424 12714 11476
rect 20654 11464 20660 11476
rect 20615 11436 20660 11464
rect 20654 11424 20660 11436
rect 20712 11424 20718 11476
rect 27462 11424 27468 11476
rect 27520 11464 27526 11476
rect 29121 11467 29179 11473
rect 29121 11464 29133 11467
rect 27520 11436 29133 11464
rect 27520 11424 27526 11436
rect 29121 11433 29133 11436
rect 29167 11464 29179 11467
rect 29578 11464 29584 11476
rect 29167 11436 29584 11464
rect 29167 11433 29179 11436
rect 29121 11427 29179 11433
rect 29578 11424 29584 11436
rect 29636 11464 29642 11476
rect 30038 11464 30044 11476
rect 29636 11436 30044 11464
rect 29636 11424 29642 11436
rect 30038 11424 30044 11436
rect 30096 11424 30102 11476
rect 1426 11396 1432 11408
rect 1387 11368 1432 11396
rect 1426 11356 1432 11368
rect 1484 11356 1490 11408
rect 6213 11399 6271 11405
rect 6213 11365 6225 11399
rect 6259 11396 6271 11399
rect 6394 11396 6400 11408
rect 6259 11368 6400 11396
rect 6259 11365 6271 11368
rect 6213 11359 6271 11365
rect 6394 11356 6400 11368
rect 6452 11356 6458 11408
rect 12742 11396 12748 11408
rect 12703 11368 12748 11396
rect 12742 11356 12748 11368
rect 12800 11356 12806 11408
rect 24334 11396 24340 11408
rect 24247 11368 24340 11396
rect 24334 11356 24340 11368
rect 24392 11396 24398 11408
rect 28658 11396 28664 11408
rect 24392 11368 28664 11396
rect 24392 11356 24398 11368
rect 28658 11356 28664 11368
rect 28716 11356 28722 11408
rect 400 11306 31680 11328
rect 400 11254 3510 11306
rect 3562 11254 3574 11306
rect 3626 11254 3638 11306
rect 3690 11254 3702 11306
rect 3754 11254 3766 11306
rect 3818 11254 31680 11306
rect 400 11232 31680 11254
rect 1334 11192 1340 11204
rect 1295 11164 1340 11192
rect 1334 11152 1340 11164
rect 1392 11152 1398 11204
rect 7682 11152 7688 11204
rect 7740 11192 7746 11204
rect 8878 11192 8884 11204
rect 7740 11164 8884 11192
rect 7740 11152 7746 11164
rect 8878 11152 8884 11164
rect 8936 11192 8942 11204
rect 8973 11195 9031 11201
rect 8973 11192 8985 11195
rect 8936 11164 8985 11192
rect 8936 11152 8942 11164
rect 8973 11161 8985 11164
rect 9019 11161 9031 11195
rect 9154 11192 9160 11204
rect 9115 11164 9160 11192
rect 8973 11155 9031 11161
rect 9154 11152 9160 11164
rect 9212 11152 9218 11204
rect 12193 11195 12251 11201
rect 12193 11161 12205 11195
rect 12239 11192 12251 11195
rect 12558 11192 12564 11204
rect 12239 11164 12564 11192
rect 12239 11161 12251 11164
rect 12193 11155 12251 11161
rect 12558 11152 12564 11164
rect 12616 11152 12622 11204
rect 12745 11195 12803 11201
rect 12745 11161 12757 11195
rect 12791 11192 12803 11195
rect 13110 11192 13116 11204
rect 12791 11164 13116 11192
rect 12791 11161 12803 11164
rect 12745 11155 12803 11161
rect 13110 11152 13116 11164
rect 13168 11192 13174 11204
rect 14950 11192 14956 11204
rect 13168 11164 14956 11192
rect 13168 11152 13174 11164
rect 14950 11152 14956 11164
rect 15008 11152 15014 11204
rect 15410 11192 15416 11204
rect 15371 11164 15416 11192
rect 15410 11152 15416 11164
rect 15468 11152 15474 11204
rect 15597 11195 15655 11201
rect 15597 11161 15609 11195
rect 15643 11192 15655 11195
rect 15686 11192 15692 11204
rect 15643 11164 15692 11192
rect 15643 11161 15655 11164
rect 15597 11155 15655 11161
rect 15686 11152 15692 11164
rect 15744 11152 15750 11204
rect 17526 11192 17532 11204
rect 17487 11164 17532 11192
rect 17526 11152 17532 11164
rect 17584 11152 17590 11204
rect 17618 11152 17624 11204
rect 17676 11192 17682 11204
rect 19829 11195 19887 11201
rect 19829 11192 19841 11195
rect 17676 11164 19841 11192
rect 17676 11152 17682 11164
rect 19829 11161 19841 11164
rect 19875 11192 19887 11195
rect 20381 11195 20439 11201
rect 20381 11192 20393 11195
rect 19875 11164 20393 11192
rect 19875 11161 19887 11164
rect 19829 11155 19887 11161
rect 20381 11161 20393 11164
rect 20427 11161 20439 11195
rect 21298 11192 21304 11204
rect 21259 11164 21304 11192
rect 20381 11155 20439 11161
rect 21298 11152 21304 11164
rect 21356 11152 21362 11204
rect 21482 11192 21488 11204
rect 21443 11164 21488 11192
rect 21482 11152 21488 11164
rect 21540 11152 21546 11204
rect 25809 11195 25867 11201
rect 25809 11161 25821 11195
rect 25855 11192 25867 11195
rect 26726 11192 26732 11204
rect 25855 11164 26732 11192
rect 25855 11161 25867 11164
rect 25809 11155 25867 11161
rect 26726 11152 26732 11164
rect 26784 11152 26790 11204
rect 29302 11152 29308 11204
rect 29360 11192 29366 11204
rect 29489 11195 29547 11201
rect 29489 11192 29501 11195
rect 29360 11164 29501 11192
rect 29360 11152 29366 11164
rect 29489 11161 29501 11164
rect 29535 11161 29547 11195
rect 29854 11192 29860 11204
rect 29815 11164 29860 11192
rect 29489 11155 29547 11161
rect 29854 11152 29860 11164
rect 29912 11152 29918 11204
rect 30038 11192 30044 11204
rect 29999 11164 30044 11192
rect 30038 11152 30044 11164
rect 30096 11152 30102 11204
rect 7590 11084 7596 11136
rect 7648 11124 7654 11136
rect 8697 11127 8755 11133
rect 8697 11124 8709 11127
rect 7648 11096 8709 11124
rect 7648 11084 7654 11096
rect 8697 11093 8709 11096
rect 8743 11124 8755 11127
rect 9706 11124 9712 11136
rect 8743 11096 9712 11124
rect 8743 11093 8755 11096
rect 8697 11087 8755 11093
rect 9706 11084 9712 11096
rect 9764 11084 9770 11136
rect 12374 11124 12380 11136
rect 12335 11096 12380 11124
rect 12374 11084 12380 11096
rect 12432 11084 12438 11136
rect 12650 11084 12656 11136
rect 12708 11124 12714 11136
rect 17434 11124 17440 11136
rect 12708 11096 17440 11124
rect 12708 11084 12714 11096
rect 17434 11084 17440 11096
rect 17492 11084 17498 11136
rect 6394 11016 6400 11068
rect 6452 11056 6458 11068
rect 6489 11059 6547 11065
rect 6489 11056 6501 11059
rect 6452 11028 6501 11056
rect 6452 11016 6458 11028
rect 6489 11025 6501 11028
rect 6535 11025 6547 11059
rect 6489 11019 6547 11025
rect 7866 11016 7872 11068
rect 7924 11056 7930 11068
rect 8881 11059 8939 11065
rect 8881 11056 8893 11059
rect 7924 11028 8893 11056
rect 7924 11016 7930 11028
rect 8881 11025 8893 11028
rect 8927 11056 8939 11059
rect 9982 11056 9988 11068
rect 8927 11028 9988 11056
rect 8927 11025 8939 11028
rect 8881 11019 8939 11025
rect 9982 11016 9988 11028
rect 10040 11016 10046 11068
rect 12558 11016 12564 11068
rect 12616 11056 12622 11068
rect 13205 11059 13263 11065
rect 13205 11056 13217 11059
rect 12616 11028 13217 11056
rect 12616 11016 12622 11028
rect 13205 11025 13217 11028
rect 13251 11025 13263 11059
rect 15686 11056 15692 11068
rect 13205 11019 13263 11025
rect 14692 11028 15692 11056
rect 2438 10988 2444 11000
rect 2399 10960 2444 10988
rect 2438 10948 2444 10960
rect 2496 10988 2502 11000
rect 3177 10991 3235 10997
rect 3177 10988 3189 10991
rect 2496 10960 3189 10988
rect 2496 10948 2502 10960
rect 3177 10957 3189 10960
rect 3223 10957 3235 10991
rect 6118 10988 6124 11000
rect 6079 10960 6124 10988
rect 3177 10951 3235 10957
rect 6118 10948 6124 10960
rect 6176 10948 6182 11000
rect 9433 10991 9491 10997
rect 9433 10988 9445 10991
rect 8252 10960 9445 10988
rect 2717 10923 2775 10929
rect 2717 10889 2729 10923
rect 2763 10889 2775 10923
rect 2717 10883 2775 10889
rect 1426 10852 1432 10864
rect 1387 10824 1432 10852
rect 1426 10812 1432 10824
rect 1484 10812 1490 10864
rect 2732 10852 2760 10883
rect 7406 10880 7412 10932
rect 7464 10880 7470 10932
rect 2990 10852 2996 10864
rect 2732 10824 2996 10852
rect 2990 10812 2996 10824
rect 3048 10812 3054 10864
rect 5658 10852 5664 10864
rect 5619 10824 5664 10852
rect 5658 10812 5664 10824
rect 5716 10812 5722 10864
rect 5934 10852 5940 10864
rect 5847 10824 5940 10852
rect 5934 10812 5940 10824
rect 5992 10852 5998 10864
rect 7424 10852 7452 10880
rect 5992 10824 7452 10852
rect 5992 10812 5998 10824
rect 7774 10812 7780 10864
rect 7832 10852 7838 10864
rect 8252 10861 8280 10960
rect 9433 10957 9445 10960
rect 9479 10988 9491 10991
rect 9893 10991 9951 10997
rect 9893 10988 9905 10991
rect 9479 10960 9905 10988
rect 9479 10957 9491 10960
rect 9433 10951 9491 10957
rect 9893 10957 9905 10960
rect 9939 10957 9951 10991
rect 9893 10951 9951 10957
rect 12009 10991 12067 10997
rect 12009 10957 12021 10991
rect 12055 10988 12067 10991
rect 13294 10988 13300 11000
rect 12055 10960 13300 10988
rect 12055 10957 12067 10960
rect 12009 10951 12067 10957
rect 13294 10948 13300 10960
rect 13352 10948 13358 11000
rect 13665 10991 13723 10997
rect 13665 10957 13677 10991
rect 13711 10957 13723 10991
rect 13665 10951 13723 10957
rect 9801 10923 9859 10929
rect 9801 10889 9813 10923
rect 9847 10920 9859 10923
rect 13680 10920 13708 10951
rect 13754 10948 13760 11000
rect 13812 10988 13818 11000
rect 14692 10997 14720 11028
rect 15686 11016 15692 11028
rect 15744 11016 15750 11068
rect 17544 11056 17572 11152
rect 17710 11124 17716 11136
rect 17671 11096 17716 11124
rect 17710 11084 17716 11096
rect 17768 11084 17774 11136
rect 17802 11084 17808 11136
rect 17860 11124 17866 11136
rect 18449 11127 18507 11133
rect 18449 11124 18461 11127
rect 17860 11096 18461 11124
rect 17860 11084 17866 11096
rect 18449 11093 18461 11096
rect 18495 11093 18507 11127
rect 18449 11087 18507 11093
rect 20841 11127 20899 11133
rect 20841 11093 20853 11127
rect 20887 11124 20899 11127
rect 21209 11127 21267 11133
rect 21209 11124 21221 11127
rect 20887 11096 21221 11124
rect 20887 11093 20899 11096
rect 20841 11087 20899 11093
rect 21209 11093 21221 11096
rect 21255 11124 21267 11127
rect 21850 11124 21856 11136
rect 21255 11096 21856 11124
rect 21255 11093 21267 11096
rect 21209 11087 21267 11093
rect 18633 11059 18691 11065
rect 18633 11056 18645 11059
rect 17544 11028 18645 11056
rect 14677 10991 14735 10997
rect 13812 10960 13857 10988
rect 13812 10948 13818 10960
rect 14677 10957 14689 10991
rect 14723 10957 14735 10991
rect 14677 10951 14735 10957
rect 14766 10948 14772 11000
rect 14824 10988 14830 11000
rect 14861 10991 14919 10997
rect 14861 10988 14873 10991
rect 14824 10960 14873 10988
rect 14824 10948 14830 10960
rect 14861 10957 14873 10960
rect 14907 10988 14919 10991
rect 15410 10988 15416 11000
rect 14907 10960 15416 10988
rect 14907 10957 14919 10960
rect 14861 10951 14919 10957
rect 15410 10948 15416 10960
rect 15468 10948 15474 11000
rect 17802 10988 17808 11000
rect 17763 10960 17808 10988
rect 17802 10948 17808 10960
rect 17860 10948 17866 11000
rect 17912 10997 17940 11028
rect 18633 11025 18645 11028
rect 18679 11025 18691 11059
rect 18633 11019 18691 11025
rect 17897 10991 17955 10997
rect 17897 10957 17909 10991
rect 17943 10957 17955 10991
rect 17897 10951 17955 10957
rect 20289 10991 20347 10997
rect 20289 10957 20301 10991
rect 20335 10988 20347 10991
rect 20856 10988 20884 11087
rect 21850 11084 21856 11096
rect 21908 11084 21914 11136
rect 25346 11084 25352 11136
rect 25404 11124 25410 11136
rect 25901 11127 25959 11133
rect 25901 11124 25913 11127
rect 25404 11096 25913 11124
rect 25404 11084 25410 11096
rect 25901 11093 25913 11096
rect 25947 11124 25959 11127
rect 26085 11127 26143 11133
rect 26085 11124 26097 11127
rect 25947 11096 26097 11124
rect 25947 11093 25959 11096
rect 25901 11087 25959 11093
rect 26085 11093 26097 11096
rect 26131 11093 26143 11127
rect 26085 11087 26143 11093
rect 26100 11056 26128 11087
rect 27002 11056 27008 11068
rect 26100 11028 27008 11056
rect 27002 11016 27008 11028
rect 27060 11056 27066 11068
rect 27373 11059 27431 11065
rect 27373 11056 27385 11059
rect 27060 11028 27385 11056
rect 27060 11016 27066 11028
rect 27373 11025 27385 11028
rect 27419 11056 27431 11059
rect 28106 11056 28112 11068
rect 27419 11028 28112 11056
rect 27419 11025 27431 11028
rect 27373 11019 27431 11025
rect 28106 11016 28112 11028
rect 28164 11016 28170 11068
rect 29118 11016 29124 11068
rect 29176 11056 29182 11068
rect 29302 11056 29308 11068
rect 29176 11028 29308 11056
rect 29176 11016 29182 11028
rect 29302 11016 29308 11028
rect 29360 11016 29366 11068
rect 20335 10960 20884 10988
rect 20335 10957 20347 10960
rect 20289 10951 20347 10957
rect 24886 10948 24892 11000
rect 24944 10988 24950 11000
rect 26634 10988 26640 11000
rect 24944 10960 26640 10988
rect 24944 10948 24950 10960
rect 26634 10948 26640 10960
rect 26692 10988 26698 11000
rect 26913 10991 26971 10997
rect 26913 10988 26925 10991
rect 26692 10960 26925 10988
rect 26692 10948 26698 10960
rect 26913 10957 26925 10960
rect 26959 10957 26971 10991
rect 27094 10988 27100 11000
rect 27055 10960 27100 10988
rect 26913 10951 26971 10957
rect 27094 10948 27100 10960
rect 27152 10948 27158 11000
rect 27462 10988 27468 11000
rect 27423 10960 27468 10988
rect 27462 10948 27468 10960
rect 27520 10948 27526 11000
rect 28750 10948 28756 11000
rect 28808 10988 28814 11000
rect 29670 10988 29676 11000
rect 28808 10960 29676 10988
rect 28808 10948 28814 10960
rect 29670 10948 29676 10960
rect 29728 10948 29734 11000
rect 9847 10892 10212 10920
rect 9847 10889 9859 10892
rect 9801 10883 9859 10889
rect 10184 10864 10212 10892
rect 12484 10892 13708 10920
rect 15229 10923 15287 10929
rect 8237 10855 8295 10861
rect 8237 10852 8249 10855
rect 7832 10824 8249 10852
rect 7832 10812 7838 10824
rect 8237 10821 8249 10824
rect 8283 10821 8295 10855
rect 10166 10852 10172 10864
rect 10127 10824 10172 10852
rect 8237 10815 8295 10821
rect 10166 10812 10172 10824
rect 10224 10812 10230 10864
rect 10258 10812 10264 10864
rect 10316 10852 10322 10864
rect 12484 10861 12512 10892
rect 15229 10889 15241 10923
rect 15275 10920 15287 10923
rect 16054 10920 16060 10932
rect 15275 10892 16060 10920
rect 15275 10889 15287 10892
rect 15229 10883 15287 10889
rect 12469 10855 12527 10861
rect 12469 10852 12481 10855
rect 10316 10824 12481 10852
rect 10316 10812 10322 10824
rect 12469 10821 12481 10824
rect 12515 10821 12527 10855
rect 12469 10815 12527 10821
rect 13570 10812 13576 10864
rect 13628 10852 13634 10864
rect 14585 10855 14643 10861
rect 14585 10852 14597 10855
rect 13628 10824 14597 10852
rect 13628 10812 13634 10824
rect 14585 10821 14597 10824
rect 14631 10852 14643 10855
rect 15244 10852 15272 10883
rect 16054 10880 16060 10892
rect 16112 10880 16118 10932
rect 18357 10923 18415 10929
rect 18357 10889 18369 10923
rect 18403 10920 18415 10923
rect 18722 10920 18728 10932
rect 18403 10892 18728 10920
rect 18403 10889 18415 10892
rect 18357 10883 18415 10889
rect 18722 10880 18728 10892
rect 18780 10880 18786 10932
rect 20013 10923 20071 10929
rect 20013 10889 20025 10923
rect 20059 10920 20071 10923
rect 20105 10923 20163 10929
rect 20105 10920 20117 10923
rect 20059 10892 20117 10920
rect 20059 10889 20071 10892
rect 20013 10883 20071 10889
rect 20105 10889 20117 10892
rect 20151 10920 20163 10923
rect 21942 10920 21948 10932
rect 20151 10892 21948 10920
rect 20151 10889 20163 10892
rect 20105 10883 20163 10889
rect 21942 10880 21948 10892
rect 22000 10880 22006 10932
rect 26269 10923 26327 10929
rect 26269 10920 26281 10923
rect 23248 10892 26281 10920
rect 23248 10864 23276 10892
rect 26269 10889 26281 10892
rect 26315 10920 26327 10923
rect 27186 10920 27192 10932
rect 26315 10892 27192 10920
rect 26315 10889 26327 10892
rect 26269 10883 26327 10889
rect 27186 10880 27192 10892
rect 27244 10880 27250 10932
rect 30222 10920 30228 10932
rect 29320 10892 30228 10920
rect 14631 10824 15272 10852
rect 14631 10821 14643 10824
rect 14585 10815 14643 10821
rect 19918 10812 19924 10864
rect 19976 10852 19982 10864
rect 20286 10852 20292 10864
rect 19976 10824 20292 10852
rect 19976 10812 19982 10824
rect 20286 10812 20292 10824
rect 20344 10852 20350 10864
rect 20933 10855 20991 10861
rect 20933 10852 20945 10855
rect 20344 10824 20945 10852
rect 20344 10812 20350 10824
rect 20933 10821 20945 10824
rect 20979 10852 20991 10855
rect 21666 10852 21672 10864
rect 20979 10824 21672 10852
rect 20979 10821 20991 10824
rect 20933 10815 20991 10821
rect 21666 10812 21672 10824
rect 21724 10852 21730 10864
rect 23230 10852 23236 10864
rect 21724 10824 23236 10852
rect 21724 10812 21730 10824
rect 23230 10812 23236 10824
rect 23288 10812 23294 10864
rect 25625 10855 25683 10861
rect 25625 10821 25637 10855
rect 25671 10852 25683 10855
rect 26910 10852 26916 10864
rect 25671 10824 26916 10852
rect 25671 10821 25683 10824
rect 25625 10815 25683 10821
rect 26910 10812 26916 10824
rect 26968 10852 26974 10864
rect 27462 10852 27468 10864
rect 26968 10824 27468 10852
rect 26968 10812 26974 10824
rect 27462 10812 27468 10824
rect 27520 10812 27526 10864
rect 29118 10812 29124 10864
rect 29176 10852 29182 10864
rect 29320 10861 29348 10892
rect 30222 10880 30228 10892
rect 30280 10880 30286 10932
rect 29305 10855 29363 10861
rect 29305 10852 29317 10855
rect 29176 10824 29317 10852
rect 29176 10812 29182 10824
rect 29305 10821 29317 10824
rect 29351 10821 29363 10855
rect 29305 10815 29363 10821
rect 400 10762 31680 10784
rect 400 10710 18870 10762
rect 18922 10710 18934 10762
rect 18986 10710 18998 10762
rect 19050 10710 19062 10762
rect 19114 10710 19126 10762
rect 19178 10710 31680 10762
rect 400 10688 31680 10710
rect 12558 10608 12564 10660
rect 12616 10648 12622 10660
rect 12653 10651 12711 10657
rect 12653 10648 12665 10651
rect 12616 10620 12665 10648
rect 12616 10608 12622 10620
rect 12653 10617 12665 10620
rect 12699 10617 12711 10651
rect 13110 10648 13116 10660
rect 13071 10620 13116 10648
rect 12653 10611 12711 10617
rect 13110 10608 13116 10620
rect 13168 10608 13174 10660
rect 14858 10608 14864 10660
rect 14916 10648 14922 10660
rect 18446 10648 18452 10660
rect 14916 10620 18452 10648
rect 14916 10608 14922 10620
rect 18446 10608 18452 10620
rect 18504 10608 18510 10660
rect 19274 10608 19280 10660
rect 19332 10648 19338 10660
rect 19369 10651 19427 10657
rect 19369 10648 19381 10651
rect 19332 10620 19381 10648
rect 19332 10608 19338 10620
rect 19369 10617 19381 10620
rect 19415 10617 19427 10651
rect 19369 10611 19427 10617
rect 26545 10651 26603 10657
rect 26545 10617 26557 10651
rect 26591 10648 26603 10651
rect 26726 10648 26732 10660
rect 26591 10620 26732 10648
rect 26591 10617 26603 10620
rect 26545 10611 26603 10617
rect 26726 10608 26732 10620
rect 26784 10608 26790 10660
rect 26913 10651 26971 10657
rect 26913 10617 26925 10651
rect 26959 10648 26971 10651
rect 27094 10648 27100 10660
rect 26959 10620 27100 10648
rect 26959 10617 26971 10620
rect 26913 10611 26971 10617
rect 27094 10608 27100 10620
rect 27152 10608 27158 10660
rect 28014 10608 28020 10660
rect 28072 10648 28078 10660
rect 28658 10648 28664 10660
rect 28072 10620 28664 10648
rect 28072 10608 28078 10620
rect 28658 10608 28664 10620
rect 28716 10648 28722 10660
rect 28753 10651 28811 10657
rect 28753 10648 28765 10651
rect 28716 10620 28765 10648
rect 28716 10608 28722 10620
rect 28753 10617 28765 10620
rect 28799 10617 28811 10651
rect 28753 10611 28811 10617
rect 6394 10540 6400 10592
rect 6452 10580 6458 10592
rect 6857 10583 6915 10589
rect 6857 10580 6869 10583
rect 6452 10552 6869 10580
rect 6452 10540 6458 10552
rect 6857 10549 6869 10552
rect 6903 10580 6915 10583
rect 7038 10580 7044 10592
rect 6903 10552 7044 10580
rect 6903 10549 6915 10552
rect 6857 10543 6915 10549
rect 7038 10540 7044 10552
rect 7096 10540 7102 10592
rect 12929 10583 12987 10589
rect 12929 10549 12941 10583
rect 12975 10580 12987 10583
rect 13665 10583 13723 10589
rect 13665 10580 13677 10583
rect 12975 10552 13677 10580
rect 12975 10549 12987 10552
rect 12929 10543 12987 10549
rect 13665 10549 13677 10552
rect 13711 10580 13723 10583
rect 13754 10580 13760 10592
rect 13711 10552 13760 10580
rect 13711 10549 13723 10552
rect 13665 10543 13723 10549
rect 13754 10540 13760 10552
rect 13812 10540 13818 10592
rect 16238 10580 16244 10592
rect 16151 10552 16244 10580
rect 16238 10540 16244 10552
rect 16296 10580 16302 10592
rect 17618 10580 17624 10592
rect 16296 10552 17624 10580
rect 16296 10540 16302 10552
rect 17618 10540 17624 10552
rect 17676 10540 17682 10592
rect 17897 10583 17955 10589
rect 17897 10549 17909 10583
rect 17943 10580 17955 10583
rect 26634 10580 26640 10592
rect 17943 10552 18860 10580
rect 26595 10552 26640 10580
rect 17943 10549 17955 10552
rect 17897 10543 17955 10549
rect 18832 10524 18860 10552
rect 26634 10540 26640 10552
rect 26692 10540 26698 10592
rect 27112 10580 27140 10608
rect 28198 10580 28204 10592
rect 27112 10552 28204 10580
rect 28198 10540 28204 10552
rect 28256 10540 28262 10592
rect 2165 10515 2223 10521
rect 2165 10481 2177 10515
rect 2211 10512 2223 10515
rect 2990 10512 2996 10524
rect 2211 10484 2996 10512
rect 2211 10481 2223 10484
rect 2165 10475 2223 10481
rect 2990 10472 2996 10484
rect 3048 10472 3054 10524
rect 3821 10515 3879 10521
rect 3821 10481 3833 10515
rect 3867 10512 3879 10515
rect 4462 10512 4468 10524
rect 3867 10484 4468 10512
rect 3867 10481 3879 10484
rect 3821 10475 3879 10481
rect 4462 10472 4468 10484
rect 4520 10472 4526 10524
rect 7501 10515 7559 10521
rect 7501 10512 7513 10515
rect 7424 10484 7513 10512
rect 7424 10456 7452 10484
rect 7501 10481 7513 10484
rect 7547 10481 7559 10515
rect 7866 10512 7872 10524
rect 7827 10484 7872 10512
rect 7501 10475 7559 10481
rect 7866 10472 7872 10484
rect 7924 10472 7930 10524
rect 12561 10515 12619 10521
rect 12561 10481 12573 10515
rect 12607 10512 12619 10515
rect 12742 10512 12748 10524
rect 12607 10484 12748 10512
rect 12607 10481 12619 10484
rect 12561 10475 12619 10481
rect 12742 10472 12748 10484
rect 12800 10472 12806 10524
rect 13570 10512 13576 10524
rect 13531 10484 13576 10512
rect 13570 10472 13576 10484
rect 13628 10472 13634 10524
rect 14585 10515 14643 10521
rect 14585 10481 14597 10515
rect 14631 10512 14643 10515
rect 14674 10512 14680 10524
rect 14631 10484 14680 10512
rect 14631 10481 14643 10484
rect 14585 10475 14643 10481
rect 14674 10472 14680 10484
rect 14732 10472 14738 10524
rect 14766 10472 14772 10524
rect 14824 10512 14830 10524
rect 14824 10484 14869 10512
rect 14824 10472 14830 10484
rect 16330 10472 16336 10524
rect 16388 10512 16394 10524
rect 16388 10484 16433 10512
rect 16388 10472 16394 10484
rect 17710 10472 17716 10524
rect 17768 10512 17774 10524
rect 18630 10512 18636 10524
rect 17768 10484 18636 10512
rect 17768 10472 17774 10484
rect 18630 10472 18636 10484
rect 18688 10512 18694 10524
rect 18725 10515 18783 10521
rect 18725 10512 18737 10515
rect 18688 10484 18737 10512
rect 18688 10472 18694 10484
rect 18725 10481 18737 10484
rect 18771 10481 18783 10515
rect 18725 10475 18783 10481
rect 18814 10472 18820 10524
rect 18872 10512 18878 10524
rect 19093 10515 19151 10521
rect 19093 10512 19105 10515
rect 18872 10484 19105 10512
rect 18872 10472 18878 10484
rect 19093 10481 19105 10484
rect 19139 10481 19151 10515
rect 26082 10512 26088 10524
rect 25995 10484 26088 10512
rect 19093 10475 19151 10481
rect 26082 10472 26088 10484
rect 26140 10512 26146 10524
rect 29762 10512 29768 10524
rect 26140 10484 29768 10512
rect 26140 10472 26146 10484
rect 29762 10472 29768 10484
rect 29820 10472 29826 10524
rect 1978 10404 1984 10456
rect 2036 10444 2042 10456
rect 3729 10447 3787 10453
rect 3729 10444 3741 10447
rect 2036 10416 3741 10444
rect 2036 10404 2042 10416
rect 3729 10413 3741 10416
rect 3775 10444 3787 10447
rect 4094 10444 4100 10456
rect 3775 10416 4100 10444
rect 3775 10413 3787 10416
rect 3729 10407 3787 10413
rect 4094 10404 4100 10416
rect 4152 10404 4158 10456
rect 7406 10404 7412 10456
rect 7464 10404 7470 10456
rect 7590 10444 7596 10456
rect 7551 10416 7596 10444
rect 7590 10404 7596 10416
rect 7648 10404 7654 10456
rect 7774 10444 7780 10456
rect 7735 10416 7780 10444
rect 7774 10404 7780 10416
rect 7832 10404 7838 10456
rect 18446 10404 18452 10456
rect 18504 10444 18510 10456
rect 18541 10447 18599 10453
rect 18541 10444 18553 10447
rect 18504 10416 18553 10444
rect 18504 10404 18510 10416
rect 18541 10413 18553 10416
rect 18587 10413 18599 10447
rect 18541 10407 18599 10413
rect 13294 10336 13300 10388
rect 13352 10376 13358 10388
rect 18556 10376 18584 10407
rect 18906 10404 18912 10456
rect 18964 10444 18970 10456
rect 19001 10447 19059 10453
rect 19001 10444 19013 10447
rect 18964 10416 19013 10444
rect 18964 10404 18970 10416
rect 19001 10413 19013 10416
rect 19047 10444 19059 10447
rect 19458 10444 19464 10456
rect 19047 10416 19464 10444
rect 19047 10413 19059 10416
rect 19001 10407 19059 10413
rect 19458 10404 19464 10416
rect 19516 10404 19522 10456
rect 22954 10444 22960 10456
rect 22915 10416 22960 10444
rect 22954 10404 22960 10416
rect 23012 10404 23018 10456
rect 23782 10404 23788 10456
rect 23840 10444 23846 10456
rect 24334 10444 24340 10456
rect 23840 10416 24340 10444
rect 23840 10404 23846 10416
rect 24334 10404 24340 10416
rect 24392 10404 24398 10456
rect 26358 10444 26364 10456
rect 24444 10416 26364 10444
rect 20102 10376 20108 10388
rect 13352 10348 16560 10376
rect 18556 10348 20108 10376
rect 13352 10336 13358 10348
rect 3910 10268 3916 10320
rect 3968 10308 3974 10320
rect 4005 10311 4063 10317
rect 4005 10308 4017 10311
rect 3968 10280 4017 10308
rect 3968 10268 3974 10280
rect 4005 10277 4017 10280
rect 4051 10308 4063 10311
rect 4554 10308 4560 10320
rect 4051 10280 4560 10308
rect 4051 10277 4063 10280
rect 4005 10271 4063 10277
rect 4554 10268 4560 10280
rect 4612 10268 4618 10320
rect 6118 10268 6124 10320
rect 6176 10308 6182 10320
rect 6213 10311 6271 10317
rect 6213 10308 6225 10311
rect 6176 10280 6225 10308
rect 6176 10268 6182 10280
rect 6213 10277 6225 10280
rect 6259 10308 6271 10311
rect 8142 10308 8148 10320
rect 6259 10280 8148 10308
rect 6259 10277 6271 10280
rect 6213 10271 6271 10277
rect 8142 10268 8148 10280
rect 8200 10268 8206 10320
rect 8970 10308 8976 10320
rect 8931 10280 8976 10308
rect 8970 10268 8976 10280
rect 9028 10268 9034 10320
rect 14122 10268 14128 10320
rect 14180 10308 14186 10320
rect 14858 10308 14864 10320
rect 14180 10280 14864 10308
rect 14180 10268 14186 10280
rect 14858 10268 14864 10280
rect 14916 10268 14922 10320
rect 16054 10308 16060 10320
rect 16015 10280 16060 10308
rect 16054 10268 16060 10280
rect 16112 10268 16118 10320
rect 16532 10317 16560 10348
rect 20102 10336 20108 10348
rect 20160 10336 20166 10388
rect 24242 10336 24248 10388
rect 24300 10376 24306 10388
rect 24444 10376 24472 10416
rect 26358 10404 26364 10416
rect 26416 10444 26422 10456
rect 27005 10447 27063 10453
rect 27005 10444 27017 10447
rect 26416 10416 27017 10444
rect 26416 10404 26422 10416
rect 27005 10413 27017 10416
rect 27051 10413 27063 10447
rect 27005 10407 27063 10413
rect 24300 10348 24472 10376
rect 24300 10336 24306 10348
rect 25622 10336 25628 10388
rect 25680 10376 25686 10388
rect 25680 10348 28704 10376
rect 25680 10336 25686 10348
rect 16517 10311 16575 10317
rect 16517 10277 16529 10311
rect 16563 10308 16575 10311
rect 16606 10308 16612 10320
rect 16563 10280 16612 10308
rect 16563 10277 16575 10280
rect 16517 10271 16575 10277
rect 16606 10268 16612 10280
rect 16664 10268 16670 10320
rect 17434 10308 17440 10320
rect 17395 10280 17440 10308
rect 17434 10268 17440 10280
rect 17492 10268 17498 10320
rect 18354 10308 18360 10320
rect 18315 10280 18360 10308
rect 18354 10268 18360 10280
rect 18412 10268 18418 10320
rect 23138 10308 23144 10320
rect 23099 10280 23144 10308
rect 23138 10268 23144 10280
rect 23196 10268 23202 10320
rect 25898 10308 25904 10320
rect 25859 10280 25904 10308
rect 25898 10268 25904 10280
rect 25956 10268 25962 10320
rect 28676 10317 28704 10348
rect 28661 10311 28719 10317
rect 28661 10277 28673 10311
rect 28707 10308 28719 10311
rect 29670 10308 29676 10320
rect 28707 10280 29676 10308
rect 28707 10277 28719 10280
rect 28661 10271 28719 10277
rect 29670 10268 29676 10280
rect 29728 10268 29734 10320
rect 400 10218 31680 10240
rect 400 10166 3510 10218
rect 3562 10166 3574 10218
rect 3626 10166 3638 10218
rect 3690 10166 3702 10218
rect 3754 10166 3766 10218
rect 3818 10166 31680 10218
rect 400 10144 31680 10166
rect 1978 10104 1984 10116
rect 1939 10076 1984 10104
rect 1978 10064 1984 10076
rect 2036 10064 2042 10116
rect 4462 10104 4468 10116
rect 4423 10076 4468 10104
rect 4462 10064 4468 10076
rect 4520 10064 4526 10116
rect 4554 10064 4560 10116
rect 4612 10104 4618 10116
rect 7038 10104 7044 10116
rect 4612 10076 4657 10104
rect 6999 10076 7044 10104
rect 4612 10064 4618 10076
rect 7038 10064 7044 10076
rect 7096 10064 7102 10116
rect 7501 10107 7559 10113
rect 7501 10073 7513 10107
rect 7547 10104 7559 10107
rect 7590 10104 7596 10116
rect 7547 10076 7596 10104
rect 7547 10073 7559 10076
rect 7501 10067 7559 10073
rect 7590 10064 7596 10076
rect 7648 10064 7654 10116
rect 8697 10107 8755 10113
rect 8697 10073 8709 10107
rect 8743 10104 8755 10107
rect 8786 10104 8792 10116
rect 8743 10076 8792 10104
rect 8743 10073 8755 10076
rect 8697 10067 8755 10073
rect 8786 10064 8792 10076
rect 8844 10104 8850 10116
rect 9522 10104 9528 10116
rect 8844 10076 9528 10104
rect 8844 10064 8850 10076
rect 9522 10064 9528 10076
rect 9580 10064 9586 10116
rect 13573 10107 13631 10113
rect 13573 10073 13585 10107
rect 13619 10104 13631 10107
rect 13754 10104 13760 10116
rect 13619 10076 13760 10104
rect 13619 10073 13631 10076
rect 13573 10067 13631 10073
rect 13754 10064 13760 10076
rect 13812 10064 13818 10116
rect 14122 10104 14128 10116
rect 14083 10076 14128 10104
rect 14122 10064 14128 10076
rect 14180 10064 14186 10116
rect 14490 10104 14496 10116
rect 14451 10076 14496 10104
rect 14490 10064 14496 10076
rect 14548 10064 14554 10116
rect 14766 10064 14772 10116
rect 14824 10104 14830 10116
rect 15229 10107 15287 10113
rect 15229 10104 15241 10107
rect 14824 10076 15241 10104
rect 14824 10064 14830 10076
rect 15229 10073 15241 10076
rect 15275 10073 15287 10107
rect 16054 10104 16060 10116
rect 16015 10076 16060 10104
rect 15229 10067 15287 10073
rect 7317 10039 7375 10045
rect 7317 10005 7329 10039
rect 7363 10036 7375 10039
rect 7866 10036 7872 10048
rect 7363 10008 7872 10036
rect 7363 10005 7375 10008
rect 7317 9999 7375 10005
rect 7866 9996 7872 10008
rect 7924 9996 7930 10048
rect 2070 9968 2076 9980
rect 2031 9940 2076 9968
rect 2070 9928 2076 9940
rect 2128 9928 2134 9980
rect 4094 9968 4100 9980
rect 4055 9940 4100 9968
rect 4094 9928 4100 9940
rect 4152 9968 4158 9980
rect 4189 9971 4247 9977
rect 4189 9968 4201 9971
rect 4152 9940 4201 9968
rect 4152 9928 4158 9940
rect 4189 9937 4201 9940
rect 4235 9937 4247 9971
rect 4189 9931 4247 9937
rect 7406 9928 7412 9980
rect 7464 9968 7470 9980
rect 7590 9968 7596 9980
rect 7464 9940 7596 9968
rect 7464 9928 7470 9940
rect 7590 9928 7596 9940
rect 7648 9928 7654 9980
rect 8142 9928 8148 9980
rect 8200 9968 8206 9980
rect 8786 9968 8792 9980
rect 8200 9940 8792 9968
rect 8200 9928 8206 9940
rect 8786 9928 8792 9940
rect 8844 9928 8850 9980
rect 13389 9971 13447 9977
rect 13389 9937 13401 9971
rect 13435 9968 13447 9971
rect 13570 9968 13576 9980
rect 13435 9940 13576 9968
rect 13435 9937 13447 9940
rect 13389 9931 13447 9937
rect 13570 9928 13576 9940
rect 13628 9928 13634 9980
rect 15244 9968 15272 10067
rect 16054 10064 16060 10076
rect 16112 10064 16118 10116
rect 16238 10104 16244 10116
rect 16199 10076 16244 10104
rect 16238 10064 16244 10076
rect 16296 10064 16302 10116
rect 16606 10104 16612 10116
rect 16567 10076 16612 10104
rect 16606 10064 16612 10076
rect 16664 10064 16670 10116
rect 17434 10064 17440 10116
rect 17492 10104 17498 10116
rect 17621 10107 17679 10113
rect 17621 10104 17633 10107
rect 17492 10076 17633 10104
rect 17492 10064 17498 10076
rect 17621 10073 17633 10076
rect 17667 10073 17679 10107
rect 18354 10104 18360 10116
rect 18315 10076 18360 10104
rect 17621 10067 17679 10073
rect 18354 10064 18360 10076
rect 18412 10064 18418 10116
rect 18909 10107 18967 10113
rect 18909 10073 18921 10107
rect 18955 10104 18967 10107
rect 19918 10104 19924 10116
rect 18955 10076 19924 10104
rect 18955 10073 18967 10076
rect 18909 10067 18967 10073
rect 19918 10064 19924 10076
rect 19976 10064 19982 10116
rect 22773 10107 22831 10113
rect 22773 10073 22785 10107
rect 22819 10104 22831 10107
rect 24610 10104 24616 10116
rect 22819 10076 24616 10104
rect 22819 10073 22831 10076
rect 22773 10067 22831 10073
rect 24610 10064 24616 10076
rect 24668 10104 24674 10116
rect 25625 10107 25683 10113
rect 25625 10104 25637 10107
rect 24668 10076 25637 10104
rect 24668 10064 24674 10076
rect 25625 10073 25637 10076
rect 25671 10104 25683 10107
rect 26082 10104 26088 10116
rect 25671 10076 26088 10104
rect 25671 10073 25683 10076
rect 25625 10067 25683 10073
rect 26082 10064 26088 10076
rect 26140 10064 26146 10116
rect 28658 10104 28664 10116
rect 28619 10076 28664 10104
rect 28658 10064 28664 10076
rect 28716 10064 28722 10116
rect 16330 9996 16336 10048
rect 16388 10036 16394 10048
rect 16517 10039 16575 10045
rect 16517 10036 16529 10039
rect 16388 10008 16529 10036
rect 16388 9996 16394 10008
rect 16517 10005 16529 10008
rect 16563 10036 16575 10039
rect 17526 10036 17532 10048
rect 16563 10008 17532 10036
rect 16563 10005 16575 10008
rect 16517 9999 16575 10005
rect 17526 9996 17532 10008
rect 17584 9996 17590 10048
rect 17069 9971 17127 9977
rect 17069 9968 17081 9971
rect 15244 9940 17081 9968
rect 17069 9937 17081 9940
rect 17115 9968 17127 9971
rect 18372 9968 18400 10064
rect 25346 9996 25352 10048
rect 25404 10036 25410 10048
rect 26174 10036 26180 10048
rect 25404 10008 26180 10036
rect 25404 9996 25410 10008
rect 26174 9996 26180 10008
rect 26232 9996 26238 10048
rect 29578 10036 29584 10048
rect 29366 10008 29584 10036
rect 19274 9968 19280 9980
rect 17115 9940 17572 9968
rect 18372 9940 19280 9968
rect 17115 9937 17127 9940
rect 17069 9931 17127 9937
rect 7498 9860 7504 9912
rect 7556 9900 7562 9912
rect 8418 9900 8424 9912
rect 7556 9872 8424 9900
rect 7556 9860 7562 9872
rect 8418 9860 8424 9872
rect 8476 9860 8482 9912
rect 14309 9903 14367 9909
rect 14309 9869 14321 9903
rect 14355 9900 14367 9903
rect 14769 9903 14827 9909
rect 14355 9872 14720 9900
rect 14355 9869 14367 9872
rect 14309 9863 14367 9869
rect 1797 9835 1855 9841
rect 1797 9801 1809 9835
rect 1843 9832 1855 9835
rect 2346 9832 2352 9844
rect 1843 9804 2352 9832
rect 1843 9801 1855 9804
rect 1797 9795 1855 9801
rect 2346 9792 2352 9804
rect 2404 9792 2410 9844
rect 2990 9792 2996 9844
rect 3048 9792 3054 9844
rect 7774 9832 7780 9844
rect 6872 9804 7780 9832
rect 5658 9724 5664 9776
rect 5716 9764 5722 9776
rect 6872 9773 6900 9804
rect 7774 9792 7780 9804
rect 7832 9792 7838 9844
rect 8329 9835 8387 9841
rect 8329 9801 8341 9835
rect 8375 9832 8387 9835
rect 9065 9835 9123 9841
rect 9065 9832 9077 9835
rect 8375 9804 9077 9832
rect 8375 9801 8387 9804
rect 8329 9795 8387 9801
rect 9065 9801 9077 9804
rect 9111 9832 9123 9835
rect 9338 9832 9344 9844
rect 9111 9804 9344 9832
rect 9111 9801 9123 9804
rect 9065 9795 9123 9801
rect 9338 9792 9344 9804
rect 9396 9792 9402 9844
rect 9522 9792 9528 9844
rect 9580 9792 9586 9844
rect 10810 9832 10816 9844
rect 10771 9804 10816 9832
rect 10810 9792 10816 9804
rect 10868 9792 10874 9844
rect 14490 9792 14496 9844
rect 14548 9832 14554 9844
rect 14585 9835 14643 9841
rect 14585 9832 14597 9835
rect 14548 9804 14597 9832
rect 14548 9792 14554 9804
rect 14585 9801 14597 9804
rect 14631 9801 14643 9835
rect 14692 9832 14720 9872
rect 14769 9869 14781 9903
rect 14815 9900 14827 9903
rect 15413 9903 15471 9909
rect 15413 9900 15425 9903
rect 14815 9872 15425 9900
rect 14815 9869 14827 9872
rect 14769 9863 14827 9869
rect 15413 9869 15425 9872
rect 15459 9900 15471 9903
rect 15870 9900 15876 9912
rect 15459 9872 15876 9900
rect 15459 9869 15471 9872
rect 15413 9863 15471 9869
rect 15870 9860 15876 9872
rect 15928 9860 15934 9912
rect 15962 9860 15968 9912
rect 16020 9900 16026 9912
rect 17544 9909 17572 9940
rect 19274 9928 19280 9940
rect 19332 9968 19338 9980
rect 19369 9971 19427 9977
rect 19369 9968 19381 9971
rect 19332 9940 19381 9968
rect 19332 9928 19338 9940
rect 19369 9937 19381 9940
rect 19415 9937 19427 9971
rect 19369 9931 19427 9937
rect 20378 9928 20384 9980
rect 20436 9968 20442 9980
rect 22313 9971 22371 9977
rect 22313 9968 22325 9971
rect 20436 9940 22325 9968
rect 20436 9928 20442 9940
rect 22313 9937 22325 9940
rect 22359 9968 22371 9971
rect 26545 9971 26603 9977
rect 26545 9968 26557 9971
rect 22359 9940 23874 9968
rect 22359 9937 22371 9940
rect 22313 9931 22371 9937
rect 16885 9903 16943 9909
rect 16885 9900 16897 9903
rect 16020 9872 16897 9900
rect 16020 9860 16026 9872
rect 16885 9869 16897 9872
rect 16931 9900 16943 9903
rect 17345 9903 17403 9909
rect 17345 9900 17357 9903
rect 16931 9872 17357 9900
rect 16931 9869 16943 9872
rect 16885 9863 16943 9869
rect 17345 9869 17357 9872
rect 17391 9869 17403 9903
rect 17345 9863 17403 9869
rect 17529 9903 17587 9909
rect 17529 9869 17541 9903
rect 17575 9869 17587 9903
rect 17529 9863 17587 9869
rect 19001 9903 19059 9909
rect 19001 9869 19013 9903
rect 19047 9900 19059 9903
rect 19090 9900 19096 9912
rect 19047 9872 19096 9900
rect 19047 9869 19059 9872
rect 19001 9863 19059 9869
rect 19090 9860 19096 9872
rect 19148 9900 19154 9912
rect 19458 9900 19464 9912
rect 19148 9872 19464 9900
rect 19148 9860 19154 9872
rect 19458 9860 19464 9872
rect 19516 9860 19522 9912
rect 23046 9860 23052 9912
rect 23104 9900 23110 9912
rect 23414 9900 23420 9912
rect 23104 9872 23420 9900
rect 23104 9860 23110 9872
rect 23414 9860 23420 9872
rect 23472 9860 23478 9912
rect 23601 9903 23659 9909
rect 23601 9869 23613 9903
rect 23647 9869 23659 9903
rect 23601 9863 23659 9869
rect 23846 9900 23874 9940
rect 25732 9940 26557 9968
rect 25732 9912 25760 9940
rect 26545 9937 26557 9940
rect 26591 9937 26603 9971
rect 26545 9931 26603 9937
rect 28290 9928 28296 9980
rect 28348 9968 28354 9980
rect 28385 9971 28443 9977
rect 28385 9968 28397 9971
rect 28348 9940 28397 9968
rect 28348 9928 28354 9940
rect 28385 9937 28397 9940
rect 28431 9968 28443 9971
rect 29366 9968 29394 10008
rect 29578 9996 29584 10008
rect 29636 9996 29642 10048
rect 28431 9940 29394 9968
rect 28431 9937 28443 9940
rect 28385 9931 28443 9937
rect 23969 9903 24027 9909
rect 23969 9900 23981 9903
rect 23846 9872 23981 9900
rect 15042 9832 15048 9844
rect 14692 9804 15048 9832
rect 14585 9795 14643 9801
rect 6857 9767 6915 9773
rect 6857 9764 6869 9767
rect 5716 9736 6869 9764
rect 5716 9724 5722 9736
rect 6857 9733 6869 9736
rect 6903 9733 6915 9767
rect 9540 9764 9568 9792
rect 11546 9764 11552 9776
rect 9540 9736 11552 9764
rect 6857 9727 6915 9733
rect 11546 9724 11552 9736
rect 11604 9724 11610 9776
rect 14600 9764 14628 9795
rect 15042 9792 15048 9804
rect 15100 9832 15106 9844
rect 15137 9835 15195 9841
rect 15137 9832 15149 9835
rect 15100 9804 15149 9832
rect 15100 9792 15106 9804
rect 15137 9801 15149 9804
rect 15183 9801 15195 9835
rect 15137 9795 15195 9801
rect 18173 9835 18231 9841
rect 18173 9801 18185 9835
rect 18219 9832 18231 9835
rect 18725 9835 18783 9841
rect 18725 9832 18737 9835
rect 18219 9804 18737 9832
rect 18219 9801 18231 9804
rect 18173 9795 18231 9801
rect 18725 9801 18737 9804
rect 18771 9832 18783 9835
rect 18906 9832 18912 9844
rect 18771 9804 18912 9832
rect 18771 9801 18783 9804
rect 18725 9795 18783 9801
rect 18906 9792 18912 9804
rect 18964 9832 18970 9844
rect 18964 9804 19136 9832
rect 18964 9792 18970 9804
rect 14766 9764 14772 9776
rect 14600 9736 14772 9764
rect 14766 9724 14772 9736
rect 14824 9724 14830 9776
rect 18354 9724 18360 9776
rect 18412 9764 18418 9776
rect 18449 9767 18507 9773
rect 18449 9764 18461 9767
rect 18412 9736 18461 9764
rect 18412 9724 18418 9736
rect 18449 9733 18461 9736
rect 18495 9733 18507 9767
rect 19108 9764 19136 9804
rect 19918 9792 19924 9844
rect 19976 9792 19982 9844
rect 22589 9835 22647 9841
rect 22589 9801 22601 9835
rect 22635 9832 22647 9835
rect 22862 9832 22868 9844
rect 22635 9804 22868 9832
rect 22635 9801 22647 9804
rect 22589 9795 22647 9801
rect 22862 9792 22868 9804
rect 22920 9832 22926 9844
rect 22957 9835 23015 9841
rect 22957 9832 22969 9835
rect 22920 9804 22969 9832
rect 22920 9792 22926 9804
rect 22957 9801 22969 9804
rect 23003 9801 23015 9835
rect 22957 9795 23015 9801
rect 23138 9792 23144 9844
rect 23196 9832 23202 9844
rect 23616 9832 23644 9863
rect 23196 9804 23644 9832
rect 23196 9792 23202 9804
rect 21117 9767 21175 9773
rect 21117 9764 21129 9767
rect 19108 9736 21129 9764
rect 18449 9727 18507 9733
rect 21117 9733 21129 9736
rect 21163 9764 21175 9767
rect 21482 9764 21488 9776
rect 21163 9736 21488 9764
rect 21163 9733 21175 9736
rect 21117 9727 21175 9733
rect 21482 9724 21488 9736
rect 21540 9724 21546 9776
rect 23690 9724 23696 9776
rect 23748 9764 23754 9776
rect 23846 9764 23874 9872
rect 23969 9869 23981 9872
rect 24015 9869 24027 9903
rect 23969 9863 24027 9869
rect 24153 9903 24211 9909
rect 24153 9869 24165 9903
rect 24199 9900 24211 9903
rect 24610 9900 24616 9912
rect 24199 9872 24616 9900
rect 24199 9869 24211 9872
rect 24153 9863 24211 9869
rect 24610 9860 24616 9872
rect 24668 9860 24674 9912
rect 25714 9900 25720 9912
rect 25675 9872 25720 9900
rect 25714 9860 25720 9872
rect 25772 9860 25778 9912
rect 26174 9900 26180 9912
rect 26135 9872 26180 9900
rect 26174 9860 26180 9872
rect 26232 9860 26238 9912
rect 28017 9903 28075 9909
rect 28017 9869 28029 9903
rect 28063 9900 28075 9903
rect 29210 9900 29216 9912
rect 28063 9872 29216 9900
rect 28063 9869 28075 9872
rect 28017 9863 28075 9869
rect 29210 9860 29216 9872
rect 29268 9860 29274 9912
rect 29305 9903 29363 9909
rect 29305 9869 29317 9903
rect 29351 9869 29363 9903
rect 29305 9863 29363 9869
rect 25257 9835 25315 9841
rect 25257 9801 25269 9835
rect 25303 9832 25315 9835
rect 25303 9804 25852 9832
rect 25303 9801 25315 9804
rect 25257 9795 25315 9801
rect 25346 9764 25352 9776
rect 23748 9736 23874 9764
rect 25307 9736 25352 9764
rect 23748 9724 23754 9736
rect 25346 9724 25352 9736
rect 25404 9724 25410 9776
rect 25824 9773 25852 9804
rect 25809 9767 25867 9773
rect 25809 9733 25821 9767
rect 25855 9764 25867 9767
rect 27094 9764 27100 9776
rect 25855 9736 27100 9764
rect 25855 9733 25867 9736
rect 25809 9727 25867 9733
rect 27094 9724 27100 9736
rect 27152 9724 27158 9776
rect 27278 9724 27284 9776
rect 27336 9764 27342 9776
rect 28201 9767 28259 9773
rect 28201 9764 28213 9767
rect 27336 9736 28213 9764
rect 27336 9724 27342 9736
rect 28201 9733 28213 9736
rect 28247 9764 28259 9767
rect 29320 9764 29348 9863
rect 29578 9860 29584 9912
rect 29636 9900 29642 9912
rect 29762 9900 29768 9912
rect 29636 9872 29681 9900
rect 29723 9872 29768 9900
rect 29636 9860 29642 9872
rect 29762 9860 29768 9872
rect 29820 9860 29826 9912
rect 28247 9736 29348 9764
rect 28247 9733 28259 9736
rect 28201 9727 28259 9733
rect 400 9674 31680 9696
rect 400 9622 18870 9674
rect 18922 9622 18934 9674
rect 18986 9622 18998 9674
rect 19050 9622 19062 9674
rect 19114 9622 19126 9674
rect 19178 9622 31680 9674
rect 400 9600 31680 9622
rect 2070 9560 2076 9572
rect 2031 9532 2076 9560
rect 2070 9520 2076 9532
rect 2128 9520 2134 9572
rect 8786 9520 8792 9572
rect 8844 9560 8850 9572
rect 8973 9563 9031 9569
rect 8973 9560 8985 9563
rect 8844 9532 8985 9560
rect 8844 9520 8850 9532
rect 8973 9529 8985 9532
rect 9019 9529 9031 9563
rect 8973 9523 9031 9529
rect 11825 9563 11883 9569
rect 11825 9529 11837 9563
rect 11871 9560 11883 9563
rect 12282 9560 12288 9572
rect 11871 9532 12288 9560
rect 11871 9529 11883 9532
rect 11825 9523 11883 9529
rect 12282 9520 12288 9532
rect 12340 9520 12346 9572
rect 14674 9560 14680 9572
rect 14635 9532 14680 9560
rect 14674 9520 14680 9532
rect 14732 9520 14738 9572
rect 18630 9560 18636 9572
rect 18591 9532 18636 9560
rect 18630 9520 18636 9532
rect 18688 9520 18694 9572
rect 18722 9520 18728 9572
rect 18780 9560 18786 9572
rect 18817 9563 18875 9569
rect 18817 9560 18829 9563
rect 18780 9532 18829 9560
rect 18780 9520 18786 9532
rect 18817 9529 18829 9532
rect 18863 9529 18875 9563
rect 18817 9523 18875 9529
rect 19093 9563 19151 9569
rect 19093 9529 19105 9563
rect 19139 9560 19151 9563
rect 19274 9560 19280 9572
rect 19139 9532 19280 9560
rect 19139 9529 19151 9532
rect 19093 9523 19151 9529
rect 19274 9520 19280 9532
rect 19332 9520 19338 9572
rect 24610 9560 24616 9572
rect 24571 9532 24616 9560
rect 24610 9520 24616 9532
rect 24668 9520 24674 9572
rect 24702 9520 24708 9572
rect 24760 9560 24766 9572
rect 24797 9563 24855 9569
rect 24797 9560 24809 9563
rect 24760 9532 24809 9560
rect 24760 9520 24766 9532
rect 24797 9529 24809 9532
rect 24843 9560 24855 9563
rect 25530 9560 25536 9572
rect 24843 9532 25536 9560
rect 24843 9529 24855 9532
rect 24797 9523 24855 9529
rect 25530 9520 25536 9532
rect 25588 9520 25594 9572
rect 25898 9560 25904 9572
rect 25859 9532 25904 9560
rect 25898 9520 25904 9532
rect 25956 9520 25962 9572
rect 2346 9452 2352 9504
rect 2404 9492 2410 9504
rect 3174 9492 3180 9504
rect 2404 9464 3180 9492
rect 2404 9452 2410 9464
rect 3174 9452 3180 9464
rect 3232 9492 3238 9504
rect 3361 9495 3419 9501
rect 3361 9492 3373 9495
rect 3232 9464 3373 9492
rect 3232 9452 3238 9464
rect 3361 9461 3373 9464
rect 3407 9461 3419 9495
rect 3361 9455 3419 9461
rect 4094 9452 4100 9504
rect 4152 9492 4158 9504
rect 5474 9492 5480 9504
rect 4152 9464 5480 9492
rect 4152 9452 4158 9464
rect 5474 9452 5480 9464
rect 5532 9452 5538 9504
rect 9338 9492 9344 9504
rect 9299 9464 9344 9492
rect 9338 9452 9344 9464
rect 9396 9452 9402 9504
rect 14766 9452 14772 9504
rect 14824 9492 14830 9504
rect 15873 9495 15931 9501
rect 15873 9492 15885 9495
rect 14824 9464 15885 9492
rect 14824 9452 14830 9464
rect 15873 9461 15885 9464
rect 15919 9461 15931 9495
rect 15873 9455 15931 9461
rect 17342 9452 17348 9504
rect 17400 9492 17406 9504
rect 17400 9464 18400 9492
rect 17400 9452 17406 9464
rect 1150 9424 1156 9436
rect 1111 9396 1156 9424
rect 1150 9384 1156 9396
rect 1208 9424 1214 9436
rect 1705 9427 1763 9433
rect 1705 9424 1717 9427
rect 1208 9396 1717 9424
rect 1208 9384 1214 9396
rect 1705 9393 1717 9396
rect 1751 9424 1763 9427
rect 2438 9424 2444 9436
rect 1751 9396 2444 9424
rect 1751 9393 1763 9396
rect 1705 9387 1763 9393
rect 2438 9384 2444 9396
rect 2496 9384 2502 9436
rect 3821 9427 3879 9433
rect 3821 9393 3833 9427
rect 3867 9424 3879 9427
rect 3910 9424 3916 9436
rect 3867 9396 3916 9424
rect 3867 9393 3879 9396
rect 3821 9387 3879 9393
rect 3910 9384 3916 9396
rect 3968 9384 3974 9436
rect 4002 9384 4008 9436
rect 4060 9424 4066 9436
rect 4186 9424 4192 9436
rect 4060 9396 4105 9424
rect 4147 9396 4192 9424
rect 4060 9384 4066 9396
rect 4186 9384 4192 9396
rect 4244 9384 4250 9436
rect 5566 9384 5572 9436
rect 5624 9424 5630 9436
rect 5661 9427 5719 9433
rect 5661 9424 5673 9427
rect 5624 9396 5673 9424
rect 5624 9384 5630 9396
rect 5661 9393 5673 9396
rect 5707 9393 5719 9427
rect 9982 9424 9988 9436
rect 9943 9396 9988 9424
rect 5661 9387 5719 9393
rect 9982 9384 9988 9396
rect 10040 9384 10046 9436
rect 10350 9424 10356 9436
rect 10311 9396 10356 9424
rect 10350 9384 10356 9396
rect 10408 9384 10414 9436
rect 15962 9384 15968 9436
rect 16020 9424 16026 9436
rect 16057 9427 16115 9433
rect 16057 9424 16069 9427
rect 16020 9396 16069 9424
rect 16020 9384 16026 9396
rect 16057 9393 16069 9396
rect 16103 9393 16115 9427
rect 17986 9424 17992 9436
rect 17947 9396 17992 9424
rect 16057 9387 16115 9393
rect 17986 9384 17992 9396
rect 18044 9384 18050 9436
rect 18372 9433 18400 9464
rect 23230 9452 23236 9504
rect 23288 9452 23294 9504
rect 26085 9495 26143 9501
rect 26085 9461 26097 9495
rect 26131 9492 26143 9495
rect 26358 9492 26364 9504
rect 26131 9464 26364 9492
rect 26131 9461 26143 9464
rect 26085 9455 26143 9461
rect 26358 9452 26364 9464
rect 26416 9492 26422 9504
rect 27554 9492 27560 9504
rect 26416 9464 27560 9492
rect 26416 9452 26422 9464
rect 27554 9452 27560 9464
rect 27612 9452 27618 9504
rect 27646 9452 27652 9504
rect 27704 9492 27710 9504
rect 28382 9492 28388 9504
rect 27704 9464 28388 9492
rect 27704 9452 27710 9464
rect 28382 9452 28388 9464
rect 28440 9452 28446 9504
rect 28566 9452 28572 9504
rect 28624 9492 28630 9504
rect 28624 9464 29072 9492
rect 28624 9452 28630 9464
rect 18357 9427 18415 9433
rect 18357 9393 18369 9427
rect 18403 9393 18415 9427
rect 18357 9387 18415 9393
rect 19277 9427 19335 9433
rect 19277 9393 19289 9427
rect 19323 9424 19335 9427
rect 19366 9424 19372 9436
rect 19323 9396 19372 9424
rect 19323 9393 19335 9396
rect 19277 9387 19335 9393
rect 19366 9384 19372 9396
rect 19424 9384 19430 9436
rect 22494 9424 22500 9436
rect 22455 9396 22500 9424
rect 22494 9384 22500 9396
rect 22552 9384 22558 9436
rect 22862 9424 22868 9436
rect 22823 9396 22868 9424
rect 22862 9384 22868 9396
rect 22920 9384 22926 9436
rect 26634 9424 26640 9436
rect 26595 9396 26640 9424
rect 26634 9384 26640 9396
rect 26692 9384 26698 9436
rect 26729 9427 26787 9433
rect 26729 9393 26741 9427
rect 26775 9393 26787 9427
rect 27002 9424 27008 9436
rect 26963 9396 27008 9424
rect 26729 9387 26787 9393
rect 969 9359 1027 9365
rect 969 9325 981 9359
rect 1015 9356 1027 9359
rect 1426 9356 1432 9368
rect 1015 9328 1432 9356
rect 1015 9325 1027 9328
rect 969 9319 1027 9325
rect 1426 9316 1432 9328
rect 1484 9316 1490 9368
rect 6026 9356 6032 9368
rect 5987 9328 6032 9356
rect 6026 9316 6032 9328
rect 6084 9316 6090 9368
rect 9430 9316 9436 9368
rect 9488 9356 9494 9368
rect 9614 9356 9620 9368
rect 9488 9328 9620 9356
rect 9488 9316 9494 9328
rect 9614 9316 9620 9328
rect 9672 9356 9678 9368
rect 9801 9359 9859 9365
rect 9801 9356 9813 9359
rect 9672 9328 9813 9356
rect 9672 9316 9678 9328
rect 9801 9325 9813 9328
rect 9847 9325 9859 9359
rect 9801 9319 9859 9325
rect 10261 9359 10319 9365
rect 10261 9325 10273 9359
rect 10307 9356 10319 9359
rect 10810 9356 10816 9368
rect 10307 9328 10816 9356
rect 10307 9325 10319 9328
rect 10261 9319 10319 9325
rect 9706 9248 9712 9300
rect 9764 9288 9770 9300
rect 10276 9288 10304 9319
rect 10810 9316 10816 9328
rect 10868 9316 10874 9368
rect 18078 9356 18084 9368
rect 18039 9328 18084 9356
rect 18078 9316 18084 9328
rect 18136 9316 18142 9368
rect 18446 9356 18452 9368
rect 18407 9328 18452 9356
rect 18446 9316 18452 9328
rect 18504 9316 18510 9368
rect 22770 9316 22776 9368
rect 22828 9356 22834 9368
rect 24610 9356 24616 9368
rect 22828 9328 24616 9356
rect 22828 9316 22834 9328
rect 24610 9316 24616 9328
rect 24668 9316 24674 9368
rect 25990 9316 25996 9368
rect 26048 9356 26054 9368
rect 26744 9356 26772 9387
rect 27002 9384 27008 9396
rect 27060 9384 27066 9436
rect 27462 9424 27468 9436
rect 27296 9396 27468 9424
rect 27186 9356 27192 9368
rect 26048 9328 26772 9356
rect 27147 9328 27192 9356
rect 26048 9316 26054 9328
rect 27186 9316 27192 9328
rect 27244 9316 27250 9368
rect 9764 9260 10304 9288
rect 9764 9248 9770 9260
rect 25714 9248 25720 9300
rect 25772 9288 25778 9300
rect 27296 9288 27324 9396
rect 27462 9384 27468 9396
rect 27520 9384 27526 9436
rect 28842 9424 28848 9436
rect 28803 9396 28848 9424
rect 28842 9384 28848 9396
rect 28900 9384 28906 9436
rect 29044 9433 29072 9464
rect 29029 9427 29087 9433
rect 29029 9393 29041 9427
rect 29075 9393 29087 9427
rect 29029 9387 29087 9393
rect 29118 9384 29124 9436
rect 29176 9424 29182 9436
rect 29213 9427 29271 9433
rect 29213 9424 29225 9427
rect 29176 9396 29225 9424
rect 29176 9384 29182 9396
rect 29213 9393 29225 9396
rect 29259 9393 29271 9427
rect 29213 9387 29271 9393
rect 28658 9316 28664 9368
rect 28716 9356 28722 9368
rect 29489 9359 29547 9365
rect 29489 9356 29501 9359
rect 28716 9328 29501 9356
rect 28716 9316 28722 9328
rect 29489 9325 29501 9328
rect 29535 9325 29547 9359
rect 29489 9319 29547 9325
rect 29765 9359 29823 9365
rect 29765 9325 29777 9359
rect 29811 9325 29823 9359
rect 29765 9319 29823 9325
rect 25772 9260 27324 9288
rect 25772 9248 25778 9260
rect 28474 9248 28480 9300
rect 28532 9288 28538 9300
rect 29780 9288 29808 9319
rect 30038 9288 30044 9300
rect 28532 9260 30044 9288
rect 28532 9248 28538 9260
rect 30038 9248 30044 9260
rect 30096 9248 30102 9300
rect 785 9223 843 9229
rect 785 9189 797 9223
rect 831 9220 843 9223
rect 1610 9220 1616 9232
rect 831 9192 1616 9220
rect 831 9189 843 9192
rect 785 9183 843 9189
rect 1610 9180 1616 9192
rect 1668 9180 1674 9232
rect 6213 9223 6271 9229
rect 6213 9189 6225 9223
rect 6259 9220 6271 9223
rect 6486 9220 6492 9232
rect 6259 9192 6492 9220
rect 6259 9189 6271 9192
rect 6213 9183 6271 9189
rect 6486 9180 6492 9192
rect 6544 9180 6550 9232
rect 12006 9220 12012 9232
rect 11967 9192 12012 9220
rect 12006 9180 12012 9192
rect 12064 9180 12070 9232
rect 16146 9220 16152 9232
rect 16107 9192 16152 9220
rect 16146 9180 16152 9192
rect 16204 9180 16210 9232
rect 17437 9223 17495 9229
rect 17437 9189 17449 9223
rect 17483 9220 17495 9223
rect 17526 9220 17532 9232
rect 17483 9192 17532 9220
rect 17483 9189 17495 9192
rect 17437 9183 17495 9189
rect 17526 9180 17532 9192
rect 17584 9180 17590 9232
rect 400 9130 31680 9152
rect 400 9078 3510 9130
rect 3562 9078 3574 9130
rect 3626 9078 3638 9130
rect 3690 9078 3702 9130
rect 3754 9078 3766 9130
rect 3818 9078 31680 9130
rect 400 9056 31680 9078
rect 2070 9016 2076 9028
rect 708 8988 2076 9016
rect 708 8892 736 8988
rect 2070 8976 2076 8988
rect 2128 8976 2134 9028
rect 3174 9016 3180 9028
rect 3135 8988 3180 9016
rect 3174 8976 3180 8988
rect 3232 8976 3238 9028
rect 4462 9016 4468 9028
rect 4423 8988 4468 9016
rect 4462 8976 4468 8988
rect 4520 8976 4526 9028
rect 5474 9016 5480 9028
rect 5435 8988 5480 9016
rect 5474 8976 5480 8988
rect 5532 8976 5538 9028
rect 9338 8976 9344 9028
rect 9396 9016 9402 9028
rect 9525 9019 9583 9025
rect 9525 9016 9537 9019
rect 9396 8988 9537 9016
rect 9396 8976 9402 8988
rect 9525 8985 9537 8988
rect 9571 8985 9583 9019
rect 9525 8979 9583 8985
rect 14582 8976 14588 9028
rect 14640 9016 14646 9028
rect 15505 9019 15563 9025
rect 15505 9016 15517 9019
rect 14640 8988 15517 9016
rect 14640 8976 14646 8988
rect 15505 8985 15517 8988
rect 15551 9016 15563 9019
rect 15686 9016 15692 9028
rect 15551 8988 15692 9016
rect 15551 8985 15563 8988
rect 15505 8979 15563 8985
rect 15686 8976 15692 8988
rect 15744 8976 15750 9028
rect 15962 9016 15968 9028
rect 15923 8988 15968 9016
rect 15962 8976 15968 8988
rect 16020 8976 16026 9028
rect 16146 8976 16152 9028
rect 16204 9016 16210 9028
rect 16241 9019 16299 9025
rect 16241 9016 16253 9019
rect 16204 8988 16253 9016
rect 16204 8976 16210 8988
rect 16241 8985 16253 8988
rect 16287 8985 16299 9019
rect 16241 8979 16299 8985
rect 16977 9019 17035 9025
rect 16977 8985 16989 9019
rect 17023 9016 17035 9019
rect 18446 9016 18452 9028
rect 17023 8988 18452 9016
rect 17023 8985 17035 8988
rect 16977 8979 17035 8985
rect 18446 8976 18452 8988
rect 18504 8976 18510 9028
rect 19093 9019 19151 9025
rect 19093 8985 19105 9019
rect 19139 9016 19151 9019
rect 19366 9016 19372 9028
rect 19139 8988 19372 9016
rect 19139 8985 19151 8988
rect 19093 8979 19151 8985
rect 19366 8976 19372 8988
rect 19424 8976 19430 9028
rect 22770 9016 22776 9028
rect 22731 8988 22776 9016
rect 22770 8976 22776 8988
rect 22828 8976 22834 9028
rect 22862 8976 22868 9028
rect 22920 9016 22926 9028
rect 22957 9019 23015 9025
rect 22957 9016 22969 9019
rect 22920 8988 22969 9016
rect 22920 8976 22926 8988
rect 22957 8985 22969 8988
rect 23003 8985 23015 9019
rect 24702 9016 24708 9028
rect 24663 8988 24708 9016
rect 22957 8979 23015 8985
rect 24702 8976 24708 8988
rect 24760 8976 24766 9028
rect 25530 8976 25536 9028
rect 25588 9016 25594 9028
rect 26361 9019 26419 9025
rect 26361 9016 26373 9019
rect 25588 8988 26373 9016
rect 25588 8976 25594 8988
rect 26361 8985 26373 8988
rect 26407 9016 26419 9019
rect 27186 9016 27192 9028
rect 26407 8988 27192 9016
rect 26407 8985 26419 8988
rect 26361 8979 26419 8985
rect 27186 8976 27192 8988
rect 27244 8976 27250 9028
rect 27462 8976 27468 9028
rect 27520 9016 27526 9028
rect 28293 9019 28351 9025
rect 28293 9016 28305 9019
rect 27520 8988 28305 9016
rect 27520 8976 27526 8988
rect 28293 8985 28305 8988
rect 28339 9016 28351 9019
rect 28474 9016 28480 9028
rect 28339 8988 28480 9016
rect 28339 8985 28351 8988
rect 28293 8979 28351 8985
rect 28474 8976 28480 8988
rect 28532 8976 28538 9028
rect 28661 9019 28719 9025
rect 28661 8985 28673 9019
rect 28707 9016 28719 9019
rect 29118 9016 29124 9028
rect 28707 8988 29124 9016
rect 28707 8985 28719 8988
rect 28661 8979 28719 8985
rect 29118 8976 29124 8988
rect 29176 8976 29182 9028
rect 29210 8976 29216 9028
rect 29268 9016 29274 9028
rect 29489 9019 29547 9025
rect 29489 9016 29501 9019
rect 29268 8988 29501 9016
rect 29268 8976 29274 8988
rect 29489 8985 29501 8988
rect 29535 9016 29547 9019
rect 30041 9019 30099 9025
rect 30041 9016 30053 9019
rect 29535 8988 30053 9016
rect 29535 8985 29547 8988
rect 29489 8979 29547 8985
rect 30041 8985 30053 8988
rect 30087 8985 30099 9019
rect 30041 8979 30099 8985
rect 5201 8951 5259 8957
rect 5201 8917 5213 8951
rect 5247 8948 5259 8951
rect 6026 8948 6032 8960
rect 5247 8920 6032 8948
rect 5247 8917 5259 8920
rect 5201 8911 5259 8917
rect 6026 8908 6032 8920
rect 6084 8908 6090 8960
rect 7866 8908 7872 8960
rect 7924 8948 7930 8960
rect 8694 8948 8700 8960
rect 7924 8920 8700 8948
rect 7924 8908 7930 8920
rect 8694 8908 8700 8920
rect 8752 8948 8758 8960
rect 9893 8951 9951 8957
rect 9893 8948 9905 8951
rect 8752 8920 9905 8948
rect 8752 8908 8758 8920
rect 9893 8917 9905 8920
rect 9939 8948 9951 8951
rect 10350 8948 10356 8960
rect 9939 8920 10356 8948
rect 9939 8917 9951 8920
rect 9893 8911 9951 8917
rect 10350 8908 10356 8920
rect 10408 8948 10414 8960
rect 11181 8951 11239 8957
rect 11181 8948 11193 8951
rect 10408 8920 11193 8948
rect 10408 8908 10414 8920
rect 11181 8917 11193 8920
rect 11227 8948 11239 8951
rect 12742 8948 12748 8960
rect 11227 8920 12748 8948
rect 11227 8917 11239 8920
rect 11181 8911 11239 8917
rect 12742 8908 12748 8920
rect 12800 8908 12806 8960
rect 18262 8908 18268 8960
rect 18320 8948 18326 8960
rect 18817 8951 18875 8957
rect 18817 8948 18829 8951
rect 18320 8920 18829 8948
rect 18320 8908 18326 8920
rect 18817 8917 18829 8920
rect 18863 8917 18875 8951
rect 18817 8911 18875 8917
rect 690 8880 696 8892
rect 603 8852 696 8880
rect 690 8840 696 8852
rect 748 8840 754 8892
rect 1610 8840 1616 8892
rect 1668 8880 1674 8892
rect 2717 8883 2775 8889
rect 2717 8880 2729 8883
rect 1668 8852 2729 8880
rect 1668 8840 1674 8852
rect 2717 8849 2729 8852
rect 2763 8880 2775 8883
rect 3361 8883 3419 8889
rect 3361 8880 3373 8883
rect 2763 8852 3373 8880
rect 2763 8849 2775 8852
rect 2717 8843 2775 8849
rect 3361 8849 3373 8852
rect 3407 8880 3419 8883
rect 3545 8883 3603 8889
rect 3545 8880 3557 8883
rect 3407 8852 3557 8880
rect 3407 8849 3419 8852
rect 3361 8843 3419 8849
rect 3545 8849 3557 8852
rect 3591 8880 3603 8883
rect 4186 8880 4192 8892
rect 3591 8852 4192 8880
rect 3591 8849 3603 8852
rect 3545 8843 3603 8849
rect 4186 8840 4192 8852
rect 4244 8840 4250 8892
rect 4738 8840 4744 8892
rect 4796 8880 4802 8892
rect 5661 8883 5719 8889
rect 5661 8880 5673 8883
rect 4796 8852 5673 8880
rect 4796 8840 4802 8852
rect 5661 8849 5673 8852
rect 5707 8880 5719 8883
rect 6486 8880 6492 8892
rect 5707 8852 6348 8880
rect 6447 8852 6492 8880
rect 5707 8849 5719 8852
rect 5661 8843 5719 8849
rect 3634 8812 3640 8824
rect 3547 8784 3640 8812
rect 3634 8772 3640 8784
rect 3692 8812 3698 8824
rect 4462 8812 4468 8824
rect 3692 8784 4468 8812
rect 3692 8772 3698 8784
rect 4462 8772 4468 8784
rect 4520 8772 4526 8824
rect 6118 8812 6124 8824
rect 6079 8784 6124 8812
rect 6118 8772 6124 8784
rect 6176 8772 6182 8824
rect 6320 8812 6348 8852
rect 6486 8840 6492 8852
rect 6544 8840 6550 8892
rect 7406 8880 7412 8892
rect 6596 8852 7412 8880
rect 6596 8812 6624 8852
rect 7406 8840 7412 8852
rect 7464 8880 7470 8892
rect 7961 8883 8019 8889
rect 7961 8880 7973 8883
rect 7464 8852 7973 8880
rect 7464 8840 7470 8852
rect 7961 8849 7973 8852
rect 8007 8849 8019 8883
rect 7961 8843 8019 8849
rect 8418 8840 8424 8892
rect 8476 8880 8482 8892
rect 9341 8883 9399 8889
rect 9341 8880 9353 8883
rect 8476 8852 9353 8880
rect 8476 8840 8482 8852
rect 9341 8849 9353 8852
rect 9387 8880 9399 8883
rect 9706 8880 9712 8892
rect 9387 8852 9712 8880
rect 9387 8849 9399 8852
rect 9341 8843 9399 8849
rect 9706 8840 9712 8852
rect 9764 8840 9770 8892
rect 9982 8840 9988 8892
rect 10040 8880 10046 8892
rect 10169 8883 10227 8889
rect 10169 8880 10181 8883
rect 10040 8852 10181 8880
rect 10040 8840 10046 8852
rect 10169 8849 10181 8852
rect 10215 8880 10227 8883
rect 12006 8880 12012 8892
rect 10215 8852 12012 8880
rect 10215 8849 10227 8852
rect 10169 8843 10227 8849
rect 12006 8840 12012 8852
rect 12064 8880 12070 8892
rect 12650 8880 12656 8892
rect 12064 8852 12420 8880
rect 12611 8852 12656 8880
rect 12064 8840 12070 8852
rect 6320 8784 6624 8812
rect 12193 8815 12251 8821
rect 12193 8781 12205 8815
rect 12239 8812 12251 8815
rect 12282 8812 12288 8824
rect 12239 8784 12288 8812
rect 12239 8781 12251 8784
rect 12193 8775 12251 8781
rect 12282 8772 12288 8784
rect 12340 8772 12346 8824
rect 12392 8821 12420 8852
rect 12650 8840 12656 8852
rect 12708 8840 12714 8892
rect 16793 8883 16851 8889
rect 16793 8849 16805 8883
rect 16839 8880 16851 8883
rect 17986 8880 17992 8892
rect 16839 8852 17992 8880
rect 16839 8849 16851 8852
rect 16793 8843 16851 8849
rect 17986 8840 17992 8852
rect 18044 8840 18050 8892
rect 18832 8880 18860 8911
rect 22494 8908 22500 8960
rect 22552 8948 22558 8960
rect 23141 8951 23199 8957
rect 23141 8948 23153 8951
rect 22552 8920 23153 8948
rect 22552 8908 22558 8920
rect 23141 8917 23153 8920
rect 23187 8917 23199 8951
rect 23141 8911 23199 8917
rect 23785 8951 23843 8957
rect 23785 8917 23797 8951
rect 23831 8948 23843 8951
rect 24337 8951 24395 8957
rect 23831 8920 24288 8948
rect 23831 8917 23843 8920
rect 23785 8911 23843 8917
rect 22589 8883 22647 8889
rect 18832 8852 20056 8880
rect 12377 8815 12435 8821
rect 12377 8781 12389 8815
rect 12423 8781 12435 8815
rect 12742 8812 12748 8824
rect 12703 8784 12748 8812
rect 12377 8775 12435 8781
rect 12742 8772 12748 8784
rect 12800 8772 12806 8824
rect 14186 8784 14720 8812
rect 966 8744 972 8756
rect 927 8716 972 8744
rect 966 8704 972 8716
rect 1024 8704 1030 8756
rect 1426 8704 1432 8756
rect 1484 8704 1490 8756
rect 2898 8744 2904 8756
rect 2811 8716 2904 8744
rect 2898 8704 2904 8716
rect 2956 8744 2962 8756
rect 4097 8747 4155 8753
rect 4097 8744 4109 8747
rect 2956 8716 4109 8744
rect 2956 8704 2962 8716
rect 4097 8713 4109 8716
rect 4143 8713 4155 8747
rect 4097 8707 4155 8713
rect 7314 8704 7320 8756
rect 7372 8704 7378 8756
rect 11178 8704 11184 8756
rect 11236 8744 11242 8756
rect 11365 8747 11423 8753
rect 11365 8744 11377 8747
rect 11236 8716 11377 8744
rect 11236 8704 11242 8716
rect 11365 8713 11377 8716
rect 11411 8744 11423 8747
rect 11733 8747 11791 8753
rect 11733 8744 11745 8747
rect 11411 8716 11745 8744
rect 11411 8713 11423 8716
rect 11365 8707 11423 8713
rect 11733 8713 11745 8716
rect 11779 8713 11791 8747
rect 11733 8707 11791 8713
rect 12650 8704 12656 8756
rect 12708 8744 12714 8756
rect 14186 8744 14214 8784
rect 14582 8744 14588 8756
rect 12708 8716 14214 8744
rect 14543 8716 14588 8744
rect 12708 8704 12714 8716
rect 14582 8704 14588 8716
rect 14640 8704 14646 8756
rect 14692 8744 14720 8784
rect 14766 8772 14772 8824
rect 14824 8812 14830 8824
rect 15229 8815 15287 8821
rect 15229 8812 15241 8815
rect 14824 8784 15241 8812
rect 14824 8772 14830 8784
rect 15229 8781 15241 8784
rect 15275 8812 15287 8815
rect 16057 8815 16115 8821
rect 16057 8812 16069 8815
rect 15275 8784 16069 8812
rect 15275 8781 15287 8784
rect 15229 8775 15287 8781
rect 16057 8781 16069 8784
rect 16103 8781 16115 8815
rect 16057 8775 16115 8781
rect 17434 8772 17440 8824
rect 17492 8812 17498 8824
rect 17529 8815 17587 8821
rect 17529 8812 17541 8815
rect 17492 8784 17541 8812
rect 17492 8772 17498 8784
rect 17529 8781 17541 8784
rect 17575 8812 17587 8815
rect 18265 8815 18323 8821
rect 18265 8812 18277 8815
rect 17575 8784 18277 8812
rect 17575 8781 17587 8784
rect 17529 8775 17587 8781
rect 18265 8781 18277 8784
rect 18311 8781 18323 8815
rect 18265 8775 18323 8781
rect 18541 8815 18599 8821
rect 18541 8781 18553 8815
rect 18587 8812 18599 8815
rect 18722 8812 18728 8824
rect 18587 8784 18728 8812
rect 18587 8781 18599 8784
rect 18541 8775 18599 8781
rect 18722 8772 18728 8784
rect 18780 8812 18786 8824
rect 20028 8821 20056 8852
rect 22589 8849 22601 8883
rect 22635 8880 22647 8883
rect 23322 8880 23328 8892
rect 22635 8852 23328 8880
rect 22635 8849 22647 8852
rect 22589 8843 22647 8849
rect 23322 8840 23328 8852
rect 23380 8840 23386 8892
rect 24260 8880 24288 8920
rect 24337 8917 24349 8951
rect 24383 8948 24395 8951
rect 24610 8948 24616 8960
rect 24383 8920 24616 8948
rect 24383 8917 24395 8920
rect 24337 8911 24395 8917
rect 24610 8908 24616 8920
rect 24668 8948 24674 8960
rect 25622 8948 25628 8960
rect 24668 8920 25628 8948
rect 24668 8908 24674 8920
rect 25622 8908 25628 8920
rect 25680 8908 25686 8960
rect 26177 8951 26235 8957
rect 26177 8917 26189 8951
rect 26223 8948 26235 8951
rect 27002 8948 27008 8960
rect 26223 8920 27008 8948
rect 26223 8917 26235 8920
rect 26177 8911 26235 8917
rect 27002 8908 27008 8920
rect 27060 8908 27066 8960
rect 29026 8908 29032 8960
rect 29084 8948 29090 8960
rect 29857 8951 29915 8957
rect 29857 8948 29869 8951
rect 29084 8920 29869 8948
rect 29084 8908 29090 8920
rect 29857 8917 29869 8920
rect 29903 8917 29915 8951
rect 29857 8911 29915 8917
rect 25165 8883 25223 8889
rect 25165 8880 25177 8883
rect 24260 8852 25177 8880
rect 25165 8849 25177 8852
rect 25211 8880 25223 8883
rect 25898 8880 25904 8892
rect 25211 8852 25904 8880
rect 25211 8849 25223 8852
rect 25165 8843 25223 8849
rect 25898 8840 25904 8852
rect 25956 8840 25962 8892
rect 26634 8840 26640 8892
rect 26692 8880 26698 8892
rect 26692 8852 28060 8880
rect 26692 8840 26698 8852
rect 19645 8815 19703 8821
rect 19645 8812 19657 8815
rect 18780 8784 19657 8812
rect 18780 8772 18786 8784
rect 19645 8781 19657 8784
rect 19691 8781 19703 8815
rect 19645 8775 19703 8781
rect 19737 8815 19795 8821
rect 19737 8781 19749 8815
rect 19783 8781 19795 8815
rect 19737 8775 19795 8781
rect 20013 8815 20071 8821
rect 20013 8781 20025 8815
rect 20059 8781 20071 8815
rect 20013 8775 20071 8781
rect 20197 8815 20255 8821
rect 20197 8781 20209 8815
rect 20243 8812 20255 8815
rect 21206 8812 21212 8824
rect 20243 8784 21212 8812
rect 20243 8781 20255 8784
rect 20197 8775 20255 8781
rect 17342 8744 17348 8756
rect 14692 8716 17348 8744
rect 17342 8704 17348 8716
rect 17400 8704 17406 8756
rect 17802 8744 17808 8756
rect 17763 8716 17808 8744
rect 17802 8704 17808 8716
rect 17860 8704 17866 8756
rect 18078 8704 18084 8756
rect 18136 8744 18142 8756
rect 18173 8747 18231 8753
rect 18173 8744 18185 8747
rect 18136 8716 18185 8744
rect 18136 8704 18142 8716
rect 18173 8713 18185 8716
rect 18219 8744 18231 8747
rect 18633 8747 18691 8753
rect 18633 8744 18645 8747
rect 18219 8716 18645 8744
rect 18219 8713 18231 8716
rect 18173 8707 18231 8713
rect 18633 8713 18645 8716
rect 18679 8744 18691 8747
rect 19752 8744 19780 8775
rect 21206 8772 21212 8784
rect 21264 8772 21270 8824
rect 24153 8815 24211 8821
rect 24153 8781 24165 8815
rect 24199 8812 24211 8815
rect 25073 8815 25131 8821
rect 25073 8812 25085 8815
rect 24199 8784 25085 8812
rect 24199 8781 24211 8784
rect 24153 8775 24211 8781
rect 25073 8781 25085 8784
rect 25119 8812 25131 8815
rect 25346 8812 25352 8824
rect 25119 8784 25352 8812
rect 25119 8781 25131 8784
rect 25073 8775 25131 8781
rect 25346 8772 25352 8784
rect 25404 8772 25410 8824
rect 25441 8815 25499 8821
rect 25441 8781 25453 8815
rect 25487 8781 25499 8815
rect 25622 8812 25628 8824
rect 25583 8784 25628 8812
rect 25441 8775 25499 8781
rect 21758 8744 21764 8756
rect 18679 8716 21764 8744
rect 18679 8713 18691 8716
rect 18633 8707 18691 8713
rect 21758 8704 21764 8716
rect 21816 8704 21822 8756
rect 23969 8747 24027 8753
rect 23969 8713 23981 8747
rect 24015 8744 24027 8747
rect 25162 8744 25168 8756
rect 24015 8716 25168 8744
rect 24015 8713 24027 8716
rect 23969 8707 24027 8713
rect 25162 8704 25168 8716
rect 25220 8744 25226 8756
rect 25456 8744 25484 8775
rect 25622 8772 25628 8784
rect 25680 8772 25686 8824
rect 27094 8812 27100 8824
rect 27055 8784 27100 8812
rect 27094 8772 27100 8784
rect 27152 8772 27158 8824
rect 27189 8815 27247 8821
rect 27189 8781 27201 8815
rect 27235 8812 27247 8815
rect 27278 8812 27284 8824
rect 27235 8784 27284 8812
rect 27235 8781 27247 8784
rect 27189 8775 27247 8781
rect 27278 8772 27284 8784
rect 27336 8772 27342 8824
rect 27462 8812 27468 8824
rect 27423 8784 27468 8812
rect 27462 8772 27468 8784
rect 27520 8772 27526 8824
rect 27646 8812 27652 8824
rect 27607 8784 27652 8812
rect 27646 8772 27652 8784
rect 27704 8772 27710 8824
rect 28032 8821 28060 8852
rect 28017 8815 28075 8821
rect 28017 8781 28029 8815
rect 28063 8812 28075 8815
rect 28842 8812 28848 8824
rect 28063 8784 28848 8812
rect 28063 8781 28075 8784
rect 28017 8775 28075 8781
rect 28842 8772 28848 8784
rect 28900 8812 28906 8824
rect 29305 8815 29363 8821
rect 29305 8812 29317 8815
rect 28900 8784 29317 8812
rect 28900 8772 28906 8784
rect 29305 8781 29317 8784
rect 29351 8812 29363 8815
rect 29394 8812 29400 8824
rect 29351 8784 29400 8812
rect 29351 8781 29363 8784
rect 29305 8775 29363 8781
rect 29394 8772 29400 8784
rect 29452 8772 29458 8824
rect 26450 8744 26456 8756
rect 25220 8716 25484 8744
rect 26411 8716 26456 8744
rect 25220 8704 25226 8716
rect 26450 8704 26456 8716
rect 26508 8704 26514 8756
rect 27480 8744 27508 8772
rect 28109 8747 28167 8753
rect 28109 8744 28121 8747
rect 27480 8716 28121 8744
rect 28109 8713 28121 8716
rect 28155 8713 28167 8747
rect 29210 8744 29216 8756
rect 29171 8716 29216 8744
rect 28109 8707 28167 8713
rect 29210 8704 29216 8716
rect 29268 8704 29274 8756
rect 3085 8679 3143 8685
rect 3085 8645 3097 8679
rect 3131 8676 3143 8679
rect 4002 8676 4008 8688
rect 3131 8648 4008 8676
rect 3131 8645 3143 8648
rect 3085 8639 3143 8645
rect 4002 8636 4008 8648
rect 4060 8636 4066 8688
rect 5385 8679 5443 8685
rect 5385 8645 5397 8679
rect 5431 8676 5443 8679
rect 5474 8676 5480 8688
rect 5431 8648 5480 8676
rect 5431 8645 5443 8648
rect 5385 8639 5443 8645
rect 5474 8636 5480 8648
rect 5532 8636 5538 8688
rect 5937 8679 5995 8685
rect 5937 8645 5949 8679
rect 5983 8676 5995 8679
rect 7332 8676 7360 8704
rect 7774 8676 7780 8688
rect 5983 8648 7780 8676
rect 5983 8645 5995 8648
rect 5937 8639 5995 8645
rect 7774 8636 7780 8648
rect 7832 8636 7838 8688
rect 9430 8636 9436 8688
rect 9488 8676 9494 8688
rect 9709 8679 9767 8685
rect 9709 8676 9721 8679
rect 9488 8648 9721 8676
rect 9488 8636 9494 8648
rect 9709 8645 9721 8648
rect 9755 8645 9767 8679
rect 11454 8676 11460 8688
rect 11415 8648 11460 8676
rect 9709 8639 9767 8645
rect 11454 8636 11460 8648
rect 11512 8636 11518 8688
rect 14493 8679 14551 8685
rect 14493 8645 14505 8679
rect 14539 8676 14551 8679
rect 14766 8676 14772 8688
rect 14539 8648 14772 8676
rect 14539 8645 14551 8648
rect 14493 8639 14551 8645
rect 14766 8636 14772 8648
rect 14824 8676 14830 8688
rect 14861 8679 14919 8685
rect 14861 8676 14873 8679
rect 14824 8648 14873 8676
rect 14824 8636 14830 8648
rect 14861 8645 14873 8648
rect 14907 8645 14919 8679
rect 14861 8639 14919 8645
rect 17161 8679 17219 8685
rect 17161 8645 17173 8679
rect 17207 8676 17219 8679
rect 17820 8676 17848 8704
rect 17207 8648 17848 8676
rect 17207 8645 17219 8648
rect 17161 8639 17219 8645
rect 24334 8636 24340 8688
rect 24392 8676 24398 8688
rect 25714 8676 25720 8688
rect 24392 8648 25720 8676
rect 24392 8636 24398 8648
rect 25714 8636 25720 8648
rect 25772 8636 25778 8688
rect 25898 8676 25904 8688
rect 25859 8648 25904 8676
rect 25898 8636 25904 8648
rect 25956 8636 25962 8688
rect 28658 8636 28664 8688
rect 28716 8676 28722 8688
rect 28753 8679 28811 8685
rect 28753 8676 28765 8679
rect 28716 8648 28765 8676
rect 28716 8636 28722 8648
rect 28753 8645 28765 8648
rect 28799 8645 28811 8679
rect 28753 8639 28811 8645
rect 400 8586 31680 8608
rect 400 8534 18870 8586
rect 18922 8534 18934 8586
rect 18986 8534 18998 8586
rect 19050 8534 19062 8586
rect 19114 8534 19126 8586
rect 19178 8534 31680 8586
rect 400 8512 31680 8534
rect 690 8432 696 8484
rect 748 8472 754 8484
rect 877 8475 935 8481
rect 877 8472 889 8475
rect 748 8444 889 8472
rect 748 8432 754 8444
rect 877 8441 889 8444
rect 923 8441 935 8475
rect 877 8435 935 8441
rect 1245 8475 1303 8481
rect 1245 8441 1257 8475
rect 1291 8472 1303 8475
rect 1426 8472 1432 8484
rect 1291 8444 1432 8472
rect 1291 8441 1303 8444
rect 1245 8435 1303 8441
rect 1426 8432 1432 8444
rect 1484 8432 1490 8484
rect 3910 8472 3916 8484
rect 3871 8444 3916 8472
rect 3910 8432 3916 8444
rect 3968 8432 3974 8484
rect 17437 8475 17495 8481
rect 17437 8441 17449 8475
rect 17483 8472 17495 8475
rect 17986 8472 17992 8484
rect 17483 8444 17992 8472
rect 17483 8441 17495 8444
rect 17437 8435 17495 8441
rect 17986 8432 17992 8444
rect 18044 8432 18050 8484
rect 26358 8472 26364 8484
rect 26319 8444 26364 8472
rect 26358 8432 26364 8444
rect 26416 8432 26422 8484
rect 27094 8472 27100 8484
rect 27055 8444 27100 8472
rect 27094 8432 27100 8444
rect 27152 8432 27158 8484
rect 28382 8472 28388 8484
rect 28343 8444 28388 8472
rect 28382 8432 28388 8444
rect 28440 8432 28446 8484
rect 29394 8472 29400 8484
rect 29355 8444 29400 8472
rect 29394 8432 29400 8444
rect 29452 8432 29458 8484
rect 30038 8472 30044 8484
rect 29999 8444 30044 8472
rect 30038 8432 30044 8444
rect 30096 8432 30102 8484
rect 2898 8404 2904 8416
rect 1904 8376 2904 8404
rect 1904 8345 1932 8376
rect 2898 8364 2904 8376
rect 2956 8364 2962 8416
rect 3729 8407 3787 8413
rect 3729 8404 3741 8407
rect 3192 8376 3741 8404
rect 1889 8339 1947 8345
rect 1889 8305 1901 8339
rect 1935 8305 1947 8339
rect 1889 8299 1947 8305
rect 2257 8339 2315 8345
rect 2257 8305 2269 8339
rect 2303 8305 2315 8339
rect 2257 8299 2315 8305
rect 1794 8228 1800 8280
rect 1852 8268 1858 8280
rect 2272 8268 2300 8299
rect 2346 8296 2352 8348
rect 2404 8336 2410 8348
rect 3192 8336 3220 8376
rect 3729 8373 3741 8376
rect 3775 8404 3787 8407
rect 4002 8404 4008 8416
rect 3775 8376 4008 8404
rect 3775 8373 3787 8376
rect 3729 8367 3787 8373
rect 4002 8364 4008 8376
rect 4060 8364 4066 8416
rect 4186 8364 4192 8416
rect 4244 8404 4250 8416
rect 5290 8404 5296 8416
rect 4244 8376 5296 8404
rect 4244 8364 4250 8376
rect 5290 8364 5296 8376
rect 5348 8364 5354 8416
rect 9982 8404 9988 8416
rect 7516 8376 9988 8404
rect 2404 8308 3220 8336
rect 2404 8296 2410 8308
rect 3358 8296 3364 8348
rect 3416 8336 3422 8348
rect 3634 8336 3640 8348
rect 3416 8308 3640 8336
rect 3416 8296 3422 8308
rect 3634 8296 3640 8308
rect 3692 8296 3698 8348
rect 5474 8336 5480 8348
rect 5435 8308 5480 8336
rect 5474 8296 5480 8308
rect 5532 8296 5538 8348
rect 6210 8296 6216 8348
rect 6268 8336 6274 8348
rect 7130 8336 7136 8348
rect 6268 8308 7136 8336
rect 6268 8296 6274 8308
rect 7130 8296 7136 8308
rect 7188 8336 7194 8348
rect 7516 8345 7544 8376
rect 9982 8364 9988 8376
rect 10040 8364 10046 8416
rect 11546 8364 11552 8416
rect 11604 8364 11610 8416
rect 17526 8404 17532 8416
rect 17487 8376 17532 8404
rect 17526 8364 17532 8376
rect 17584 8364 17590 8416
rect 19093 8407 19151 8413
rect 19093 8373 19105 8407
rect 19139 8404 19151 8407
rect 24610 8404 24616 8416
rect 19139 8376 24616 8404
rect 19139 8373 19151 8376
rect 19093 8367 19151 8373
rect 21224 8348 21252 8376
rect 22880 8348 22908 8376
rect 24610 8364 24616 8376
rect 24668 8404 24674 8416
rect 24705 8407 24763 8413
rect 24705 8404 24717 8407
rect 24668 8376 24717 8404
rect 24668 8364 24674 8376
rect 24705 8373 24717 8376
rect 24751 8373 24763 8407
rect 24705 8367 24763 8373
rect 26450 8364 26456 8416
rect 26508 8404 26514 8416
rect 27189 8407 27247 8413
rect 27189 8404 27201 8407
rect 26508 8376 27201 8404
rect 26508 8364 26514 8376
rect 27189 8373 27201 8376
rect 27235 8404 27247 8407
rect 27370 8404 27376 8416
rect 27235 8376 27376 8404
rect 27235 8373 27247 8376
rect 27189 8367 27247 8373
rect 27370 8364 27376 8376
rect 27428 8364 27434 8416
rect 7501 8339 7559 8345
rect 7501 8336 7513 8339
rect 7188 8308 7513 8336
rect 7188 8296 7194 8308
rect 7501 8305 7513 8308
rect 7547 8305 7559 8339
rect 7866 8336 7872 8348
rect 7827 8308 7872 8336
rect 7501 8299 7559 8305
rect 7866 8296 7872 8308
rect 7924 8296 7930 8348
rect 7961 8339 8019 8345
rect 7961 8305 7973 8339
rect 8007 8305 8019 8339
rect 7961 8299 8019 8305
rect 5842 8268 5848 8280
rect 1852 8240 2300 8268
rect 5803 8240 5848 8268
rect 1852 8228 1858 8240
rect 5842 8228 5848 8240
rect 5900 8228 5906 8280
rect 6854 8268 6860 8280
rect 6815 8240 6860 8268
rect 6854 8228 6860 8240
rect 6912 8228 6918 8280
rect 6946 8228 6952 8280
rect 7004 8268 7010 8280
rect 7317 8271 7375 8277
rect 7317 8268 7329 8271
rect 7004 8240 7329 8268
rect 7004 8228 7010 8240
rect 7317 8237 7329 8240
rect 7363 8237 7375 8271
rect 7317 8231 7375 8237
rect 785 8203 843 8209
rect 785 8169 797 8203
rect 831 8200 843 8203
rect 966 8200 972 8212
rect 831 8172 972 8200
rect 831 8169 843 8172
rect 785 8163 843 8169
rect 966 8160 972 8172
rect 1024 8200 1030 8212
rect 1702 8200 1708 8212
rect 1024 8172 1708 8200
rect 1024 8160 1030 8172
rect 1702 8160 1708 8172
rect 1760 8160 1766 8212
rect 6394 8160 6400 8212
rect 6452 8200 6458 8212
rect 7884 8200 7912 8296
rect 6452 8172 7912 8200
rect 7976 8200 8004 8299
rect 8786 8296 8792 8348
rect 8844 8336 8850 8348
rect 10810 8336 10816 8348
rect 8844 8308 10816 8336
rect 8844 8296 8850 8308
rect 10810 8296 10816 8308
rect 10868 8296 10874 8348
rect 11178 8336 11184 8348
rect 11139 8308 11184 8336
rect 11178 8296 11184 8308
rect 11236 8296 11242 8348
rect 20930 8336 20936 8348
rect 20891 8308 20936 8336
rect 20930 8296 20936 8308
rect 20988 8296 20994 8348
rect 21206 8336 21212 8348
rect 21119 8308 21212 8336
rect 21206 8296 21212 8308
rect 21264 8296 21270 8348
rect 21758 8336 21764 8348
rect 21719 8308 21764 8336
rect 21758 8296 21764 8308
rect 21816 8296 21822 8348
rect 22862 8336 22868 8348
rect 22775 8308 22868 8336
rect 22862 8296 22868 8308
rect 22920 8296 22926 8348
rect 24334 8296 24340 8348
rect 24392 8336 24398 8348
rect 24429 8339 24487 8345
rect 24429 8336 24441 8339
rect 24392 8308 24441 8336
rect 24392 8296 24398 8308
rect 24429 8305 24441 8308
rect 24475 8336 24487 8339
rect 24518 8336 24524 8348
rect 24475 8308 24524 8336
rect 24475 8305 24487 8308
rect 24429 8299 24487 8305
rect 24518 8296 24524 8308
rect 24576 8296 24582 8348
rect 25346 8296 25352 8348
rect 25404 8336 25410 8348
rect 26637 8339 26695 8345
rect 26637 8336 26649 8339
rect 25404 8308 26649 8336
rect 25404 8296 25410 8308
rect 26637 8305 26649 8308
rect 26683 8336 26695 8339
rect 27462 8336 27468 8348
rect 26683 8308 27468 8336
rect 26683 8305 26695 8308
rect 26637 8299 26695 8305
rect 27462 8296 27468 8308
rect 27520 8296 27526 8348
rect 28661 8339 28719 8345
rect 28661 8336 28673 8339
rect 28400 8308 28673 8336
rect 11454 8228 11460 8280
rect 11512 8268 11518 8280
rect 12561 8271 12619 8277
rect 12561 8268 12573 8271
rect 11512 8240 12573 8268
rect 11512 8228 11518 8240
rect 12561 8237 12573 8240
rect 12607 8268 12619 8271
rect 12650 8268 12656 8280
rect 12607 8240 12656 8268
rect 12607 8237 12619 8240
rect 12561 8231 12619 8237
rect 12650 8228 12656 8240
rect 12708 8228 12714 8280
rect 21485 8271 21543 8277
rect 21485 8237 21497 8271
rect 21531 8237 21543 8271
rect 21485 8231 21543 8237
rect 8602 8200 8608 8212
rect 7976 8172 8608 8200
rect 6452 8160 6458 8172
rect 8602 8160 8608 8172
rect 8660 8160 8666 8212
rect 20562 8160 20568 8212
rect 20620 8200 20626 8212
rect 21500 8200 21528 8231
rect 22034 8228 22040 8280
rect 22092 8268 22098 8280
rect 22773 8271 22831 8277
rect 22773 8268 22785 8271
rect 22092 8240 22785 8268
rect 22092 8228 22098 8240
rect 22773 8237 22785 8240
rect 22819 8268 22831 8271
rect 23506 8268 23512 8280
rect 22819 8240 23512 8268
rect 22819 8237 22831 8240
rect 22773 8231 22831 8237
rect 23506 8228 23512 8240
rect 23564 8228 23570 8280
rect 25898 8228 25904 8280
rect 25956 8268 25962 8280
rect 28400 8268 28428 8308
rect 28661 8305 28673 8308
rect 28707 8336 28719 8339
rect 29210 8336 29216 8348
rect 28707 8308 29216 8336
rect 28707 8305 28719 8308
rect 28661 8299 28719 8305
rect 29210 8296 29216 8308
rect 29268 8336 29274 8348
rect 29949 8339 30007 8345
rect 29949 8336 29961 8339
rect 29268 8308 29961 8336
rect 29268 8296 29274 8308
rect 29949 8305 29961 8308
rect 29995 8305 30007 8339
rect 29949 8299 30007 8305
rect 25956 8240 28428 8268
rect 25956 8228 25962 8240
rect 28566 8228 28572 8280
rect 28624 8268 28630 8280
rect 28845 8271 28903 8277
rect 28845 8268 28857 8271
rect 28624 8240 28857 8268
rect 28624 8228 28630 8240
rect 28845 8237 28857 8240
rect 28891 8237 28903 8271
rect 28845 8231 28903 8237
rect 20620 8172 21528 8200
rect 20620 8160 20626 8172
rect 21574 8160 21580 8212
rect 21632 8200 21638 8212
rect 21669 8203 21727 8209
rect 21669 8200 21681 8203
rect 21632 8172 21681 8200
rect 21632 8160 21638 8172
rect 21669 8169 21681 8172
rect 21715 8169 21727 8203
rect 21669 8163 21727 8169
rect 6118 8092 6124 8144
rect 6176 8132 6182 8144
rect 6213 8135 6271 8141
rect 6213 8132 6225 8135
rect 6176 8104 6225 8132
rect 6176 8092 6182 8104
rect 6213 8101 6225 8104
rect 6259 8132 6271 8135
rect 7038 8132 7044 8144
rect 6259 8104 7044 8132
rect 6259 8101 6271 8104
rect 6213 8095 6271 8101
rect 7038 8092 7044 8104
rect 7096 8092 7102 8144
rect 14306 8092 14312 8144
rect 14364 8132 14370 8144
rect 22052 8132 22080 8228
rect 26177 8203 26235 8209
rect 26177 8169 26189 8203
rect 26223 8200 26235 8203
rect 26634 8200 26640 8212
rect 26223 8172 26640 8200
rect 26223 8169 26235 8172
rect 26177 8163 26235 8169
rect 26634 8160 26640 8172
rect 26692 8160 26698 8212
rect 26913 8203 26971 8209
rect 26913 8169 26925 8203
rect 26959 8200 26971 8203
rect 27646 8200 27652 8212
rect 26959 8172 27652 8200
rect 26959 8169 26971 8172
rect 26913 8163 26971 8169
rect 27646 8160 27652 8172
rect 27704 8160 27710 8212
rect 23046 8132 23052 8144
rect 14364 8104 22080 8132
rect 23007 8104 23052 8132
rect 14364 8092 14370 8104
rect 23046 8092 23052 8104
rect 23104 8092 23110 8144
rect 25070 8132 25076 8144
rect 25031 8104 25076 8132
rect 25070 8092 25076 8104
rect 25128 8092 25134 8144
rect 26545 8135 26603 8141
rect 26545 8101 26557 8135
rect 26591 8132 26603 8135
rect 27278 8132 27284 8144
rect 26591 8104 27284 8132
rect 26591 8101 26603 8104
rect 26545 8095 26603 8101
rect 27278 8092 27284 8104
rect 27336 8092 27342 8144
rect 400 8042 31680 8064
rect 400 7990 3510 8042
rect 3562 7990 3574 8042
rect 3626 7990 3638 8042
rect 3690 7990 3702 8042
rect 3754 7990 3766 8042
rect 3818 7990 31680 8042
rect 400 7968 31680 7990
rect 1702 7888 1708 7940
rect 1760 7928 1766 7940
rect 1889 7931 1947 7937
rect 1889 7928 1901 7931
rect 1760 7900 1901 7928
rect 1760 7888 1766 7900
rect 1889 7897 1901 7900
rect 1935 7897 1947 7931
rect 1889 7891 1947 7897
rect 2349 7931 2407 7937
rect 2349 7897 2361 7931
rect 2395 7928 2407 7931
rect 2898 7928 2904 7940
rect 2395 7900 2904 7928
rect 2395 7897 2407 7900
rect 2349 7891 2407 7897
rect 2898 7888 2904 7900
rect 2956 7888 2962 7940
rect 3358 7928 3364 7940
rect 3319 7900 3364 7928
rect 3358 7888 3364 7900
rect 3416 7888 3422 7940
rect 3637 7931 3695 7937
rect 3637 7897 3649 7931
rect 3683 7928 3695 7931
rect 4002 7928 4008 7940
rect 3683 7900 4008 7928
rect 3683 7897 3695 7900
rect 3637 7891 3695 7897
rect 4002 7888 4008 7900
rect 4060 7888 4066 7940
rect 5290 7928 5296 7940
rect 5251 7900 5296 7928
rect 5290 7888 5296 7900
rect 5348 7888 5354 7940
rect 5753 7931 5811 7937
rect 5753 7897 5765 7931
rect 5799 7928 5811 7931
rect 5842 7928 5848 7940
rect 5799 7900 5848 7928
rect 5799 7897 5811 7900
rect 5753 7891 5811 7897
rect 5842 7888 5848 7900
rect 5900 7888 5906 7940
rect 6210 7928 6216 7940
rect 6171 7900 6216 7928
rect 6210 7888 6216 7900
rect 6268 7888 6274 7940
rect 6394 7928 6400 7940
rect 6355 7900 6400 7928
rect 6394 7888 6400 7900
rect 6452 7888 6458 7940
rect 6581 7931 6639 7937
rect 6581 7897 6593 7931
rect 6627 7928 6639 7931
rect 6854 7928 6860 7940
rect 6627 7900 6860 7928
rect 6627 7897 6639 7900
rect 6581 7891 6639 7897
rect 6854 7888 6860 7900
rect 6912 7888 6918 7940
rect 11178 7928 11184 7940
rect 11139 7900 11184 7928
rect 11178 7888 11184 7900
rect 11236 7888 11242 7940
rect 14306 7928 14312 7940
rect 14267 7900 14312 7928
rect 14306 7888 14312 7900
rect 14364 7888 14370 7940
rect 17345 7931 17403 7937
rect 17345 7897 17357 7931
rect 17391 7928 17403 7931
rect 17434 7928 17440 7940
rect 17391 7900 17440 7928
rect 17391 7897 17403 7900
rect 17345 7891 17403 7897
rect 17434 7888 17440 7900
rect 17492 7888 17498 7940
rect 17805 7931 17863 7937
rect 17805 7897 17817 7931
rect 17851 7928 17863 7931
rect 17986 7928 17992 7940
rect 17851 7900 17992 7928
rect 17851 7897 17863 7900
rect 17805 7891 17863 7897
rect 17986 7888 17992 7900
rect 18044 7888 18050 7940
rect 20841 7931 20899 7937
rect 20841 7897 20853 7931
rect 20887 7928 20899 7931
rect 21206 7928 21212 7940
rect 20887 7900 21212 7928
rect 20887 7897 20899 7900
rect 20841 7891 20899 7897
rect 21206 7888 21212 7900
rect 21264 7888 21270 7940
rect 21393 7931 21451 7937
rect 21393 7897 21405 7931
rect 21439 7928 21451 7931
rect 21574 7928 21580 7940
rect 21439 7900 21580 7928
rect 21439 7897 21451 7900
rect 21393 7891 21451 7897
rect 21574 7888 21580 7900
rect 21632 7888 21638 7940
rect 22405 7931 22463 7937
rect 22405 7897 22417 7931
rect 22451 7928 22463 7931
rect 23046 7928 23052 7940
rect 22451 7900 23052 7928
rect 22451 7897 22463 7900
rect 22405 7891 22463 7897
rect 23046 7888 23052 7900
rect 23104 7888 23110 7940
rect 23966 7888 23972 7940
rect 24024 7928 24030 7940
rect 24245 7931 24303 7937
rect 24245 7928 24257 7931
rect 24024 7900 24257 7928
rect 24024 7888 24030 7900
rect 24245 7897 24257 7900
rect 24291 7928 24303 7931
rect 25530 7928 25536 7940
rect 24291 7900 25536 7928
rect 24291 7897 24303 7900
rect 24245 7891 24303 7897
rect 25530 7888 25536 7900
rect 25588 7888 25594 7940
rect 27462 7888 27468 7940
rect 27520 7928 27526 7940
rect 28293 7931 28351 7937
rect 28293 7928 28305 7931
rect 27520 7900 28305 7928
rect 27520 7888 27526 7900
rect 28293 7897 28305 7900
rect 28339 7897 28351 7931
rect 29210 7928 29216 7940
rect 29171 7900 29216 7928
rect 28293 7891 28351 7897
rect 2165 7795 2223 7801
rect 2165 7761 2177 7795
rect 2211 7792 2223 7795
rect 2346 7792 2352 7804
rect 2211 7764 2352 7792
rect 2211 7761 2223 7764
rect 2165 7755 2223 7761
rect 2346 7752 2352 7764
rect 2404 7752 2410 7804
rect 6872 7792 6900 7888
rect 10810 7820 10816 7872
rect 10868 7860 10874 7872
rect 11365 7863 11423 7869
rect 11365 7860 11377 7863
rect 10868 7832 11377 7860
rect 10868 7820 10874 7832
rect 11365 7829 11377 7832
rect 11411 7829 11423 7863
rect 17452 7860 17480 7888
rect 18173 7863 18231 7869
rect 18173 7860 18185 7863
rect 17452 7832 18185 7860
rect 11365 7823 11423 7829
rect 18173 7829 18185 7832
rect 18219 7829 18231 7863
rect 20930 7860 20936 7872
rect 20891 7832 20936 7860
rect 18173 7823 18231 7829
rect 20930 7820 20936 7832
rect 20988 7820 20994 7872
rect 22773 7863 22831 7869
rect 22773 7829 22785 7863
rect 22819 7860 22831 7863
rect 22862 7860 22868 7872
rect 22819 7832 22868 7860
rect 22819 7829 22831 7832
rect 22773 7823 22831 7829
rect 22862 7820 22868 7832
rect 22920 7820 22926 7872
rect 23506 7860 23512 7872
rect 23467 7832 23512 7860
rect 23506 7820 23512 7832
rect 23564 7820 23570 7872
rect 23782 7860 23788 7872
rect 23743 7832 23788 7860
rect 23782 7820 23788 7832
rect 23840 7820 23846 7872
rect 23874 7820 23880 7872
rect 23932 7860 23938 7872
rect 24794 7860 24800 7872
rect 23932 7832 24800 7860
rect 23932 7820 23938 7832
rect 24794 7820 24800 7832
rect 24852 7860 24858 7872
rect 24852 7832 25116 7860
rect 24852 7820 24858 7832
rect 7222 7792 7228 7804
rect 6872 7764 7228 7792
rect 7222 7752 7228 7764
rect 7280 7792 7286 7804
rect 7409 7795 7467 7801
rect 7409 7792 7421 7795
rect 7280 7764 7421 7792
rect 7280 7752 7286 7764
rect 7409 7761 7421 7764
rect 7455 7761 7467 7795
rect 7409 7755 7467 7761
rect 8602 7752 8608 7804
rect 8660 7792 8666 7804
rect 8789 7795 8847 7801
rect 8789 7792 8801 7795
rect 8660 7764 8801 7792
rect 8660 7752 8666 7764
rect 8789 7761 8801 7764
rect 8835 7761 8847 7795
rect 8789 7755 8847 7761
rect 10350 7752 10356 7804
rect 10408 7792 10414 7804
rect 10905 7795 10963 7801
rect 10905 7792 10917 7795
rect 10408 7764 10917 7792
rect 10408 7752 10414 7764
rect 10905 7761 10917 7764
rect 10951 7792 10963 7795
rect 11546 7792 11552 7804
rect 10951 7764 11552 7792
rect 10951 7761 10963 7764
rect 10905 7755 10963 7761
rect 11546 7752 11552 7764
rect 11604 7752 11610 7804
rect 15597 7795 15655 7801
rect 15597 7792 15609 7795
rect 15060 7764 15609 7792
rect 877 7727 935 7733
rect 877 7693 889 7727
rect 923 7724 935 7727
rect 1150 7724 1156 7736
rect 923 7696 1156 7724
rect 923 7693 935 7696
rect 877 7687 935 7693
rect 1150 7684 1156 7696
rect 1208 7684 1214 7736
rect 7038 7724 7044 7736
rect 6951 7696 7044 7724
rect 7038 7684 7044 7696
rect 7096 7724 7102 7736
rect 7498 7724 7504 7736
rect 7096 7696 7504 7724
rect 7096 7684 7102 7696
rect 7498 7684 7504 7696
rect 7556 7684 7562 7736
rect 12282 7684 12288 7736
rect 12340 7724 12346 7736
rect 13665 7727 13723 7733
rect 13665 7724 13677 7727
rect 12340 7696 13677 7724
rect 12340 7684 12346 7696
rect 13665 7693 13677 7696
rect 13711 7724 13723 7727
rect 14306 7724 14312 7736
rect 13711 7696 14312 7724
rect 13711 7693 13723 7696
rect 13665 7687 13723 7693
rect 14306 7684 14312 7696
rect 14364 7684 14370 7736
rect 14858 7684 14864 7736
rect 14916 7724 14922 7736
rect 15060 7733 15088 7764
rect 15597 7761 15609 7764
rect 15643 7792 15655 7795
rect 15778 7792 15784 7804
rect 15643 7764 15784 7792
rect 15643 7761 15655 7764
rect 15597 7755 15655 7761
rect 15778 7752 15784 7764
rect 15836 7752 15842 7804
rect 23230 7792 23236 7804
rect 17084 7764 17756 7792
rect 23191 7764 23236 7792
rect 15045 7727 15103 7733
rect 15045 7724 15057 7727
rect 14916 7696 15057 7724
rect 14916 7684 14922 7696
rect 15045 7693 15057 7696
rect 15091 7693 15103 7727
rect 15045 7687 15103 7693
rect 15134 7684 15140 7736
rect 15192 7724 15198 7736
rect 17084 7733 17112 7764
rect 17069 7727 17127 7733
rect 17069 7724 17081 7727
rect 15192 7696 17081 7724
rect 15192 7684 15198 7696
rect 17069 7693 17081 7696
rect 17115 7693 17127 7727
rect 17621 7727 17679 7733
rect 17621 7724 17633 7727
rect 17069 7687 17127 7693
rect 17452 7696 17633 7724
rect 1061 7659 1119 7665
rect 1061 7625 1073 7659
rect 1107 7656 1119 7659
rect 1426 7656 1432 7668
rect 1107 7628 1432 7656
rect 1107 7625 1119 7628
rect 1061 7619 1119 7625
rect 1426 7616 1432 7628
rect 1484 7616 1490 7668
rect 7774 7616 7780 7668
rect 7832 7616 7838 7668
rect 8786 7616 8792 7668
rect 8844 7656 8850 7668
rect 10997 7659 11055 7665
rect 10997 7656 11009 7659
rect 8844 7628 11009 7656
rect 8844 7616 8850 7628
rect 10997 7625 11009 7628
rect 11043 7656 11055 7659
rect 11454 7656 11460 7668
rect 11043 7628 11460 7656
rect 11043 7625 11055 7628
rect 10997 7619 11055 7625
rect 11454 7616 11460 7628
rect 11512 7616 11518 7668
rect 13941 7659 13999 7665
rect 13941 7625 13953 7659
rect 13987 7625 13999 7659
rect 15321 7659 15379 7665
rect 13941 7619 13999 7625
rect 14186 7628 14444 7656
rect 1794 7588 1800 7600
rect 1755 7560 1800 7588
rect 1794 7548 1800 7560
rect 1852 7548 1858 7600
rect 5474 7588 5480 7600
rect 5435 7560 5480 7588
rect 5474 7548 5480 7560
rect 5532 7548 5538 7600
rect 6762 7588 6768 7600
rect 6723 7560 6768 7588
rect 6762 7548 6768 7560
rect 6820 7548 6826 7600
rect 6949 7591 7007 7597
rect 6949 7557 6961 7591
rect 6995 7588 7007 7591
rect 7792 7588 7820 7616
rect 13956 7588 13984 7619
rect 14030 7588 14036 7600
rect 6995 7560 7820 7588
rect 13943 7560 14036 7588
rect 6995 7557 7007 7560
rect 6949 7551 7007 7557
rect 14030 7548 14036 7560
rect 14088 7588 14094 7600
rect 14186 7588 14214 7628
rect 14416 7600 14444 7628
rect 15321 7625 15333 7659
rect 15367 7625 15379 7659
rect 17452 7656 17480 7696
rect 17621 7693 17633 7696
rect 17667 7693 17679 7727
rect 17621 7687 17679 7693
rect 15321 7619 15379 7625
rect 16900 7628 17480 7656
rect 17529 7659 17587 7665
rect 14398 7588 14404 7600
rect 14088 7560 14214 7588
rect 14359 7560 14404 7588
rect 14088 7548 14094 7560
rect 14398 7548 14404 7560
rect 14456 7548 14462 7600
rect 14674 7548 14680 7600
rect 14732 7588 14738 7600
rect 15336 7588 15364 7619
rect 15781 7591 15839 7597
rect 15781 7588 15793 7591
rect 14732 7560 15793 7588
rect 14732 7548 14738 7560
rect 15781 7557 15793 7560
rect 15827 7557 15839 7591
rect 15781 7551 15839 7557
rect 16790 7548 16796 7600
rect 16848 7588 16854 7600
rect 16900 7597 16928 7628
rect 17529 7625 17541 7659
rect 17575 7656 17587 7659
rect 17728 7656 17756 7764
rect 23230 7752 23236 7764
rect 23288 7752 23294 7804
rect 24886 7792 24892 7804
rect 23846 7764 24892 7792
rect 21209 7727 21267 7733
rect 21209 7693 21221 7727
rect 21255 7724 21267 7727
rect 21758 7724 21764 7736
rect 21255 7696 21764 7724
rect 21255 7693 21267 7696
rect 21209 7687 21267 7693
rect 21758 7684 21764 7696
rect 21816 7724 21822 7736
rect 22589 7727 22647 7733
rect 22589 7724 22601 7727
rect 21816 7696 22601 7724
rect 21816 7684 21822 7696
rect 22589 7693 22601 7696
rect 22635 7724 22647 7727
rect 22957 7727 23015 7733
rect 22957 7724 22969 7727
rect 22635 7696 22969 7724
rect 22635 7693 22647 7696
rect 22589 7687 22647 7693
rect 22957 7693 22969 7696
rect 23003 7724 23015 7727
rect 23846 7724 23874 7764
rect 24886 7752 24892 7764
rect 24944 7792 24950 7804
rect 25088 7801 25116 7832
rect 25073 7795 25131 7801
rect 24944 7764 25024 7792
rect 24944 7752 24950 7764
rect 24996 7733 25024 7764
rect 25073 7761 25085 7795
rect 25119 7761 25131 7795
rect 25073 7755 25131 7761
rect 23003 7696 23874 7724
rect 24981 7727 25039 7733
rect 23003 7693 23015 7696
rect 22957 7687 23015 7693
rect 24981 7693 24993 7727
rect 25027 7693 25039 7727
rect 24981 7687 25039 7693
rect 25349 7727 25407 7733
rect 25349 7693 25361 7727
rect 25395 7693 25407 7727
rect 25530 7724 25536 7736
rect 25491 7696 25536 7724
rect 25349 7687 25407 7693
rect 17575 7628 17756 7656
rect 17575 7625 17587 7628
rect 17529 7619 17587 7625
rect 23598 7616 23604 7668
rect 23656 7656 23662 7668
rect 23966 7656 23972 7668
rect 23656 7628 23972 7656
rect 23656 7616 23662 7628
rect 23966 7616 23972 7628
rect 24024 7616 24030 7668
rect 24061 7659 24119 7665
rect 24061 7625 24073 7659
rect 24107 7656 24119 7659
rect 24334 7656 24340 7668
rect 24107 7628 24340 7656
rect 24107 7625 24119 7628
rect 24061 7619 24119 7625
rect 24334 7616 24340 7628
rect 24392 7616 24398 7668
rect 24610 7616 24616 7668
rect 24668 7656 24674 7668
rect 25070 7656 25076 7668
rect 24668 7628 25076 7656
rect 24668 7616 24674 7628
rect 25070 7616 25076 7628
rect 25128 7656 25134 7668
rect 25364 7656 25392 7687
rect 25530 7684 25536 7696
rect 25588 7684 25594 7736
rect 28308 7724 28336 7891
rect 29210 7888 29216 7900
rect 29268 7928 29274 7940
rect 29949 7931 30007 7937
rect 29949 7928 29961 7931
rect 29268 7900 29961 7928
rect 29268 7888 29274 7900
rect 29949 7897 29961 7900
rect 29995 7897 30007 7931
rect 29949 7891 30007 7897
rect 30038 7888 30044 7940
rect 30096 7928 30102 7940
rect 30133 7931 30191 7937
rect 30133 7928 30145 7931
rect 30096 7900 30145 7928
rect 30096 7888 30102 7900
rect 30133 7897 30145 7900
rect 30179 7897 30191 7931
rect 30133 7891 30191 7897
rect 28566 7724 28572 7736
rect 28308 7696 28572 7724
rect 28566 7684 28572 7696
rect 28624 7724 28630 7736
rect 29305 7727 29363 7733
rect 29305 7724 29317 7727
rect 28624 7696 29317 7724
rect 28624 7684 28630 7696
rect 29305 7693 29317 7696
rect 29351 7693 29363 7727
rect 29305 7687 29363 7693
rect 28845 7659 28903 7665
rect 28845 7656 28857 7659
rect 25128 7628 25392 7656
rect 28124 7628 28857 7656
rect 25128 7616 25134 7628
rect 28124 7600 28152 7628
rect 28845 7625 28857 7628
rect 28891 7625 28903 7659
rect 28845 7619 28903 7625
rect 16885 7591 16943 7597
rect 16885 7588 16897 7591
rect 16848 7560 16897 7588
rect 16848 7548 16854 7560
rect 16885 7557 16897 7560
rect 16931 7557 16943 7591
rect 20562 7588 20568 7600
rect 20523 7560 20568 7588
rect 16885 7551 16943 7557
rect 20562 7548 20568 7560
rect 20620 7548 20626 7600
rect 28106 7588 28112 7600
rect 28067 7560 28112 7588
rect 28106 7548 28112 7560
rect 28164 7548 28170 7600
rect 400 7498 31680 7520
rect 400 7446 18870 7498
rect 18922 7446 18934 7498
rect 18986 7446 18998 7498
rect 19050 7446 19062 7498
rect 19114 7446 19126 7498
rect 19178 7446 31680 7498
rect 400 7424 31680 7446
rect 6946 7384 6952 7396
rect 6907 7356 6952 7384
rect 6946 7344 6952 7356
rect 7004 7344 7010 7396
rect 7222 7384 7228 7396
rect 7183 7356 7228 7384
rect 7222 7344 7228 7356
rect 7280 7344 7286 7396
rect 7498 7384 7504 7396
rect 7411 7356 7504 7384
rect 7498 7344 7504 7356
rect 7556 7384 7562 7396
rect 8878 7384 8884 7396
rect 7556 7356 8884 7384
rect 7556 7344 7562 7356
rect 8878 7344 8884 7356
rect 8936 7344 8942 7396
rect 23049 7387 23107 7393
rect 23049 7353 23061 7387
rect 23095 7384 23107 7387
rect 23230 7384 23236 7396
rect 23095 7356 23236 7384
rect 23095 7353 23107 7356
rect 23049 7347 23107 7353
rect 23230 7344 23236 7356
rect 23288 7344 23294 7396
rect 24334 7384 24340 7396
rect 24295 7356 24340 7384
rect 24334 7344 24340 7356
rect 24392 7344 24398 7396
rect 24518 7384 24524 7396
rect 24479 7356 24524 7384
rect 24518 7344 24524 7356
rect 24576 7344 24582 7396
rect 24702 7384 24708 7396
rect 24663 7356 24708 7384
rect 24702 7344 24708 7356
rect 24760 7344 24766 7396
rect 24886 7384 24892 7396
rect 24847 7356 24892 7384
rect 24886 7344 24892 7356
rect 24944 7344 24950 7396
rect 5845 7319 5903 7325
rect 5845 7285 5857 7319
rect 5891 7316 5903 7319
rect 5934 7316 5940 7328
rect 5891 7288 5940 7316
rect 5891 7285 5903 7288
rect 5845 7279 5903 7285
rect 5934 7276 5940 7288
rect 5992 7276 5998 7328
rect 6762 7276 6768 7328
rect 6820 7316 6826 7328
rect 7133 7319 7191 7325
rect 7133 7316 7145 7319
rect 6820 7288 7145 7316
rect 6820 7276 6826 7288
rect 7133 7285 7145 7288
rect 7179 7316 7191 7319
rect 8602 7316 8608 7328
rect 7179 7288 8608 7316
rect 7179 7285 7191 7288
rect 7133 7279 7191 7285
rect 8602 7276 8608 7288
rect 8660 7276 8666 7328
rect 18722 7316 18728 7328
rect 18683 7288 18728 7316
rect 18722 7276 18728 7288
rect 18780 7276 18786 7328
rect 23601 7319 23659 7325
rect 23601 7285 23613 7319
rect 23647 7316 23659 7319
rect 23690 7316 23696 7328
rect 23647 7288 23696 7316
rect 23647 7285 23659 7288
rect 23601 7279 23659 7285
rect 23690 7276 23696 7288
rect 23748 7276 23754 7328
rect 26634 7276 26640 7328
rect 26692 7316 26698 7328
rect 26692 7288 26772 7316
rect 26692 7276 26698 7288
rect 3358 7208 3364 7260
rect 3416 7248 3422 7260
rect 3545 7251 3603 7257
rect 3545 7248 3557 7251
rect 3416 7220 3557 7248
rect 3416 7208 3422 7220
rect 3545 7217 3557 7220
rect 3591 7217 3603 7251
rect 5290 7248 5296 7260
rect 5251 7220 5296 7248
rect 3545 7211 3603 7217
rect 5290 7208 5296 7220
rect 5348 7208 5354 7260
rect 5474 7248 5480 7260
rect 5435 7220 5480 7248
rect 5474 7208 5480 7220
rect 5532 7208 5538 7260
rect 12282 7248 12288 7260
rect 12243 7220 12288 7248
rect 12282 7208 12288 7220
rect 12340 7208 12346 7260
rect 14674 7208 14680 7260
rect 14732 7248 14738 7260
rect 14861 7251 14919 7257
rect 14861 7248 14873 7251
rect 14732 7220 14873 7248
rect 14732 7208 14738 7220
rect 14861 7217 14873 7220
rect 14907 7217 14919 7251
rect 14861 7211 14919 7217
rect 14950 7208 14956 7260
rect 15008 7248 15014 7260
rect 15045 7251 15103 7257
rect 15045 7248 15057 7251
rect 15008 7220 15057 7248
rect 15008 7208 15014 7220
rect 15045 7217 15057 7220
rect 15091 7217 15103 7251
rect 15045 7211 15103 7217
rect 17802 7208 17808 7260
rect 17860 7248 17866 7260
rect 17989 7251 18047 7257
rect 17989 7248 18001 7251
rect 17860 7220 18001 7248
rect 17860 7208 17866 7220
rect 17989 7217 18001 7220
rect 18035 7217 18047 7251
rect 18170 7248 18176 7260
rect 18131 7220 18176 7248
rect 17989 7211 18047 7217
rect 18170 7208 18176 7220
rect 18228 7208 18234 7260
rect 18265 7251 18323 7257
rect 18265 7217 18277 7251
rect 18311 7248 18323 7251
rect 18446 7248 18452 7260
rect 18311 7220 18452 7248
rect 18311 7217 18323 7220
rect 18265 7211 18323 7217
rect 18446 7208 18452 7220
rect 18504 7208 18510 7260
rect 23046 7208 23052 7260
rect 23104 7248 23110 7260
rect 26744 7257 26772 7288
rect 28658 7276 28664 7328
rect 28716 7316 28722 7328
rect 28716 7288 29348 7316
rect 28716 7276 28722 7288
rect 23325 7251 23383 7257
rect 23325 7248 23337 7251
rect 23104 7220 23337 7248
rect 23104 7208 23110 7220
rect 23325 7217 23337 7220
rect 23371 7217 23383 7251
rect 23325 7211 23383 7217
rect 26729 7251 26787 7257
rect 26729 7217 26741 7251
rect 26775 7217 26787 7251
rect 26729 7211 26787 7217
rect 28106 7208 28112 7260
rect 28164 7248 28170 7260
rect 29320 7257 29348 7288
rect 28845 7251 28903 7257
rect 28845 7248 28857 7251
rect 28164 7220 28857 7248
rect 28164 7208 28170 7220
rect 28845 7217 28857 7220
rect 28891 7217 28903 7251
rect 28845 7211 28903 7217
rect 29213 7251 29271 7257
rect 29213 7217 29225 7251
rect 29259 7217 29271 7251
rect 29213 7211 29271 7217
rect 29305 7251 29363 7257
rect 29305 7217 29317 7251
rect 29351 7217 29363 7251
rect 29305 7211 29363 7217
rect 3821 7183 3879 7189
rect 3821 7149 3833 7183
rect 3867 7180 3879 7183
rect 3910 7180 3916 7192
rect 3867 7152 3916 7180
rect 3867 7149 3879 7152
rect 3821 7143 3879 7149
rect 3910 7140 3916 7152
rect 3968 7140 3974 7192
rect 26542 7140 26548 7192
rect 26600 7180 26606 7192
rect 26637 7183 26695 7189
rect 26637 7180 26649 7183
rect 26600 7152 26649 7180
rect 26600 7140 26606 7152
rect 26637 7149 26649 7152
rect 26683 7149 26695 7183
rect 26637 7143 26695 7149
rect 27830 7140 27836 7192
rect 27888 7180 27894 7192
rect 28661 7183 28719 7189
rect 28661 7180 28673 7183
rect 27888 7152 28673 7180
rect 27888 7140 27894 7152
rect 28661 7149 28673 7152
rect 28707 7180 28719 7183
rect 28750 7180 28756 7192
rect 28707 7152 28756 7180
rect 28707 7149 28719 7152
rect 28661 7143 28719 7149
rect 28750 7140 28756 7152
rect 28808 7140 28814 7192
rect 28014 7072 28020 7124
rect 28072 7112 28078 7124
rect 29228 7112 29256 7211
rect 29578 7112 29584 7124
rect 28072 7084 29584 7112
rect 28072 7072 28078 7084
rect 29578 7072 29584 7084
rect 29636 7072 29642 7124
rect 7777 7047 7835 7053
rect 7777 7013 7789 7047
rect 7823 7044 7835 7047
rect 8142 7044 8148 7056
rect 7823 7016 8148 7044
rect 7823 7013 7835 7016
rect 7777 7007 7835 7013
rect 8142 7004 8148 7016
rect 8200 7004 8206 7056
rect 11546 7004 11552 7056
rect 11604 7044 11610 7056
rect 12285 7047 12343 7053
rect 12285 7044 12297 7047
rect 11604 7016 12297 7044
rect 11604 7004 11610 7016
rect 12285 7013 12297 7016
rect 12331 7044 12343 7047
rect 12742 7044 12748 7056
rect 12331 7016 12748 7044
rect 12331 7013 12343 7016
rect 12285 7007 12343 7013
rect 12742 7004 12748 7016
rect 12800 7004 12806 7056
rect 15134 7044 15140 7056
rect 15095 7016 15140 7044
rect 15134 7004 15140 7016
rect 15192 7004 15198 7056
rect 20194 7004 20200 7056
rect 20252 7044 20258 7056
rect 20289 7047 20347 7053
rect 20289 7044 20301 7047
rect 20252 7016 20301 7044
rect 20252 7004 20258 7016
rect 20289 7013 20301 7016
rect 20335 7013 20347 7047
rect 20289 7007 20347 7013
rect 20565 7047 20623 7053
rect 20565 7013 20577 7047
rect 20611 7044 20623 7047
rect 20930 7044 20936 7056
rect 20611 7016 20936 7044
rect 20611 7013 20623 7016
rect 20565 7007 20623 7013
rect 20930 7004 20936 7016
rect 20988 7004 20994 7056
rect 26910 7044 26916 7056
rect 26871 7016 26916 7044
rect 26910 7004 26916 7016
rect 26968 7004 26974 7056
rect 28474 7044 28480 7056
rect 28435 7016 28480 7044
rect 28474 7004 28480 7016
rect 28532 7004 28538 7056
rect 400 6954 31680 6976
rect 400 6902 3510 6954
rect 3562 6902 3574 6954
rect 3626 6902 3638 6954
rect 3690 6902 3702 6954
rect 3754 6902 3766 6954
rect 3818 6902 31680 6954
rect 400 6880 31680 6902
rect 3358 6800 3364 6852
rect 3416 6840 3422 6852
rect 3545 6843 3603 6849
rect 3545 6840 3557 6843
rect 3416 6812 3557 6840
rect 3416 6800 3422 6812
rect 3545 6809 3557 6812
rect 3591 6809 3603 6843
rect 3545 6803 3603 6809
rect 3821 6843 3879 6849
rect 3821 6809 3833 6843
rect 3867 6840 3879 6843
rect 4002 6840 4008 6852
rect 3867 6812 4008 6840
rect 3867 6809 3879 6812
rect 3821 6803 3879 6809
rect 2993 6639 3051 6645
rect 2993 6605 3005 6639
rect 3039 6636 3051 6639
rect 3836 6636 3864 6803
rect 4002 6800 4008 6812
rect 4060 6800 4066 6852
rect 4830 6840 4836 6852
rect 4480 6812 4836 6840
rect 4480 6645 4508 6812
rect 4830 6800 4836 6812
rect 4888 6800 4894 6852
rect 5290 6840 5296 6852
rect 5251 6812 5296 6840
rect 5290 6800 5296 6812
rect 5348 6800 5354 6852
rect 5753 6843 5811 6849
rect 5753 6809 5765 6843
rect 5799 6840 5811 6843
rect 5934 6840 5940 6852
rect 5799 6812 5940 6840
rect 5799 6809 5811 6812
rect 5753 6803 5811 6809
rect 5934 6800 5940 6812
rect 5992 6800 5998 6852
rect 6486 6800 6492 6852
rect 6544 6840 6550 6852
rect 7317 6843 7375 6849
rect 7317 6840 7329 6843
rect 6544 6812 7329 6840
rect 6544 6800 6550 6812
rect 7317 6809 7329 6812
rect 7363 6840 7375 6843
rect 7961 6843 8019 6849
rect 7961 6840 7973 6843
rect 7363 6812 7973 6840
rect 7363 6809 7375 6812
rect 7317 6803 7375 6809
rect 7961 6809 7973 6812
rect 8007 6809 8019 6843
rect 8878 6840 8884 6852
rect 7961 6803 8019 6809
rect 8436 6812 8884 6840
rect 7130 6772 7136 6784
rect 7091 6744 7136 6772
rect 7130 6732 7136 6744
rect 7188 6732 7194 6784
rect 7406 6732 7412 6784
rect 7464 6772 7470 6784
rect 7501 6775 7559 6781
rect 7501 6772 7513 6775
rect 7464 6744 7513 6772
rect 7464 6732 7470 6744
rect 7501 6741 7513 6744
rect 7547 6772 7559 6775
rect 8436 6772 8464 6812
rect 7547 6744 8464 6772
rect 7547 6741 7559 6744
rect 7501 6735 7559 6741
rect 4465 6639 4523 6645
rect 4465 6636 4477 6639
rect 3039 6608 3864 6636
rect 4296 6608 4477 6636
rect 3039 6605 3051 6608
rect 2993 6599 3051 6605
rect 3269 6571 3327 6577
rect 3269 6568 3281 6571
rect 2916 6540 3281 6568
rect 2916 6512 2944 6540
rect 3269 6537 3281 6540
rect 3315 6537 3327 6571
rect 3269 6531 3327 6537
rect 2898 6500 2904 6512
rect 2859 6472 2904 6500
rect 2898 6460 2904 6472
rect 2956 6460 2962 6512
rect 3082 6460 3088 6512
rect 3140 6500 3146 6512
rect 3910 6500 3916 6512
rect 3140 6472 3916 6500
rect 3140 6460 3146 6472
rect 3910 6460 3916 6472
rect 3968 6460 3974 6512
rect 4094 6460 4100 6512
rect 4152 6500 4158 6512
rect 4296 6509 4324 6608
rect 4465 6605 4477 6608
rect 4511 6605 4523 6639
rect 7148 6636 7176 6732
rect 8142 6704 8148 6716
rect 8103 6676 8148 6704
rect 8142 6664 8148 6676
rect 8200 6664 8206 6716
rect 8329 6639 8387 6645
rect 8329 6636 8341 6639
rect 7148 6608 8341 6636
rect 4465 6599 4523 6605
rect 8329 6605 8341 6608
rect 8375 6605 8387 6639
rect 8694 6636 8700 6648
rect 8655 6608 8700 6636
rect 8329 6599 8387 6605
rect 8694 6596 8700 6608
rect 8752 6596 8758 6648
rect 8804 6645 8832 6812
rect 8878 6800 8884 6812
rect 8936 6800 8942 6852
rect 11365 6843 11423 6849
rect 11365 6809 11377 6843
rect 11411 6840 11423 6843
rect 12009 6843 12067 6849
rect 12009 6840 12021 6843
rect 11411 6812 12021 6840
rect 11411 6809 11423 6812
rect 11365 6803 11423 6809
rect 12009 6809 12021 6812
rect 12055 6809 12067 6843
rect 12009 6803 12067 6809
rect 11546 6772 11552 6784
rect 11507 6744 11552 6772
rect 11546 6732 11552 6744
rect 11604 6732 11610 6784
rect 8789 6639 8847 6645
rect 8789 6605 8801 6639
rect 8835 6605 8847 6639
rect 11917 6639 11975 6645
rect 11917 6636 11929 6639
rect 8789 6599 8847 6605
rect 8896 6608 11929 6636
rect 4370 6528 4376 6580
rect 4428 6568 4434 6580
rect 4741 6571 4799 6577
rect 4741 6568 4753 6571
rect 4428 6540 4753 6568
rect 4428 6528 4434 6540
rect 4741 6537 4753 6540
rect 4787 6568 4799 6571
rect 5017 6571 5075 6577
rect 5017 6568 5029 6571
rect 4787 6540 5029 6568
rect 4787 6537 4799 6540
rect 4741 6531 4799 6537
rect 5017 6537 5029 6540
rect 5063 6537 5075 6571
rect 5017 6531 5075 6537
rect 5474 6528 5480 6580
rect 5532 6568 5538 6580
rect 5569 6571 5627 6577
rect 5569 6568 5581 6571
rect 5532 6540 5581 6568
rect 5532 6528 5538 6540
rect 5569 6537 5581 6540
rect 5615 6568 5627 6571
rect 6578 6568 6584 6580
rect 5615 6540 6584 6568
rect 5615 6537 5627 6540
rect 5569 6531 5627 6537
rect 6578 6528 6584 6540
rect 6636 6528 6642 6580
rect 6670 6528 6676 6580
rect 6728 6568 6734 6580
rect 8896 6568 8924 6608
rect 11917 6605 11929 6608
rect 11963 6605 11975 6639
rect 12024 6636 12052 6803
rect 12282 6800 12288 6852
rect 12340 6840 12346 6852
rect 12377 6843 12435 6849
rect 12377 6840 12389 6843
rect 12340 6812 12389 6840
rect 12340 6800 12346 6812
rect 12377 6809 12389 6812
rect 12423 6809 12435 6843
rect 12742 6840 12748 6852
rect 12703 6812 12748 6840
rect 12377 6803 12435 6809
rect 12742 6800 12748 6812
rect 12800 6800 12806 6852
rect 14585 6843 14643 6849
rect 14585 6809 14597 6843
rect 14631 6840 14643 6843
rect 15134 6840 15140 6852
rect 14631 6812 15140 6840
rect 14631 6809 14643 6812
rect 14585 6803 14643 6809
rect 15134 6800 15140 6812
rect 15192 6800 15198 6852
rect 15226 6800 15232 6852
rect 15284 6840 15290 6852
rect 15413 6843 15471 6849
rect 15413 6840 15425 6843
rect 15284 6812 15425 6840
rect 15284 6800 15290 6812
rect 15413 6809 15425 6812
rect 15459 6840 15471 6843
rect 18170 6840 18176 6852
rect 15459 6812 18176 6840
rect 15459 6809 15471 6812
rect 15413 6803 15471 6809
rect 18170 6800 18176 6812
rect 18228 6800 18234 6852
rect 18633 6843 18691 6849
rect 18633 6809 18645 6843
rect 18679 6840 18691 6843
rect 18722 6840 18728 6852
rect 18679 6812 18728 6840
rect 18679 6809 18691 6812
rect 18633 6803 18691 6809
rect 18722 6800 18728 6812
rect 18780 6800 18786 6852
rect 23046 6800 23052 6852
rect 23104 6840 23110 6852
rect 23325 6843 23383 6849
rect 23325 6840 23337 6843
rect 23104 6812 23337 6840
rect 23104 6800 23110 6812
rect 23325 6809 23337 6812
rect 23371 6840 23383 6843
rect 24610 6840 24616 6852
rect 23371 6812 24616 6840
rect 23371 6809 23383 6812
rect 23325 6803 23383 6809
rect 17802 6732 17808 6784
rect 17860 6772 17866 6784
rect 17989 6775 18047 6781
rect 17989 6772 18001 6775
rect 17860 6744 18001 6772
rect 17860 6732 17866 6744
rect 17989 6741 18001 6744
rect 18035 6741 18047 6775
rect 17989 6735 18047 6741
rect 19829 6775 19887 6781
rect 19829 6741 19841 6775
rect 19875 6772 19887 6775
rect 23601 6775 23659 6781
rect 19875 6744 21160 6772
rect 19875 6741 19887 6744
rect 19829 6735 19887 6741
rect 12190 6664 12196 6716
rect 12248 6704 12254 6716
rect 13297 6707 13355 6713
rect 13297 6704 13309 6707
rect 12248 6676 13309 6704
rect 12248 6664 12254 6676
rect 13297 6673 13309 6676
rect 13343 6704 13355 6707
rect 13849 6707 13907 6713
rect 13849 6704 13861 6707
rect 13343 6676 13861 6704
rect 13343 6673 13355 6676
rect 13297 6667 13355 6673
rect 13849 6673 13861 6676
rect 13895 6704 13907 6707
rect 13938 6704 13944 6716
rect 13895 6676 13944 6704
rect 13895 6673 13907 6676
rect 13849 6667 13907 6673
rect 13938 6664 13944 6676
rect 13996 6664 14002 6716
rect 19553 6707 19611 6713
rect 19553 6704 19565 6707
rect 19016 6676 19565 6704
rect 13113 6639 13171 6645
rect 13113 6636 13125 6639
rect 12024 6608 13125 6636
rect 11917 6599 11975 6605
rect 13113 6605 13125 6608
rect 13159 6636 13171 6639
rect 13202 6636 13208 6648
rect 13159 6608 13208 6636
rect 13159 6605 13171 6608
rect 13113 6599 13171 6605
rect 6728 6540 8924 6568
rect 6728 6528 6734 6540
rect 11546 6528 11552 6580
rect 11604 6568 11610 6580
rect 11733 6571 11791 6577
rect 11733 6568 11745 6571
rect 11604 6540 11745 6568
rect 11604 6528 11610 6540
rect 11733 6537 11745 6540
rect 11779 6537 11791 6571
rect 11932 6568 11960 6599
rect 13202 6596 13208 6608
rect 13260 6636 13266 6648
rect 13665 6639 13723 6645
rect 13665 6636 13677 6639
rect 13260 6608 13677 6636
rect 13260 6596 13266 6608
rect 13665 6605 13677 6608
rect 13711 6605 13723 6639
rect 15321 6639 15379 6645
rect 15321 6636 15333 6639
rect 13665 6599 13723 6605
rect 14186 6608 15333 6636
rect 12561 6571 12619 6577
rect 12561 6568 12573 6571
rect 11932 6540 12573 6568
rect 11733 6531 11791 6537
rect 12561 6537 12573 6540
rect 12607 6537 12619 6571
rect 12561 6531 12619 6537
rect 4281 6503 4339 6509
rect 4281 6500 4293 6503
rect 4152 6472 4293 6500
rect 4152 6460 4158 6472
rect 4281 6469 4293 6472
rect 4327 6469 4339 6503
rect 4281 6463 4339 6469
rect 10810 6460 10816 6512
rect 10868 6500 10874 6512
rect 14186 6500 14214 6608
rect 15321 6605 15333 6608
rect 15367 6636 15379 6639
rect 15781 6639 15839 6645
rect 15781 6636 15793 6639
rect 15367 6608 15793 6636
rect 15367 6605 15379 6608
rect 15321 6599 15379 6605
rect 15781 6605 15793 6608
rect 15827 6605 15839 6639
rect 15781 6599 15839 6605
rect 18262 6596 18268 6648
rect 18320 6636 18326 6648
rect 19016 6645 19044 6676
rect 19553 6673 19565 6676
rect 19599 6673 19611 6707
rect 19553 6667 19611 6673
rect 20194 6664 20200 6716
rect 20252 6704 20258 6716
rect 20749 6707 20807 6713
rect 20749 6704 20761 6707
rect 20252 6676 20761 6704
rect 20252 6664 20258 6676
rect 20749 6673 20761 6676
rect 20795 6673 20807 6707
rect 20749 6667 20807 6673
rect 21132 6648 21160 6744
rect 23601 6741 23613 6775
rect 23647 6772 23659 6775
rect 23690 6772 23696 6784
rect 23647 6744 23696 6772
rect 23647 6741 23659 6744
rect 23601 6735 23659 6741
rect 23690 6732 23696 6744
rect 23748 6732 23754 6784
rect 24260 6704 24288 6812
rect 24610 6800 24616 6812
rect 24668 6800 24674 6852
rect 24886 6800 24892 6852
rect 24944 6840 24950 6852
rect 27557 6843 27615 6849
rect 27557 6840 27569 6843
rect 24944 6812 27569 6840
rect 24944 6800 24950 6812
rect 27557 6809 27569 6812
rect 27603 6840 27615 6843
rect 28106 6840 28112 6852
rect 27603 6812 28112 6840
rect 27603 6809 27615 6812
rect 27557 6803 27615 6809
rect 28106 6800 28112 6812
rect 28164 6800 28170 6852
rect 28290 6840 28296 6852
rect 28251 6812 28296 6840
rect 28290 6800 28296 6812
rect 28348 6800 28354 6852
rect 25530 6732 25536 6784
rect 25588 6772 25594 6784
rect 26361 6775 26419 6781
rect 26361 6772 26373 6775
rect 25588 6744 26373 6772
rect 25588 6732 25594 6744
rect 26361 6741 26373 6744
rect 26407 6741 26419 6775
rect 26361 6735 26419 6741
rect 26634 6732 26640 6784
rect 26692 6772 26698 6784
rect 26821 6775 26879 6781
rect 26821 6772 26833 6775
rect 26692 6744 26833 6772
rect 26692 6732 26698 6744
rect 26821 6741 26833 6744
rect 26867 6741 26879 6775
rect 26821 6735 26879 6741
rect 26910 6732 26916 6784
rect 26968 6772 26974 6784
rect 27005 6775 27063 6781
rect 27005 6772 27017 6775
rect 26968 6744 27017 6772
rect 26968 6732 26974 6744
rect 27005 6741 27017 6744
rect 27051 6741 27063 6775
rect 27830 6772 27836 6784
rect 27791 6744 27836 6772
rect 27005 6735 27063 6741
rect 27830 6732 27836 6744
rect 27888 6732 27894 6784
rect 27373 6707 27431 6713
rect 27373 6704 27385 6707
rect 24260 6676 27385 6704
rect 27373 6673 27385 6676
rect 27419 6704 27431 6707
rect 28014 6704 28020 6716
rect 27419 6676 28020 6704
rect 27419 6673 27431 6676
rect 27373 6667 27431 6673
rect 28014 6664 28020 6676
rect 28072 6664 28078 6716
rect 28124 6704 28152 6800
rect 28308 6772 28336 6800
rect 28308 6744 29532 6772
rect 28124 6676 29256 6704
rect 29228 6648 29256 6676
rect 29302 6664 29308 6716
rect 29360 6704 29366 6716
rect 29504 6713 29532 6744
rect 29489 6707 29547 6713
rect 29360 6676 29405 6704
rect 29360 6664 29366 6676
rect 29489 6673 29501 6707
rect 29535 6673 29547 6707
rect 29489 6667 29547 6673
rect 19001 6639 19059 6645
rect 19001 6636 19013 6639
rect 18320 6608 19013 6636
rect 18320 6596 18326 6608
rect 19001 6605 19013 6608
rect 19047 6605 19059 6639
rect 19001 6599 19059 6605
rect 19277 6639 19335 6645
rect 19277 6605 19289 6639
rect 19323 6636 19335 6639
rect 20930 6636 20936 6648
rect 19323 6608 20700 6636
rect 20843 6608 20936 6636
rect 19323 6605 19335 6608
rect 19277 6599 19335 6605
rect 14674 6528 14680 6580
rect 14732 6568 14738 6580
rect 14769 6571 14827 6577
rect 14769 6568 14781 6571
rect 14732 6540 14781 6568
rect 14732 6528 14738 6540
rect 14769 6537 14781 6540
rect 14815 6568 14827 6571
rect 15137 6571 15195 6577
rect 15137 6568 15149 6571
rect 14815 6540 15149 6568
rect 14815 6537 14827 6540
rect 14769 6531 14827 6537
rect 15137 6537 15149 6540
rect 15183 6537 15195 6571
rect 15137 6531 15195 6537
rect 14858 6500 14864 6512
rect 10868 6472 14214 6500
rect 14819 6472 14864 6500
rect 10868 6460 10874 6472
rect 14858 6460 14864 6472
rect 14916 6460 14922 6512
rect 15152 6500 15180 6531
rect 15410 6528 15416 6580
rect 15468 6568 15474 6580
rect 18909 6571 18967 6577
rect 15468 6540 18676 6568
rect 15468 6528 15474 6540
rect 16057 6503 16115 6509
rect 16057 6500 16069 6503
rect 15152 6472 16069 6500
rect 16057 6469 16069 6472
rect 16103 6500 16115 6503
rect 16330 6500 16336 6512
rect 16103 6472 16336 6500
rect 16103 6469 16115 6472
rect 16057 6463 16115 6469
rect 16330 6460 16336 6472
rect 16388 6460 16394 6512
rect 18446 6500 18452 6512
rect 18407 6472 18452 6500
rect 18446 6460 18452 6472
rect 18504 6460 18510 6512
rect 18648 6500 18676 6540
rect 18909 6537 18921 6571
rect 18955 6568 18967 6571
rect 19292 6568 19320 6599
rect 20013 6571 20071 6577
rect 18955 6540 19320 6568
rect 19706 6540 19872 6568
rect 18955 6537 18967 6540
rect 18909 6531 18967 6537
rect 19706 6500 19734 6540
rect 18648 6472 19734 6500
rect 19844 6500 19872 6540
rect 20013 6537 20025 6571
rect 20059 6568 20071 6571
rect 20289 6571 20347 6577
rect 20289 6568 20301 6571
rect 20059 6540 20301 6568
rect 20059 6537 20071 6540
rect 20013 6531 20071 6537
rect 20289 6537 20301 6540
rect 20335 6568 20347 6571
rect 20562 6568 20568 6580
rect 20335 6540 20568 6568
rect 20335 6537 20347 6540
rect 20289 6531 20347 6537
rect 20562 6528 20568 6540
rect 20620 6528 20626 6580
rect 20672 6568 20700 6608
rect 20930 6596 20936 6608
rect 20988 6596 20994 6648
rect 21114 6636 21120 6648
rect 21027 6608 21120 6636
rect 21114 6596 21120 6608
rect 21172 6636 21178 6648
rect 21255 6639 21313 6645
rect 21255 6636 21267 6639
rect 21172 6608 21267 6636
rect 21172 6596 21178 6608
rect 21255 6605 21267 6608
rect 21301 6605 21313 6639
rect 21255 6599 21313 6605
rect 21485 6639 21543 6645
rect 21485 6605 21497 6639
rect 21531 6636 21543 6639
rect 21942 6636 21948 6648
rect 21531 6608 21948 6636
rect 21531 6605 21543 6608
rect 21485 6599 21543 6605
rect 21942 6596 21948 6608
rect 22000 6596 22006 6648
rect 23414 6596 23420 6648
rect 23472 6636 23478 6648
rect 23690 6636 23696 6648
rect 23472 6608 23696 6636
rect 23472 6596 23478 6608
rect 23690 6596 23696 6608
rect 23748 6596 23754 6648
rect 24242 6636 24248 6648
rect 24203 6608 24248 6636
rect 24242 6596 24248 6608
rect 24300 6596 24306 6648
rect 24334 6596 24340 6648
rect 24392 6636 24398 6648
rect 24613 6639 24671 6645
rect 24613 6636 24625 6639
rect 24392 6608 24625 6636
rect 24392 6596 24398 6608
rect 24613 6605 24625 6608
rect 24659 6605 24671 6639
rect 24613 6599 24671 6605
rect 25438 6596 25444 6648
rect 25496 6636 25502 6648
rect 26542 6636 26548 6648
rect 25496 6608 26548 6636
rect 25496 6596 25502 6608
rect 26542 6596 26548 6608
rect 26600 6636 26606 6648
rect 26637 6639 26695 6645
rect 26637 6636 26649 6639
rect 26600 6608 26649 6636
rect 26600 6596 26606 6608
rect 26637 6605 26649 6608
rect 26683 6605 26695 6639
rect 29210 6636 29216 6648
rect 29123 6608 29216 6636
rect 26637 6599 26695 6605
rect 29210 6596 29216 6608
rect 29268 6596 29274 6648
rect 29578 6636 29584 6648
rect 29539 6608 29584 6636
rect 29578 6596 29584 6608
rect 29636 6636 29642 6648
rect 29857 6639 29915 6645
rect 29857 6636 29869 6639
rect 29636 6608 29869 6636
rect 29636 6596 29642 6608
rect 29857 6605 29869 6608
rect 29903 6605 29915 6639
rect 29857 6599 29915 6605
rect 20948 6568 20976 6596
rect 21666 6568 21672 6580
rect 20672 6540 21672 6568
rect 21666 6528 21672 6540
rect 21724 6528 21730 6580
rect 23322 6528 23328 6580
rect 23380 6568 23386 6580
rect 28017 6571 28075 6577
rect 23380 6540 24196 6568
rect 23380 6528 23386 6540
rect 20197 6503 20255 6509
rect 20197 6500 20209 6503
rect 19844 6472 20209 6500
rect 20197 6469 20209 6472
rect 20243 6500 20255 6503
rect 20378 6500 20384 6512
rect 20243 6472 20384 6500
rect 20243 6469 20255 6472
rect 20197 6463 20255 6469
rect 20378 6460 20384 6472
rect 20436 6460 20442 6512
rect 21574 6460 21580 6512
rect 21632 6500 21638 6512
rect 22126 6500 22132 6512
rect 21632 6472 22132 6500
rect 21632 6460 21638 6472
rect 22126 6460 22132 6472
rect 22184 6500 22190 6512
rect 23340 6500 23368 6528
rect 22184 6472 23368 6500
rect 22184 6460 22190 6472
rect 23598 6460 23604 6512
rect 23656 6500 23662 6512
rect 24168 6509 24196 6540
rect 23877 6503 23935 6509
rect 23877 6500 23889 6503
rect 23656 6472 23889 6500
rect 23656 6460 23662 6472
rect 23877 6469 23889 6472
rect 23923 6469 23935 6503
rect 23877 6463 23935 6469
rect 24153 6503 24211 6509
rect 24153 6469 24165 6503
rect 24199 6500 24211 6503
rect 24996 6500 25024 6568
rect 28017 6537 28029 6571
rect 28063 6568 28075 6571
rect 28474 6568 28480 6580
rect 28063 6540 28480 6568
rect 28063 6537 28075 6540
rect 28017 6531 28075 6537
rect 28474 6528 28480 6540
rect 28532 6568 28538 6580
rect 28934 6568 28940 6580
rect 28532 6540 28940 6568
rect 28532 6528 28538 6540
rect 28934 6528 28940 6540
rect 28992 6528 28998 6580
rect 24199 6472 25024 6500
rect 28201 6503 28259 6509
rect 24199 6469 24211 6472
rect 24153 6463 24211 6469
rect 28201 6469 28213 6503
rect 28247 6500 28259 6503
rect 28658 6500 28664 6512
rect 28247 6472 28664 6500
rect 28247 6469 28259 6472
rect 28201 6463 28259 6469
rect 28658 6460 28664 6472
rect 28716 6460 28722 6512
rect 28842 6500 28848 6512
rect 28803 6472 28848 6500
rect 28842 6460 28848 6472
rect 28900 6460 28906 6512
rect 400 6410 31680 6432
rect 400 6358 18870 6410
rect 18922 6358 18934 6410
rect 18986 6358 18998 6410
rect 19050 6358 19062 6410
rect 19114 6358 19126 6410
rect 19178 6358 31680 6410
rect 400 6336 31680 6358
rect 874 6296 880 6308
rect 835 6268 880 6296
rect 874 6256 880 6268
rect 932 6256 938 6308
rect 7777 6299 7835 6305
rect 7777 6265 7789 6299
rect 7823 6296 7835 6299
rect 8694 6296 8700 6308
rect 7823 6268 8700 6296
rect 7823 6265 7835 6268
rect 7777 6259 7835 6265
rect 8694 6256 8700 6268
rect 8752 6256 8758 6308
rect 9154 6256 9160 6308
rect 9212 6296 9218 6308
rect 11270 6296 11276 6308
rect 9212 6268 11276 6296
rect 9212 6256 9218 6268
rect 10368 6240 10396 6268
rect 11270 6256 11276 6268
rect 11328 6256 11334 6308
rect 11825 6299 11883 6305
rect 11825 6265 11837 6299
rect 11871 6296 11883 6299
rect 12190 6296 12196 6308
rect 11871 6268 12196 6296
rect 11871 6265 11883 6268
rect 11825 6259 11883 6265
rect 12190 6256 12196 6268
rect 12248 6256 12254 6308
rect 15226 6296 15232 6308
rect 15187 6268 15232 6296
rect 15226 6256 15232 6268
rect 15284 6256 15290 6308
rect 24242 6296 24248 6308
rect 24203 6268 24248 6296
rect 24242 6256 24248 6268
rect 24300 6296 24306 6308
rect 28014 6296 28020 6308
rect 24300 6268 28020 6296
rect 24300 6256 24306 6268
rect 28014 6256 28020 6268
rect 28072 6256 28078 6308
rect 29210 6296 29216 6308
rect 29171 6268 29216 6296
rect 29210 6256 29216 6268
rect 29268 6256 29274 6308
rect 690 6188 696 6240
rect 748 6228 754 6240
rect 1153 6231 1211 6237
rect 1153 6228 1165 6231
rect 748 6200 1165 6228
rect 748 6188 754 6200
rect 1153 6197 1165 6200
rect 1199 6228 1211 6231
rect 3358 6228 3364 6240
rect 1199 6200 3364 6228
rect 1199 6197 1211 6200
rect 1153 6191 1211 6197
rect 3358 6188 3364 6200
rect 3416 6228 3422 6240
rect 3416 6200 3680 6228
rect 3416 6188 3422 6200
rect 1981 6163 2039 6169
rect 1981 6129 1993 6163
rect 2027 6160 2039 6163
rect 3082 6160 3088 6172
rect 2027 6132 3088 6160
rect 2027 6129 2039 6132
rect 1981 6123 2039 6129
rect 3082 6120 3088 6132
rect 3140 6120 3146 6172
rect 3652 6169 3680 6200
rect 4370 6188 4376 6240
rect 4428 6188 4434 6240
rect 10350 6188 10356 6240
rect 10408 6188 10414 6240
rect 21574 6188 21580 6240
rect 21632 6188 21638 6240
rect 29121 6231 29179 6237
rect 29121 6197 29133 6231
rect 29167 6228 29179 6231
rect 29302 6228 29308 6240
rect 29167 6200 29308 6228
rect 29167 6197 29179 6200
rect 29121 6191 29179 6197
rect 29302 6188 29308 6200
rect 29360 6188 29366 6240
rect 3637 6163 3695 6169
rect 3637 6129 3649 6163
rect 3683 6129 3695 6163
rect 6762 6160 6768 6172
rect 6723 6132 6768 6160
rect 3637 6123 3695 6129
rect 6762 6120 6768 6132
rect 6820 6120 6826 6172
rect 9433 6163 9491 6169
rect 9433 6129 9445 6163
rect 9479 6160 9491 6163
rect 9522 6160 9528 6172
rect 9479 6132 9528 6160
rect 9479 6129 9491 6132
rect 9433 6123 9491 6129
rect 9522 6120 9528 6132
rect 9580 6120 9586 6172
rect 13202 6160 13208 6172
rect 13163 6132 13208 6160
rect 13202 6120 13208 6132
rect 13260 6120 13266 6172
rect 14766 6120 14772 6172
rect 14824 6160 14830 6172
rect 15781 6163 15839 6169
rect 15781 6160 15793 6163
rect 14824 6132 15793 6160
rect 14824 6120 14830 6132
rect 15781 6129 15793 6132
rect 15827 6160 15839 6163
rect 15962 6160 15968 6172
rect 15827 6132 15968 6160
rect 15827 6129 15839 6132
rect 15781 6123 15839 6129
rect 15962 6120 15968 6132
rect 16020 6120 16026 6172
rect 16146 6120 16152 6172
rect 16204 6160 16210 6172
rect 18262 6160 18268 6172
rect 16204 6132 18268 6160
rect 16204 6120 16210 6132
rect 18262 6120 18268 6132
rect 18320 6120 18326 6172
rect 19458 6120 19464 6172
rect 19516 6160 19522 6172
rect 19826 6160 19832 6172
rect 19516 6132 19832 6160
rect 19516 6120 19522 6132
rect 19826 6120 19832 6132
rect 19884 6160 19890 6172
rect 20197 6163 20255 6169
rect 20197 6160 20209 6163
rect 19884 6132 20209 6160
rect 19884 6120 19890 6132
rect 20197 6129 20209 6132
rect 20243 6129 20255 6163
rect 20562 6160 20568 6172
rect 20523 6132 20568 6160
rect 20197 6123 20255 6129
rect 20562 6120 20568 6132
rect 20620 6120 20626 6172
rect 26634 6120 26640 6172
rect 26692 6160 26698 6172
rect 27373 6163 27431 6169
rect 27373 6160 27385 6163
rect 26692 6132 27385 6160
rect 26692 6120 26698 6132
rect 27373 6129 27385 6132
rect 27419 6129 27431 6163
rect 27738 6160 27744 6172
rect 27699 6132 27744 6160
rect 27373 6123 27431 6129
rect 27738 6120 27744 6132
rect 27796 6120 27802 6172
rect 28198 6120 28204 6172
rect 28256 6160 28262 6172
rect 28385 6163 28443 6169
rect 28385 6160 28397 6163
rect 28256 6132 28397 6160
rect 28256 6120 28262 6132
rect 28385 6129 28397 6132
rect 28431 6129 28443 6163
rect 28385 6123 28443 6129
rect 785 6095 843 6101
rect 785 6061 797 6095
rect 831 6092 843 6095
rect 1794 6092 1800 6104
rect 831 6064 1800 6092
rect 831 6061 843 6064
rect 785 6055 843 6061
rect 1794 6052 1800 6064
rect 1852 6092 1858 6104
rect 1889 6095 1947 6101
rect 1889 6092 1901 6095
rect 1852 6064 1901 6092
rect 1852 6052 1858 6064
rect 1889 6061 1901 6064
rect 1935 6061 1947 6095
rect 1889 6055 1947 6061
rect 1904 6024 1932 6055
rect 2162 6052 2168 6104
rect 2220 6092 2226 6104
rect 2441 6095 2499 6101
rect 2441 6092 2453 6095
rect 2220 6064 2453 6092
rect 2220 6052 2226 6064
rect 2441 6061 2453 6064
rect 2487 6092 2499 6095
rect 2533 6095 2591 6101
rect 2533 6092 2545 6095
rect 2487 6064 2545 6092
rect 2487 6061 2499 6064
rect 2441 6055 2499 6061
rect 2533 6061 2545 6064
rect 2579 6061 2591 6095
rect 3910 6092 3916 6104
rect 3871 6064 3916 6092
rect 2533 6055 2591 6061
rect 3910 6052 3916 6064
rect 3968 6052 3974 6104
rect 5658 6092 5664 6104
rect 5619 6064 5664 6092
rect 5658 6052 5664 6064
rect 5716 6052 5722 6104
rect 6578 6052 6584 6104
rect 6636 6092 6642 6104
rect 6949 6095 7007 6101
rect 6949 6092 6961 6095
rect 6636 6064 6961 6092
rect 6636 6052 6642 6064
rect 6949 6061 6961 6064
rect 6995 6061 7007 6095
rect 6949 6055 7007 6061
rect 8418 6052 8424 6104
rect 8476 6092 8482 6104
rect 9065 6095 9123 6101
rect 9065 6092 9077 6095
rect 8476 6064 9077 6092
rect 8476 6052 8482 6064
rect 9065 6061 9077 6064
rect 9111 6092 9123 6095
rect 10718 6092 10724 6104
rect 9111 6064 10724 6092
rect 9111 6061 9123 6064
rect 9065 6055 9123 6061
rect 10718 6052 10724 6064
rect 10776 6052 10782 6104
rect 10810 6052 10816 6104
rect 10868 6092 10874 6104
rect 13478 6092 13484 6104
rect 10868 6064 10913 6092
rect 13439 6064 13484 6092
rect 10868 6052 10874 6064
rect 13478 6052 13484 6064
rect 13536 6052 13542 6104
rect 16057 6095 16115 6101
rect 16057 6061 16069 6095
rect 16103 6092 16115 6095
rect 16238 6092 16244 6104
rect 16103 6064 16244 6092
rect 16103 6061 16115 6064
rect 16057 6055 16115 6061
rect 16238 6052 16244 6064
rect 16296 6052 16302 6104
rect 20378 6052 20384 6104
rect 20436 6092 20442 6104
rect 21942 6092 21948 6104
rect 20436 6064 21948 6092
rect 20436 6052 20442 6064
rect 21942 6052 21948 6064
rect 22000 6052 22006 6104
rect 28290 6092 28296 6104
rect 28251 6064 28296 6092
rect 28290 6052 28296 6064
rect 28348 6052 28354 6104
rect 1904 5996 3036 6024
rect 3008 5968 3036 5996
rect 12282 5984 12288 6036
rect 12340 6024 12346 6036
rect 20194 6024 20200 6036
rect 12340 5996 20200 6024
rect 12340 5984 12346 5996
rect 20194 5984 20200 5996
rect 20252 5984 20258 6036
rect 27646 5984 27652 6036
rect 27704 6024 27710 6036
rect 27741 6027 27799 6033
rect 27741 6024 27753 6027
rect 27704 5996 27753 6024
rect 27704 5984 27710 5996
rect 27741 5993 27753 5996
rect 27787 5993 27799 6027
rect 27741 5987 27799 5993
rect 2990 5916 2996 5968
rect 3048 5956 3054 5968
rect 5290 5956 5296 5968
rect 3048 5928 5296 5956
rect 3048 5916 3054 5928
rect 5290 5916 5296 5928
rect 5348 5916 5354 5968
rect 12009 5959 12067 5965
rect 12009 5925 12021 5959
rect 12055 5956 12067 5959
rect 12374 5956 12380 5968
rect 12055 5928 12380 5956
rect 12055 5925 12067 5928
rect 12009 5919 12067 5925
rect 12374 5916 12380 5928
rect 12432 5916 12438 5968
rect 18541 5959 18599 5965
rect 18541 5925 18553 5959
rect 18587 5956 18599 5959
rect 18630 5956 18636 5968
rect 18587 5928 18636 5956
rect 18587 5925 18599 5928
rect 18541 5919 18599 5925
rect 18630 5916 18636 5928
rect 18688 5916 18694 5968
rect 28842 5956 28848 5968
rect 28803 5928 28848 5956
rect 28842 5916 28848 5928
rect 28900 5916 28906 5968
rect 400 5866 31680 5888
rect 400 5814 3510 5866
rect 3562 5814 3574 5866
rect 3626 5814 3638 5866
rect 3690 5814 3702 5866
rect 3754 5814 3766 5866
rect 3818 5814 31680 5866
rect 400 5792 31680 5814
rect 2901 5755 2959 5761
rect 2901 5721 2913 5755
rect 2947 5752 2959 5755
rect 2990 5752 2996 5764
rect 2947 5724 2996 5752
rect 2947 5721 2959 5724
rect 2901 5715 2959 5721
rect 690 5616 696 5628
rect 651 5588 696 5616
rect 690 5576 696 5588
rect 748 5576 754 5628
rect 2717 5619 2775 5625
rect 2717 5585 2729 5619
rect 2763 5616 2775 5619
rect 2916 5616 2944 5715
rect 2990 5712 2996 5724
rect 3048 5712 3054 5764
rect 3082 5712 3088 5764
rect 3140 5752 3146 5764
rect 3910 5752 3916 5764
rect 3140 5724 3185 5752
rect 3871 5724 3916 5752
rect 3140 5712 3146 5724
rect 3910 5712 3916 5724
rect 3968 5712 3974 5764
rect 6946 5712 6952 5764
rect 7004 5752 7010 5764
rect 7041 5755 7099 5761
rect 7041 5752 7053 5755
rect 7004 5724 7053 5752
rect 7004 5712 7010 5724
rect 7041 5721 7053 5724
rect 7087 5752 7099 5755
rect 7501 5755 7559 5761
rect 7501 5752 7513 5755
rect 7087 5724 7513 5752
rect 7087 5721 7099 5724
rect 7041 5715 7099 5721
rect 7501 5721 7513 5724
rect 7547 5721 7559 5755
rect 7501 5715 7559 5721
rect 8145 5755 8203 5761
rect 8145 5721 8157 5755
rect 8191 5752 8203 5755
rect 8237 5755 8295 5761
rect 8237 5752 8249 5755
rect 8191 5724 8249 5752
rect 8191 5721 8203 5724
rect 8145 5715 8203 5721
rect 8237 5721 8249 5724
rect 8283 5752 8295 5755
rect 11546 5752 11552 5764
rect 8283 5724 11552 5752
rect 8283 5721 8295 5724
rect 8237 5715 8295 5721
rect 2763 5588 2944 5616
rect 3545 5619 3603 5625
rect 2763 5585 2775 5588
rect 2717 5579 2775 5585
rect 3545 5585 3557 5619
rect 3591 5616 3603 5619
rect 3928 5616 3956 5712
rect 4005 5619 4063 5625
rect 4005 5616 4017 5619
rect 3591 5588 4017 5616
rect 3591 5585 3603 5588
rect 3545 5579 3603 5585
rect 4005 5585 4017 5588
rect 4051 5585 4063 5619
rect 7516 5616 7544 5715
rect 11546 5712 11552 5724
rect 11604 5712 11610 5764
rect 13202 5752 13208 5764
rect 13163 5724 13208 5752
rect 13202 5712 13208 5724
rect 13260 5712 13266 5764
rect 13757 5755 13815 5761
rect 13757 5721 13769 5755
rect 13803 5752 13815 5755
rect 14125 5755 14183 5761
rect 14125 5752 14137 5755
rect 13803 5724 14137 5752
rect 13803 5721 13815 5724
rect 13757 5715 13815 5721
rect 14125 5721 14137 5724
rect 14171 5752 14183 5755
rect 14674 5752 14680 5764
rect 14171 5724 14680 5752
rect 14171 5721 14183 5724
rect 14125 5715 14183 5721
rect 14674 5712 14680 5724
rect 14732 5712 14738 5764
rect 15778 5752 15784 5764
rect 15739 5724 15784 5752
rect 15778 5712 15784 5724
rect 15836 5712 15842 5764
rect 15962 5752 15968 5764
rect 15923 5724 15968 5752
rect 15962 5712 15968 5724
rect 16020 5712 16026 5764
rect 18262 5752 18268 5764
rect 18223 5724 18268 5752
rect 18262 5712 18268 5724
rect 18320 5712 18326 5764
rect 19826 5752 19832 5764
rect 19787 5724 19832 5752
rect 19826 5712 19832 5724
rect 19884 5712 19890 5764
rect 20105 5755 20163 5761
rect 20105 5721 20117 5755
rect 20151 5752 20163 5755
rect 20562 5752 20568 5764
rect 20151 5724 20568 5752
rect 20151 5721 20163 5724
rect 20105 5715 20163 5721
rect 20562 5712 20568 5724
rect 20620 5712 20626 5764
rect 21114 5712 21120 5764
rect 21172 5752 21178 5764
rect 21850 5752 21856 5764
rect 21172 5724 21856 5752
rect 21172 5712 21178 5724
rect 21850 5712 21856 5724
rect 21908 5712 21914 5764
rect 23877 5755 23935 5761
rect 23877 5721 23889 5755
rect 23923 5752 23935 5755
rect 24242 5752 24248 5764
rect 23923 5724 24248 5752
rect 23923 5721 23935 5724
rect 23877 5715 23935 5721
rect 24242 5712 24248 5724
rect 24300 5712 24306 5764
rect 24705 5755 24763 5761
rect 24705 5721 24717 5755
rect 24751 5752 24763 5755
rect 25438 5752 25444 5764
rect 24751 5724 25444 5752
rect 24751 5721 24763 5724
rect 24705 5715 24763 5721
rect 8418 5684 8424 5696
rect 8379 5656 8424 5684
rect 8418 5644 8424 5656
rect 8476 5644 8482 5696
rect 8605 5687 8663 5693
rect 8605 5653 8617 5687
rect 8651 5684 8663 5687
rect 8651 5656 10488 5684
rect 8651 5653 8663 5656
rect 8605 5647 8663 5653
rect 9706 5616 9712 5628
rect 7516 5588 9712 5616
rect 4005 5579 4063 5585
rect 9706 5576 9712 5588
rect 9764 5616 9770 5628
rect 9893 5619 9951 5625
rect 9893 5616 9905 5619
rect 9764 5588 9905 5616
rect 9764 5576 9770 5588
rect 9893 5585 9905 5588
rect 9939 5585 9951 5619
rect 9893 5579 9951 5585
rect 10460 5616 10488 5656
rect 10534 5644 10540 5696
rect 10592 5684 10598 5696
rect 11454 5684 11460 5696
rect 10592 5656 11460 5684
rect 10592 5644 10598 5656
rect 11454 5644 11460 5656
rect 11512 5684 11518 5696
rect 14858 5684 14864 5696
rect 11512 5656 14864 5684
rect 11512 5644 11518 5656
rect 11181 5619 11239 5625
rect 11181 5616 11193 5619
rect 10460 5588 11193 5616
rect 3361 5551 3419 5557
rect 3361 5517 3373 5551
rect 3407 5548 3419 5551
rect 4462 5548 4468 5560
rect 3407 5520 4468 5548
rect 3407 5517 3419 5520
rect 3361 5511 3419 5517
rect 4462 5508 4468 5520
rect 4520 5508 4526 5560
rect 4646 5548 4652 5560
rect 4607 5520 4652 5548
rect 4646 5508 4652 5520
rect 4704 5508 4710 5560
rect 4830 5548 4836 5560
rect 4743 5520 4836 5548
rect 4830 5508 4836 5520
rect 4888 5548 4894 5560
rect 6670 5548 6676 5560
rect 4888 5520 6676 5548
rect 4888 5508 4894 5520
rect 6670 5508 6676 5520
rect 6728 5508 6734 5560
rect 6762 5508 6768 5560
rect 6820 5548 6826 5560
rect 6857 5551 6915 5557
rect 6857 5548 6869 5551
rect 6820 5520 6869 5548
rect 6820 5508 6826 5520
rect 6857 5517 6869 5520
rect 6903 5548 6915 5551
rect 7409 5551 7467 5557
rect 7409 5548 7421 5551
rect 6903 5520 7421 5548
rect 6903 5517 6915 5520
rect 6857 5511 6915 5517
rect 7409 5517 7421 5520
rect 7455 5548 7467 5551
rect 7498 5548 7504 5560
rect 7455 5520 7504 5548
rect 7455 5517 7467 5520
rect 7409 5511 7467 5517
rect 7498 5508 7504 5520
rect 7556 5548 7562 5560
rect 8237 5551 8295 5557
rect 8237 5548 8249 5551
rect 7556 5520 8249 5548
rect 7556 5508 7562 5520
rect 8237 5517 8249 5520
rect 8283 5517 8295 5551
rect 8237 5511 8295 5517
rect 8973 5551 9031 5557
rect 8973 5517 8985 5551
rect 9019 5548 9031 5551
rect 9246 5548 9252 5560
rect 9019 5520 9252 5548
rect 9019 5517 9031 5520
rect 8973 5511 9031 5517
rect 9246 5508 9252 5520
rect 9304 5548 9310 5560
rect 10074 5548 10080 5560
rect 9304 5520 9936 5548
rect 10035 5520 10080 5548
rect 9304 5508 9310 5520
rect 966 5480 972 5492
rect 927 5452 972 5480
rect 966 5440 972 5452
rect 1024 5440 1030 5492
rect 1426 5440 1432 5492
rect 1484 5440 1490 5492
rect 3729 5483 3787 5489
rect 3729 5449 3741 5483
rect 3775 5480 3787 5483
rect 3775 5452 3956 5480
rect 3775 5449 3787 5452
rect 3729 5443 3787 5449
rect 3928 5412 3956 5452
rect 5658 5440 5664 5492
rect 5716 5480 5722 5492
rect 5934 5480 5940 5492
rect 5716 5452 5940 5480
rect 5716 5440 5722 5452
rect 5934 5440 5940 5452
rect 5992 5480 5998 5492
rect 7225 5483 7283 5489
rect 7225 5480 7237 5483
rect 5992 5452 7237 5480
rect 5992 5440 5998 5452
rect 7225 5449 7237 5452
rect 7271 5480 7283 5483
rect 7869 5483 7927 5489
rect 7869 5480 7881 5483
rect 7271 5452 7881 5480
rect 7271 5449 7283 5452
rect 7225 5443 7283 5449
rect 7869 5449 7881 5452
rect 7915 5449 7927 5483
rect 7869 5443 7927 5449
rect 8789 5483 8847 5489
rect 8789 5449 8801 5483
rect 8835 5480 8847 5483
rect 9433 5483 9491 5489
rect 9433 5480 9445 5483
rect 8835 5452 9445 5480
rect 8835 5449 8847 5452
rect 8789 5443 8847 5449
rect 9433 5449 9445 5452
rect 9479 5480 9491 5483
rect 9522 5480 9528 5492
rect 9479 5452 9528 5480
rect 9479 5449 9491 5452
rect 9433 5443 9491 5449
rect 9522 5440 9528 5452
rect 9580 5440 9586 5492
rect 9908 5480 9936 5520
rect 10074 5508 10080 5520
rect 10132 5508 10138 5560
rect 10350 5508 10356 5560
rect 10408 5548 10414 5560
rect 10460 5557 10488 5588
rect 11181 5585 11193 5588
rect 11227 5616 11239 5619
rect 11227 5588 12788 5616
rect 11227 5585 11239 5588
rect 11181 5579 11239 5585
rect 10445 5551 10503 5557
rect 10445 5548 10457 5551
rect 10408 5520 10457 5548
rect 10408 5508 10414 5520
rect 10445 5517 10457 5520
rect 10491 5517 10503 5551
rect 10445 5511 10503 5517
rect 10537 5551 10595 5557
rect 10537 5517 10549 5551
rect 10583 5548 10595 5551
rect 10810 5548 10816 5560
rect 10583 5520 10816 5548
rect 10583 5517 10595 5520
rect 10537 5511 10595 5517
rect 10552 5480 10580 5511
rect 10810 5508 10816 5520
rect 10868 5508 10874 5560
rect 12190 5548 12196 5560
rect 12151 5520 12196 5548
rect 12190 5508 12196 5520
rect 12248 5508 12254 5560
rect 12374 5548 12380 5560
rect 12335 5520 12380 5548
rect 12374 5508 12380 5520
rect 12432 5508 12438 5560
rect 12760 5557 12788 5588
rect 12852 5557 12880 5656
rect 14858 5644 14864 5656
rect 14916 5644 14922 5696
rect 20378 5684 20384 5696
rect 20339 5656 20384 5684
rect 20378 5644 20384 5656
rect 20436 5644 20442 5696
rect 21574 5684 21580 5696
rect 20580 5656 21580 5684
rect 12926 5576 12932 5628
rect 12984 5616 12990 5628
rect 13570 5616 13576 5628
rect 12984 5588 13576 5616
rect 12984 5576 12990 5588
rect 13570 5576 13576 5588
rect 13628 5616 13634 5628
rect 13849 5619 13907 5625
rect 13849 5616 13861 5619
rect 13628 5588 13861 5616
rect 13628 5576 13634 5588
rect 13849 5585 13861 5588
rect 13895 5616 13907 5619
rect 14493 5619 14551 5625
rect 14493 5616 14505 5619
rect 13895 5588 14505 5616
rect 13895 5585 13907 5588
rect 13849 5579 13907 5585
rect 14493 5585 14505 5588
rect 14539 5585 14551 5619
rect 19366 5616 19372 5628
rect 14493 5579 14551 5585
rect 18556 5588 19372 5616
rect 12745 5551 12803 5557
rect 12745 5517 12757 5551
rect 12791 5517 12803 5551
rect 12745 5511 12803 5517
rect 12837 5551 12895 5557
rect 12837 5517 12849 5551
rect 12883 5517 12895 5551
rect 12837 5511 12895 5517
rect 13941 5551 13999 5557
rect 13941 5517 13953 5551
rect 13987 5548 13999 5551
rect 14582 5548 14588 5560
rect 13987 5520 14588 5548
rect 13987 5517 13999 5520
rect 13941 5511 13999 5517
rect 9908 5452 10580 5480
rect 10902 5440 10908 5492
rect 10960 5480 10966 5492
rect 11365 5483 11423 5489
rect 11365 5480 11377 5483
rect 10960 5452 11377 5480
rect 10960 5440 10966 5452
rect 11365 5449 11377 5452
rect 11411 5480 11423 5483
rect 11733 5483 11791 5489
rect 11733 5480 11745 5483
rect 11411 5452 11745 5480
rect 11411 5449 11423 5452
rect 11365 5443 11423 5449
rect 11733 5449 11745 5452
rect 11779 5449 11791 5483
rect 12760 5480 12788 5511
rect 14582 5508 14588 5520
rect 14640 5548 14646 5560
rect 14677 5551 14735 5557
rect 14677 5548 14689 5551
rect 14640 5520 14689 5548
rect 14640 5508 14646 5520
rect 14677 5517 14689 5520
rect 14723 5517 14735 5551
rect 14677 5511 14735 5517
rect 15597 5551 15655 5557
rect 15597 5517 15609 5551
rect 15643 5548 15655 5551
rect 15778 5548 15784 5560
rect 15643 5520 15784 5548
rect 15643 5517 15655 5520
rect 15597 5511 15655 5517
rect 15778 5508 15784 5520
rect 15836 5508 15842 5560
rect 18556 5480 18584 5588
rect 19366 5576 19372 5588
rect 19424 5576 19430 5628
rect 19458 5576 19464 5628
rect 19516 5616 19522 5628
rect 20289 5619 20347 5625
rect 20289 5616 20301 5619
rect 19516 5588 20301 5616
rect 19516 5576 19522 5588
rect 20289 5585 20301 5588
rect 20335 5616 20347 5619
rect 20580 5616 20608 5656
rect 21574 5644 21580 5656
rect 21632 5644 21638 5696
rect 21666 5644 21672 5696
rect 21724 5684 21730 5696
rect 22129 5687 22187 5693
rect 22129 5684 22141 5687
rect 21724 5656 22141 5684
rect 21724 5644 21730 5656
rect 22129 5653 22141 5656
rect 22175 5653 22187 5687
rect 22129 5647 22187 5653
rect 20335 5588 20608 5616
rect 20335 5585 20347 5588
rect 20289 5579 20347 5585
rect 20654 5576 20660 5628
rect 20712 5616 20718 5628
rect 21761 5619 21819 5625
rect 21761 5616 21773 5619
rect 20712 5588 21773 5616
rect 20712 5576 20718 5588
rect 21761 5585 21773 5588
rect 21807 5616 21819 5619
rect 23414 5616 23420 5628
rect 21807 5588 23420 5616
rect 21807 5585 21819 5588
rect 21761 5579 21819 5585
rect 23414 5576 23420 5588
rect 23472 5576 23478 5628
rect 23969 5619 24027 5625
rect 23969 5585 23981 5619
rect 24015 5616 24027 5619
rect 24720 5616 24748 5715
rect 25438 5712 25444 5724
rect 25496 5712 25502 5764
rect 26453 5755 26511 5761
rect 26453 5721 26465 5755
rect 26499 5752 26511 5755
rect 26634 5752 26640 5764
rect 26499 5724 26640 5752
rect 26499 5721 26511 5724
rect 26453 5715 26511 5721
rect 26634 5712 26640 5724
rect 26692 5712 26698 5764
rect 27557 5755 27615 5761
rect 27557 5721 27569 5755
rect 27603 5752 27615 5755
rect 28290 5752 28296 5764
rect 27603 5724 28296 5752
rect 27603 5721 27615 5724
rect 27557 5715 27615 5721
rect 28290 5712 28296 5724
rect 28348 5712 28354 5764
rect 26174 5644 26180 5696
rect 26232 5684 26238 5696
rect 27738 5684 27744 5696
rect 26232 5656 27744 5684
rect 26232 5644 26238 5656
rect 27738 5644 27744 5656
rect 27796 5684 27802 5696
rect 28017 5687 28075 5693
rect 28017 5684 28029 5687
rect 27796 5656 28029 5684
rect 27796 5644 27802 5656
rect 28017 5653 28029 5656
rect 28063 5653 28075 5687
rect 28198 5684 28204 5696
rect 28159 5656 28204 5684
rect 28017 5647 28075 5653
rect 28198 5644 28204 5656
rect 28256 5644 28262 5696
rect 24015 5588 24748 5616
rect 25901 5619 25959 5625
rect 24015 5585 24027 5588
rect 23969 5579 24027 5585
rect 25901 5585 25913 5619
rect 25947 5616 25959 5619
rect 26634 5616 26640 5628
rect 25947 5588 26640 5616
rect 25947 5585 25959 5588
rect 25901 5579 25959 5585
rect 26634 5576 26640 5588
rect 26692 5616 26698 5628
rect 27833 5619 27891 5625
rect 27833 5616 27845 5619
rect 26692 5588 27845 5616
rect 26692 5576 26698 5588
rect 27833 5585 27845 5588
rect 27879 5585 27891 5619
rect 27833 5579 27891 5585
rect 18725 5551 18783 5557
rect 18725 5548 18737 5551
rect 12760 5452 18584 5480
rect 18648 5520 18737 5548
rect 11733 5443 11791 5449
rect 18648 5424 18676 5520
rect 18725 5517 18737 5520
rect 18771 5548 18783 5551
rect 19277 5551 19335 5557
rect 19277 5548 19289 5551
rect 18771 5520 19289 5548
rect 18771 5517 18783 5520
rect 18725 5511 18783 5517
rect 19277 5517 19289 5520
rect 19323 5517 19335 5551
rect 19277 5511 19335 5517
rect 21206 5508 21212 5560
rect 21264 5548 21270 5560
rect 21301 5551 21359 5557
rect 21301 5548 21313 5551
rect 21264 5520 21313 5548
rect 21264 5508 21270 5520
rect 21301 5517 21313 5520
rect 21347 5517 21359 5551
rect 21301 5511 21359 5517
rect 21485 5551 21543 5557
rect 21485 5517 21497 5551
rect 21531 5548 21543 5551
rect 21666 5548 21672 5560
rect 21531 5520 21672 5548
rect 21531 5517 21543 5520
rect 21485 5511 21543 5517
rect 21666 5508 21672 5520
rect 21724 5508 21730 5560
rect 21850 5548 21856 5560
rect 21811 5520 21856 5548
rect 21850 5508 21856 5520
rect 21908 5508 21914 5560
rect 24061 5551 24119 5557
rect 24061 5517 24073 5551
rect 24107 5548 24119 5551
rect 24107 5520 24840 5548
rect 24107 5517 24119 5520
rect 24061 5511 24119 5517
rect 19001 5483 19059 5489
rect 19001 5449 19013 5483
rect 19047 5480 19059 5483
rect 19553 5483 19611 5489
rect 19553 5480 19565 5483
rect 19047 5452 19565 5480
rect 19047 5449 19059 5452
rect 19001 5443 19059 5449
rect 19292 5424 19320 5452
rect 19553 5449 19565 5452
rect 19599 5480 19611 5483
rect 24076 5480 24104 5511
rect 19599 5452 21068 5480
rect 19599 5449 19611 5452
rect 19553 5443 19611 5449
rect 4554 5412 4560 5424
rect 3928 5384 4560 5412
rect 4554 5372 4560 5384
rect 4612 5372 4618 5424
rect 6578 5412 6584 5424
rect 6539 5384 6584 5412
rect 6578 5372 6584 5384
rect 6636 5372 6642 5424
rect 9154 5412 9160 5424
rect 9115 5384 9160 5412
rect 9154 5372 9160 5384
rect 9212 5372 9218 5424
rect 13478 5412 13484 5424
rect 13391 5384 13484 5412
rect 13478 5372 13484 5384
rect 13536 5412 13542 5424
rect 13846 5412 13852 5424
rect 13536 5384 13852 5412
rect 13536 5372 13542 5384
rect 13846 5372 13852 5384
rect 13904 5412 13910 5424
rect 15134 5412 15140 5424
rect 13904 5384 15140 5412
rect 13904 5372 13910 5384
rect 15134 5372 15140 5384
rect 15192 5372 15198 5424
rect 15229 5415 15287 5421
rect 15229 5381 15241 5415
rect 15275 5412 15287 5415
rect 15410 5412 15416 5424
rect 15275 5384 15416 5412
rect 15275 5381 15287 5384
rect 15229 5375 15287 5381
rect 15410 5372 15416 5384
rect 15468 5372 15474 5424
rect 16238 5412 16244 5424
rect 16199 5384 16244 5412
rect 16238 5372 16244 5384
rect 16296 5372 16302 5424
rect 18541 5415 18599 5421
rect 18541 5381 18553 5415
rect 18587 5412 18599 5415
rect 18630 5412 18636 5424
rect 18587 5384 18636 5412
rect 18587 5381 18599 5384
rect 18541 5375 18599 5381
rect 18630 5372 18636 5384
rect 18688 5372 18694 5424
rect 19274 5372 19280 5424
rect 19332 5372 19338 5424
rect 20654 5412 20660 5424
rect 20615 5384 20660 5412
rect 20654 5372 20660 5384
rect 20712 5372 20718 5424
rect 20930 5412 20936 5424
rect 20891 5384 20936 5412
rect 20930 5372 20936 5384
rect 20988 5372 20994 5424
rect 21040 5412 21068 5452
rect 21960 5452 24104 5480
rect 21960 5412 21988 5452
rect 24812 5424 24840 5520
rect 24886 5508 24892 5560
rect 24944 5548 24950 5560
rect 25625 5551 25683 5557
rect 25625 5548 25637 5551
rect 24944 5520 25637 5548
rect 24944 5508 24950 5520
rect 25625 5517 25637 5520
rect 25671 5548 25683 5551
rect 26177 5551 26235 5557
rect 26177 5548 26189 5551
rect 25671 5520 26189 5548
rect 25671 5517 25683 5520
rect 25625 5511 25683 5517
rect 26177 5517 26189 5520
rect 26223 5517 26235 5551
rect 26177 5511 26235 5517
rect 26542 5508 26548 5560
rect 26600 5548 26606 5560
rect 26913 5551 26971 5557
rect 26913 5548 26925 5551
rect 26600 5520 26925 5548
rect 26600 5508 26606 5520
rect 26913 5517 26925 5520
rect 26959 5548 26971 5551
rect 27649 5551 27707 5557
rect 27649 5548 27661 5551
rect 26959 5520 27661 5548
rect 26959 5517 26971 5520
rect 26913 5511 26971 5517
rect 27649 5517 27661 5520
rect 27695 5517 27707 5551
rect 27649 5511 27707 5517
rect 28569 5551 28627 5557
rect 28569 5517 28581 5551
rect 28615 5517 28627 5551
rect 28569 5511 28627 5517
rect 26821 5483 26879 5489
rect 26821 5449 26833 5483
rect 26867 5480 26879 5483
rect 27094 5480 27100 5492
rect 26867 5452 27100 5480
rect 26867 5449 26879 5452
rect 26821 5443 26879 5449
rect 27094 5440 27100 5452
rect 27152 5480 27158 5492
rect 27189 5483 27247 5489
rect 27189 5480 27201 5483
rect 27152 5452 27201 5480
rect 27152 5440 27158 5452
rect 27189 5449 27201 5452
rect 27235 5480 27247 5483
rect 28198 5480 28204 5492
rect 27235 5452 28204 5480
rect 27235 5449 27247 5452
rect 27189 5443 27247 5449
rect 28198 5440 28204 5452
rect 28256 5440 28262 5492
rect 24794 5412 24800 5424
rect 21040 5384 21988 5412
rect 24755 5384 24800 5412
rect 24794 5372 24800 5384
rect 24852 5372 24858 5424
rect 26910 5372 26916 5424
rect 26968 5412 26974 5424
rect 28584 5412 28612 5511
rect 28750 5440 28756 5492
rect 28808 5480 28814 5492
rect 28845 5483 28903 5489
rect 28845 5480 28857 5483
rect 28808 5452 28857 5480
rect 28808 5440 28814 5452
rect 28845 5449 28857 5452
rect 28891 5480 28903 5483
rect 29302 5480 29308 5492
rect 28891 5452 29308 5480
rect 28891 5449 28903 5452
rect 28845 5443 28903 5449
rect 29302 5440 29308 5452
rect 29360 5440 29366 5492
rect 29121 5415 29179 5421
rect 29121 5412 29133 5415
rect 26968 5384 29133 5412
rect 26968 5372 26974 5384
rect 29121 5381 29133 5384
rect 29167 5381 29179 5415
rect 29121 5375 29179 5381
rect 400 5322 31680 5344
rect 400 5270 18870 5322
rect 18922 5270 18934 5322
rect 18986 5270 18998 5322
rect 19050 5270 19062 5322
rect 19114 5270 19126 5322
rect 19178 5270 31680 5322
rect 400 5248 31680 5270
rect 874 5208 880 5220
rect 835 5180 880 5208
rect 874 5168 880 5180
rect 932 5168 938 5220
rect 1153 5211 1211 5217
rect 1153 5177 1165 5211
rect 1199 5208 1211 5211
rect 1426 5208 1432 5220
rect 1199 5180 1432 5208
rect 1199 5177 1211 5180
rect 1153 5171 1211 5177
rect 1426 5168 1432 5180
rect 1484 5168 1490 5220
rect 3729 5211 3787 5217
rect 3729 5177 3741 5211
rect 3775 5208 3787 5211
rect 4370 5208 4376 5220
rect 3775 5180 4376 5208
rect 3775 5177 3787 5180
rect 3729 5171 3787 5177
rect 4370 5168 4376 5180
rect 4428 5168 4434 5220
rect 9522 5208 9528 5220
rect 9483 5180 9528 5208
rect 9522 5168 9528 5180
rect 9580 5168 9586 5220
rect 9706 5208 9712 5220
rect 9667 5180 9712 5208
rect 9706 5168 9712 5180
rect 9764 5168 9770 5220
rect 20746 5208 20752 5220
rect 16992 5180 20752 5208
rect 785 5143 843 5149
rect 785 5109 797 5143
rect 831 5140 843 5143
rect 966 5140 972 5152
rect 831 5112 972 5140
rect 831 5109 843 5112
rect 785 5103 843 5109
rect 966 5100 972 5112
rect 1024 5140 1030 5152
rect 4097 5143 4155 5149
rect 1024 5112 1472 5140
rect 1024 5100 1030 5112
rect 1444 5081 1472 5112
rect 4097 5109 4109 5143
rect 4143 5140 4155 5143
rect 4830 5140 4836 5152
rect 4143 5112 4836 5140
rect 4143 5109 4155 5112
rect 4097 5103 4155 5109
rect 4830 5100 4836 5112
rect 4888 5100 4894 5152
rect 7869 5143 7927 5149
rect 7869 5109 7881 5143
rect 7915 5140 7927 5143
rect 8142 5140 8148 5152
rect 7915 5112 8148 5140
rect 7915 5109 7927 5112
rect 7869 5103 7927 5109
rect 8142 5100 8148 5112
rect 8200 5140 8206 5152
rect 8200 5112 9016 5140
rect 8200 5100 8206 5112
rect 1429 5075 1487 5081
rect 1429 5041 1441 5075
rect 1475 5072 1487 5075
rect 1610 5072 1616 5084
rect 1475 5044 1616 5072
rect 1475 5041 1487 5044
rect 1429 5035 1487 5041
rect 1610 5032 1616 5044
rect 1668 5032 1674 5084
rect 1889 5075 1947 5081
rect 1889 5041 1901 5075
rect 1935 5072 1947 5075
rect 2162 5072 2168 5084
rect 1935 5044 2168 5072
rect 1935 5041 1947 5044
rect 1889 5035 1947 5041
rect 2162 5032 2168 5044
rect 2220 5032 2226 5084
rect 2257 5075 2315 5081
rect 2257 5041 2269 5075
rect 2303 5072 2315 5075
rect 3266 5072 3272 5084
rect 2303 5044 3272 5072
rect 2303 5041 2315 5044
rect 2257 5035 2315 5041
rect 3266 5032 3272 5044
rect 3324 5032 3330 5084
rect 4002 5032 4008 5084
rect 4060 5072 4066 5084
rect 4649 5075 4707 5081
rect 4649 5072 4661 5075
rect 4060 5044 4661 5072
rect 4060 5032 4066 5044
rect 4649 5041 4661 5044
rect 4695 5072 4707 5075
rect 4738 5072 4744 5084
rect 4695 5044 4744 5072
rect 4695 5041 4707 5044
rect 4649 5035 4707 5041
rect 4738 5032 4744 5044
rect 4796 5032 4802 5084
rect 7314 5072 7320 5084
rect 7275 5044 7320 5072
rect 7314 5032 7320 5044
rect 7372 5032 7378 5084
rect 7498 5072 7504 5084
rect 7459 5044 7504 5072
rect 7498 5032 7504 5044
rect 7556 5032 7562 5084
rect 8988 5081 9016 5112
rect 11270 5100 11276 5152
rect 11328 5100 11334 5152
rect 16882 5100 16888 5152
rect 16940 5140 16946 5152
rect 16992 5149 17020 5180
rect 20746 5168 20752 5180
rect 20804 5168 20810 5220
rect 20930 5208 20936 5220
rect 20891 5180 20936 5208
rect 20930 5168 20936 5180
rect 20988 5208 20994 5220
rect 20988 5180 21712 5208
rect 20988 5168 20994 5180
rect 16977 5143 17035 5149
rect 16977 5140 16989 5143
rect 16940 5112 16989 5140
rect 16940 5100 16946 5112
rect 16977 5109 16989 5112
rect 17023 5109 17035 5143
rect 16977 5103 17035 5109
rect 17618 5100 17624 5152
rect 17676 5140 17682 5152
rect 20654 5140 20660 5152
rect 17676 5112 20660 5140
rect 17676 5100 17682 5112
rect 8973 5075 9031 5081
rect 8973 5041 8985 5075
rect 9019 5072 9031 5075
rect 9798 5072 9804 5084
rect 9019 5044 9804 5072
rect 9019 5041 9031 5044
rect 8973 5035 9031 5041
rect 9798 5032 9804 5044
rect 9856 5032 9862 5084
rect 10902 5072 10908 5084
rect 10863 5044 10908 5072
rect 10902 5032 10908 5044
rect 10960 5032 10966 5084
rect 15410 5072 15416 5084
rect 15371 5044 15416 5072
rect 15410 5032 15416 5044
rect 15468 5032 15474 5084
rect 15597 5075 15655 5081
rect 15597 5041 15609 5075
rect 15643 5041 15655 5075
rect 15870 5072 15876 5084
rect 15831 5044 15876 5072
rect 15597 5035 15655 5041
rect 1978 4964 1984 5016
rect 2036 5004 2042 5016
rect 2346 5004 2352 5016
rect 2036 4976 2352 5004
rect 2036 4964 2042 4976
rect 2346 4964 2352 4976
rect 2404 5004 2410 5016
rect 2898 5004 2904 5016
rect 2404 4976 2904 5004
rect 2404 4964 2410 4976
rect 2898 4964 2904 4976
rect 2956 5004 2962 5016
rect 4189 5007 4247 5013
rect 4189 5004 4201 5007
rect 2956 4976 4201 5004
rect 2956 4964 2962 4976
rect 4189 4973 4201 4976
rect 4235 4973 4247 5007
rect 4189 4967 4247 4973
rect 3358 4896 3364 4948
rect 3416 4936 3422 4948
rect 3821 4939 3879 4945
rect 3821 4936 3833 4939
rect 3416 4908 3833 4936
rect 3416 4896 3422 4908
rect 3821 4905 3833 4908
rect 3867 4936 3879 4939
rect 4002 4936 4008 4948
rect 3867 4908 4008 4936
rect 3867 4905 3879 4908
rect 3821 4899 3879 4905
rect 4002 4896 4008 4908
rect 4060 4896 4066 4948
rect 4204 4936 4232 4967
rect 4554 4964 4560 5016
rect 4612 5004 4618 5016
rect 9154 5004 9160 5016
rect 4612 4976 4657 5004
rect 9115 4976 9160 5004
rect 4612 4964 4618 4976
rect 9154 4964 9160 4976
rect 9212 4964 9218 5016
rect 10537 5007 10595 5013
rect 10537 4973 10549 5007
rect 10583 5004 10595 5007
rect 10718 5004 10724 5016
rect 10583 4976 10724 5004
rect 10583 4973 10595 4976
rect 10537 4967 10595 4973
rect 10718 4964 10724 4976
rect 10776 4964 10782 5016
rect 11454 4964 11460 5016
rect 11512 5004 11518 5016
rect 12285 5007 12343 5013
rect 12285 5004 12297 5007
rect 11512 4976 12297 5004
rect 11512 4964 11518 4976
rect 12285 4973 12297 4976
rect 12331 4973 12343 5007
rect 12285 4967 12343 4973
rect 14674 4964 14680 5016
rect 14732 5004 14738 5016
rect 15612 5004 15640 5035
rect 15870 5032 15876 5044
rect 15928 5032 15934 5084
rect 16149 5075 16207 5081
rect 16149 5041 16161 5075
rect 16195 5041 16207 5075
rect 16330 5072 16336 5084
rect 16388 5081 16394 5084
rect 16300 5044 16336 5072
rect 16149 5035 16207 5041
rect 14732 4976 15640 5004
rect 14732 4964 14738 4976
rect 4646 4936 4652 4948
rect 4204 4908 4652 4936
rect 4646 4896 4652 4908
rect 4704 4896 4710 4948
rect 15318 4896 15324 4948
rect 15376 4936 15382 4948
rect 16164 4936 16192 5035
rect 16330 5032 16336 5044
rect 16388 5035 16400 5081
rect 18354 5072 18360 5084
rect 18315 5044 18360 5072
rect 16388 5032 16394 5035
rect 18354 5032 18360 5044
rect 18412 5032 18418 5084
rect 18740 5081 18768 5112
rect 20654 5100 20660 5112
rect 20712 5100 20718 5152
rect 21114 5100 21120 5152
rect 21172 5140 21178 5152
rect 21684 5149 21712 5180
rect 25254 5168 25260 5220
rect 25312 5208 25318 5220
rect 25806 5208 25812 5220
rect 25312 5180 25812 5208
rect 25312 5168 25318 5180
rect 25806 5168 25812 5180
rect 25864 5168 25870 5220
rect 27646 5208 27652 5220
rect 27607 5180 27652 5208
rect 27646 5168 27652 5180
rect 27704 5168 27710 5220
rect 28750 5168 28756 5220
rect 28808 5208 28814 5220
rect 30501 5211 30559 5217
rect 30501 5208 30513 5211
rect 28808 5180 30513 5208
rect 28808 5168 28814 5180
rect 30501 5177 30513 5180
rect 30547 5177 30559 5211
rect 30501 5171 30559 5177
rect 21209 5143 21267 5149
rect 21209 5140 21221 5143
rect 21172 5112 21221 5140
rect 21172 5100 21178 5112
rect 21209 5109 21221 5112
rect 21255 5109 21267 5143
rect 21209 5103 21267 5109
rect 21669 5143 21727 5149
rect 21669 5109 21681 5143
rect 21715 5140 21727 5143
rect 21758 5140 21764 5152
rect 21715 5112 21764 5140
rect 21715 5109 21727 5112
rect 21669 5103 21727 5109
rect 21758 5100 21764 5112
rect 21816 5100 21822 5152
rect 22126 5100 22132 5152
rect 22184 5100 22190 5152
rect 23414 5140 23420 5152
rect 23375 5112 23420 5140
rect 23414 5100 23420 5112
rect 23472 5140 23478 5152
rect 24426 5140 24432 5152
rect 23472 5112 24432 5140
rect 23472 5100 23478 5112
rect 24426 5100 24432 5112
rect 24484 5100 24490 5152
rect 29118 5100 29124 5152
rect 29176 5100 29182 5152
rect 18725 5075 18783 5081
rect 18725 5041 18737 5075
rect 18771 5041 18783 5075
rect 18725 5035 18783 5041
rect 19826 5032 19832 5084
rect 19884 5072 19890 5084
rect 21390 5072 21396 5084
rect 19884 5044 21396 5072
rect 19884 5032 19890 5044
rect 21390 5032 21396 5044
rect 21448 5032 21454 5084
rect 24242 5072 24248 5084
rect 24203 5044 24248 5072
rect 24242 5032 24248 5044
rect 24300 5032 24306 5084
rect 27094 5072 27100 5084
rect 27055 5044 27100 5072
rect 27094 5032 27100 5044
rect 27152 5032 27158 5084
rect 28014 5032 28020 5084
rect 28072 5072 28078 5084
rect 28385 5075 28443 5081
rect 28385 5072 28397 5075
rect 28072 5044 28397 5072
rect 28072 5032 28078 5044
rect 28385 5041 28397 5044
rect 28431 5041 28443 5075
rect 28385 5035 28443 5041
rect 17066 4964 17072 5016
rect 17124 5004 17130 5016
rect 17897 5007 17955 5013
rect 17897 5004 17909 5007
rect 17124 4976 17909 5004
rect 17124 4964 17130 4976
rect 17897 4973 17909 4976
rect 17943 5004 17955 5007
rect 18538 5004 18544 5016
rect 17943 4976 18544 5004
rect 17943 4973 17955 4976
rect 17897 4967 17955 4973
rect 18538 4964 18544 4976
rect 18596 4964 18602 5016
rect 18630 4964 18636 5016
rect 18688 5004 18694 5016
rect 18817 5007 18875 5013
rect 18817 5004 18829 5007
rect 18688 4976 18829 5004
rect 18688 4964 18694 4976
rect 18817 4973 18829 4976
rect 18863 4973 18875 5007
rect 24426 5004 24432 5016
rect 24387 4976 24432 5004
rect 18817 4967 18875 4973
rect 24426 4964 24432 4976
rect 24484 4964 24490 5016
rect 27278 5004 27284 5016
rect 27239 4976 27284 5004
rect 27278 4964 27284 4976
rect 27336 4964 27342 5016
rect 28753 5007 28811 5013
rect 28753 4973 28765 5007
rect 28799 5004 28811 5007
rect 28934 5004 28940 5016
rect 28799 4976 28940 5004
rect 28799 4973 28811 4976
rect 28753 4967 28811 4973
rect 28934 4964 28940 4976
rect 28992 4964 28998 5016
rect 15376 4908 16192 4936
rect 15376 4896 15382 4908
rect 4462 4828 4468 4880
rect 4520 4868 4526 4880
rect 4833 4871 4891 4877
rect 4833 4868 4845 4871
rect 4520 4840 4845 4868
rect 4520 4828 4526 4840
rect 4833 4837 4845 4840
rect 4879 4868 4891 4871
rect 4922 4868 4928 4880
rect 4879 4840 4928 4868
rect 4879 4837 4891 4840
rect 4833 4831 4891 4837
rect 4922 4828 4928 4840
rect 4980 4828 4986 4880
rect 9985 4871 10043 4877
rect 9985 4837 9997 4871
rect 10031 4868 10043 4871
rect 10074 4868 10080 4880
rect 10031 4840 10080 4868
rect 10031 4837 10043 4840
rect 9985 4831 10043 4837
rect 10074 4828 10080 4840
rect 10132 4868 10138 4880
rect 12374 4868 12380 4880
rect 10132 4840 12380 4868
rect 10132 4828 10138 4840
rect 12374 4828 12380 4840
rect 12432 4828 12438 4880
rect 15134 4828 15140 4880
rect 15192 4868 15198 4880
rect 18262 4868 18268 4880
rect 15192 4840 18268 4868
rect 15192 4828 15198 4840
rect 18262 4828 18268 4840
rect 18320 4868 18326 4880
rect 21025 4871 21083 4877
rect 21025 4868 21037 4871
rect 18320 4840 21037 4868
rect 18320 4828 18326 4840
rect 21025 4837 21037 4840
rect 21071 4868 21083 4871
rect 21206 4868 21212 4880
rect 21071 4840 21212 4868
rect 21071 4837 21083 4840
rect 21025 4831 21083 4837
rect 21206 4828 21212 4840
rect 21264 4828 21270 4880
rect 400 4778 31680 4800
rect 400 4726 3510 4778
rect 3562 4726 3574 4778
rect 3626 4726 3638 4778
rect 3690 4726 3702 4778
rect 3754 4726 3766 4778
rect 3818 4726 31680 4778
rect 400 4704 31680 4726
rect 1610 4664 1616 4676
rect 1571 4636 1616 4664
rect 1610 4624 1616 4636
rect 1668 4624 1674 4676
rect 1889 4667 1947 4673
rect 1889 4633 1901 4667
rect 1935 4664 1947 4667
rect 1978 4664 1984 4676
rect 1935 4636 1984 4664
rect 1935 4633 1947 4636
rect 1889 4627 1947 4633
rect 1978 4624 1984 4636
rect 2036 4624 2042 4676
rect 2073 4667 2131 4673
rect 2073 4633 2085 4667
rect 2119 4664 2131 4667
rect 2162 4664 2168 4676
rect 2119 4636 2168 4664
rect 2119 4633 2131 4636
rect 2073 4627 2131 4633
rect 2162 4624 2168 4636
rect 2220 4624 2226 4676
rect 4738 4664 4744 4676
rect 4699 4636 4744 4664
rect 4738 4624 4744 4636
rect 4796 4624 4802 4676
rect 4922 4664 4928 4676
rect 4883 4636 4928 4664
rect 4922 4624 4928 4636
rect 4980 4624 4986 4676
rect 7498 4664 7504 4676
rect 7459 4636 7504 4664
rect 7498 4624 7504 4636
rect 7556 4624 7562 4676
rect 7777 4667 7835 4673
rect 7777 4633 7789 4667
rect 7823 4664 7835 4667
rect 8142 4664 8148 4676
rect 7823 4636 8148 4664
rect 7823 4633 7835 4636
rect 7777 4627 7835 4633
rect 8142 4624 8148 4636
rect 8200 4624 8206 4676
rect 8789 4667 8847 4673
rect 8789 4633 8801 4667
rect 8835 4664 8847 4667
rect 9154 4664 9160 4676
rect 8835 4636 9160 4664
rect 8835 4633 8847 4636
rect 8789 4627 8847 4633
rect 9154 4624 9160 4636
rect 9212 4624 9218 4676
rect 9525 4667 9583 4673
rect 9525 4633 9537 4667
rect 9571 4664 9583 4667
rect 9706 4664 9712 4676
rect 9571 4636 9712 4664
rect 9571 4633 9583 4636
rect 9525 4627 9583 4633
rect 4554 4556 4560 4608
rect 4612 4596 4618 4608
rect 4649 4599 4707 4605
rect 4649 4596 4661 4599
rect 4612 4568 4661 4596
rect 4612 4556 4618 4568
rect 4649 4565 4661 4568
rect 4695 4596 4707 4599
rect 5934 4596 5940 4608
rect 4695 4568 5940 4596
rect 4695 4565 4707 4568
rect 4649 4559 4707 4565
rect 5934 4556 5940 4568
rect 5992 4556 5998 4608
rect 6305 4463 6363 4469
rect 6305 4429 6317 4463
rect 6351 4460 6363 4463
rect 6578 4460 6584 4472
rect 6351 4432 6584 4460
rect 6351 4429 6363 4432
rect 6305 4423 6363 4429
rect 6578 4420 6584 4432
rect 6636 4420 6642 4472
rect 8881 4463 8939 4469
rect 8881 4429 8893 4463
rect 8927 4460 8939 4463
rect 9540 4460 9568 4627
rect 9706 4624 9712 4636
rect 9764 4624 9770 4676
rect 10442 4624 10448 4676
rect 10500 4664 10506 4676
rect 10721 4667 10779 4673
rect 10721 4664 10733 4667
rect 10500 4636 10733 4664
rect 10500 4624 10506 4636
rect 10721 4633 10733 4636
rect 10767 4633 10779 4667
rect 10902 4664 10908 4676
rect 10863 4636 10908 4664
rect 10721 4627 10779 4633
rect 10902 4624 10908 4636
rect 10960 4624 10966 4676
rect 11270 4624 11276 4676
rect 11328 4664 11334 4676
rect 11914 4664 11920 4676
rect 11328 4636 11920 4664
rect 11328 4624 11334 4636
rect 11914 4624 11920 4636
rect 11972 4624 11978 4676
rect 15318 4664 15324 4676
rect 14186 4636 15324 4664
rect 9798 4596 9804 4608
rect 9759 4568 9804 4596
rect 9798 4556 9804 4568
rect 9856 4556 9862 4608
rect 10534 4556 10540 4608
rect 10592 4596 10598 4608
rect 14186 4596 14214 4636
rect 15318 4624 15324 4636
rect 15376 4624 15382 4676
rect 15870 4664 15876 4676
rect 15831 4636 15876 4664
rect 15870 4624 15876 4636
rect 15928 4664 15934 4676
rect 16425 4667 16483 4673
rect 16425 4664 16437 4667
rect 15928 4636 16437 4664
rect 15928 4624 15934 4636
rect 16425 4633 16437 4636
rect 16471 4664 16483 4667
rect 16609 4667 16667 4673
rect 16609 4664 16621 4667
rect 16471 4636 16621 4664
rect 16471 4633 16483 4636
rect 16425 4627 16483 4633
rect 16609 4633 16621 4636
rect 16655 4633 16667 4667
rect 16882 4664 16888 4676
rect 16843 4636 16888 4664
rect 16609 4627 16667 4633
rect 16882 4624 16888 4636
rect 16940 4624 16946 4676
rect 17437 4667 17495 4673
rect 17437 4633 17449 4667
rect 17483 4664 17495 4667
rect 18630 4664 18636 4676
rect 17483 4636 18636 4664
rect 17483 4633 17495 4636
rect 17437 4627 17495 4633
rect 18630 4624 18636 4636
rect 18688 4624 18694 4676
rect 18722 4624 18728 4676
rect 18780 4664 18786 4676
rect 21206 4664 21212 4676
rect 18780 4636 21212 4664
rect 18780 4624 18786 4636
rect 21206 4624 21212 4636
rect 21264 4624 21270 4676
rect 21758 4664 21764 4676
rect 21719 4636 21764 4664
rect 21758 4624 21764 4636
rect 21816 4624 21822 4676
rect 24242 4664 24248 4676
rect 24203 4636 24248 4664
rect 24242 4624 24248 4636
rect 24300 4624 24306 4676
rect 27094 4664 27100 4676
rect 27055 4636 27100 4664
rect 27094 4624 27100 4636
rect 27152 4624 27158 4676
rect 28934 4664 28940 4676
rect 28895 4636 28940 4664
rect 28934 4624 28940 4636
rect 28992 4624 28998 4676
rect 14582 4596 14588 4608
rect 10592 4568 14214 4596
rect 14543 4568 14588 4596
rect 10592 4556 10598 4568
rect 14582 4556 14588 4568
rect 14640 4556 14646 4608
rect 14674 4556 14680 4608
rect 14732 4596 14738 4608
rect 14732 4568 14777 4596
rect 14732 4556 14738 4568
rect 15226 4556 15232 4608
rect 15284 4596 15290 4608
rect 15413 4599 15471 4605
rect 15413 4596 15425 4599
rect 15284 4568 15425 4596
rect 15284 4556 15290 4568
rect 15413 4565 15425 4568
rect 15459 4596 15471 4599
rect 16241 4599 16299 4605
rect 16241 4596 16253 4599
rect 15459 4568 16253 4596
rect 15459 4565 15471 4568
rect 15413 4559 15471 4565
rect 16241 4565 16253 4568
rect 16287 4565 16299 4599
rect 17618 4596 17624 4608
rect 17579 4568 17624 4596
rect 16241 4559 16299 4565
rect 17618 4556 17624 4568
rect 17676 4556 17682 4608
rect 18170 4596 18176 4608
rect 18131 4568 18176 4596
rect 18170 4556 18176 4568
rect 18228 4556 18234 4608
rect 18538 4556 18544 4608
rect 18596 4596 18602 4608
rect 19185 4599 19243 4605
rect 19185 4596 19197 4599
rect 18596 4568 19197 4596
rect 18596 4556 18602 4568
rect 19185 4565 19197 4568
rect 19231 4565 19243 4599
rect 19185 4559 19243 4565
rect 20654 4556 20660 4608
rect 20712 4596 20718 4608
rect 21577 4599 21635 4605
rect 21577 4596 21589 4599
rect 20712 4568 21589 4596
rect 20712 4556 20718 4568
rect 21577 4565 21589 4568
rect 21623 4565 21635 4599
rect 21577 4559 21635 4565
rect 10629 4531 10687 4537
rect 10629 4497 10641 4531
rect 10675 4528 10687 4531
rect 11086 4528 11092 4540
rect 10675 4500 11092 4528
rect 10675 4497 10687 4500
rect 10629 4491 10687 4497
rect 11086 4488 11092 4500
rect 11144 4528 11150 4540
rect 11914 4528 11920 4540
rect 11144 4500 11920 4528
rect 11144 4488 11150 4500
rect 11914 4488 11920 4500
rect 11972 4488 11978 4540
rect 13665 4531 13723 4537
rect 13665 4497 13677 4531
rect 13711 4528 13723 4531
rect 14398 4528 14404 4540
rect 13711 4500 14404 4528
rect 13711 4497 13723 4500
rect 13665 4491 13723 4497
rect 14398 4488 14404 4500
rect 14456 4488 14462 4540
rect 19001 4531 19059 4537
rect 19001 4528 19013 4531
rect 18372 4500 19013 4528
rect 18372 4472 18400 4500
rect 19001 4497 19013 4500
rect 19047 4497 19059 4531
rect 19001 4491 19059 4497
rect 21114 4488 21120 4540
rect 21172 4528 21178 4540
rect 21390 4528 21396 4540
rect 21172 4500 21396 4528
rect 21172 4488 21178 4500
rect 21390 4488 21396 4500
rect 21448 4528 21454 4540
rect 21945 4531 22003 4537
rect 21945 4528 21957 4531
rect 21448 4500 21957 4528
rect 21448 4488 21454 4500
rect 21945 4497 21957 4500
rect 21991 4497 22003 4531
rect 21945 4491 22003 4497
rect 8927 4432 9568 4460
rect 8927 4429 8939 4432
rect 8881 4423 8939 4429
rect 10166 4420 10172 4472
rect 10224 4460 10230 4472
rect 12282 4460 12288 4472
rect 10224 4432 12288 4460
rect 10224 4420 10230 4432
rect 12282 4420 12288 4432
rect 12340 4420 12346 4472
rect 13757 4463 13815 4469
rect 13757 4429 13769 4463
rect 13803 4460 13815 4463
rect 14490 4460 14496 4472
rect 13803 4432 14496 4460
rect 13803 4429 13815 4432
rect 13757 4423 13815 4429
rect 14490 4420 14496 4432
rect 14548 4420 14554 4472
rect 15137 4463 15195 4469
rect 15137 4429 15149 4463
rect 15183 4460 15195 4463
rect 15183 4432 15640 4460
rect 15183 4429 15195 4432
rect 15137 4423 15195 4429
rect 6121 4395 6179 4401
rect 6121 4392 6133 4395
rect 4526 4364 6133 4392
rect 1521 4327 1579 4333
rect 1521 4293 1533 4327
rect 1567 4324 1579 4327
rect 3266 4324 3272 4336
rect 1567 4296 3272 4324
rect 1567 4293 1579 4296
rect 1521 4287 1579 4293
rect 3266 4284 3272 4296
rect 3324 4324 3330 4336
rect 4526 4324 4554 4364
rect 6121 4361 6133 4364
rect 6167 4392 6179 4395
rect 6765 4395 6823 4401
rect 6765 4392 6777 4395
rect 6167 4364 6777 4392
rect 6167 4361 6179 4364
rect 6121 4355 6179 4361
rect 6765 4361 6777 4364
rect 6811 4361 6823 4395
rect 6765 4355 6823 4361
rect 8970 4352 8976 4404
rect 9028 4392 9034 4404
rect 9157 4395 9215 4401
rect 9157 4392 9169 4395
rect 9028 4364 9169 4392
rect 9028 4352 9034 4364
rect 9157 4361 9169 4364
rect 9203 4392 9215 4395
rect 9709 4395 9767 4401
rect 9709 4392 9721 4395
rect 9203 4364 9721 4392
rect 9203 4361 9215 4364
rect 9157 4355 9215 4361
rect 9709 4361 9721 4364
rect 9755 4392 9767 4395
rect 11730 4392 11736 4404
rect 9755 4364 11736 4392
rect 9755 4361 9767 4364
rect 9709 4355 9767 4361
rect 11730 4352 11736 4364
rect 11788 4352 11794 4404
rect 15612 4401 15640 4432
rect 15686 4420 15692 4472
rect 15744 4460 15750 4472
rect 15744 4432 15789 4460
rect 15744 4420 15750 4432
rect 16054 4420 16060 4472
rect 16112 4460 16118 4472
rect 18354 4460 18360 4472
rect 16112 4432 18360 4460
rect 16112 4420 16118 4432
rect 18354 4420 18360 4432
rect 18412 4420 18418 4472
rect 18541 4463 18599 4469
rect 18541 4429 18553 4463
rect 18587 4460 18599 4463
rect 18630 4460 18636 4472
rect 18587 4432 18636 4460
rect 18587 4429 18599 4432
rect 18541 4423 18599 4429
rect 14217 4395 14275 4401
rect 14217 4392 14229 4395
rect 13496 4364 14229 4392
rect 3324 4296 4554 4324
rect 5937 4327 5995 4333
rect 3324 4284 3330 4296
rect 5937 4293 5949 4327
rect 5983 4324 5995 4327
rect 6394 4324 6400 4336
rect 5983 4296 6400 4324
rect 5983 4293 5995 4296
rect 5937 4287 5995 4293
rect 6394 4284 6400 4296
rect 6452 4284 6458 4336
rect 6578 4284 6584 4336
rect 6636 4324 6642 4336
rect 7041 4327 7099 4333
rect 7041 4324 7053 4327
rect 6636 4296 7053 4324
rect 6636 4284 6642 4296
rect 7041 4293 7053 4296
rect 7087 4324 7099 4327
rect 7130 4324 7136 4336
rect 7087 4296 7136 4324
rect 7087 4293 7099 4296
rect 7041 4287 7099 4293
rect 7130 4284 7136 4296
rect 7188 4284 7194 4336
rect 7314 4284 7320 4336
rect 7372 4324 7378 4336
rect 7409 4327 7467 4333
rect 7409 4324 7421 4327
rect 7372 4296 7421 4324
rect 7372 4284 7378 4296
rect 7409 4293 7421 4296
rect 7455 4324 7467 4327
rect 7498 4324 7504 4336
rect 7455 4296 7504 4324
rect 7455 4293 7467 4296
rect 7409 4287 7467 4293
rect 7498 4284 7504 4296
rect 7556 4284 7562 4336
rect 10718 4284 10724 4336
rect 10776 4324 10782 4336
rect 11178 4324 11184 4336
rect 10776 4296 11184 4324
rect 10776 4284 10782 4296
rect 11178 4284 11184 4296
rect 11236 4284 11242 4336
rect 13386 4284 13392 4336
rect 13444 4324 13450 4336
rect 13496 4333 13524 4364
rect 14217 4361 14229 4364
rect 14263 4361 14275 4395
rect 14217 4355 14275 4361
rect 14953 4395 15011 4401
rect 14953 4361 14965 4395
rect 14999 4392 15011 4395
rect 15597 4395 15655 4401
rect 14999 4364 15548 4392
rect 14999 4361 15011 4364
rect 14953 4355 15011 4361
rect 13481 4327 13539 4333
rect 13481 4324 13493 4327
rect 13444 4296 13493 4324
rect 13444 4284 13450 4296
rect 13481 4293 13493 4296
rect 13527 4293 13539 4327
rect 14398 4324 14404 4336
rect 14311 4296 14404 4324
rect 13481 4287 13539 4293
rect 14398 4284 14404 4296
rect 14456 4324 14462 4336
rect 15042 4324 15048 4336
rect 14456 4296 15048 4324
rect 14456 4284 14462 4296
rect 15042 4284 15048 4296
rect 15100 4284 15106 4336
rect 15520 4324 15548 4364
rect 15597 4361 15609 4395
rect 15643 4392 15655 4395
rect 17161 4395 17219 4401
rect 17161 4392 17173 4395
rect 15643 4364 17173 4392
rect 15643 4361 15655 4364
rect 15597 4355 15655 4361
rect 17161 4361 17173 4364
rect 17207 4392 17219 4395
rect 18556 4392 18584 4423
rect 18630 4420 18636 4432
rect 18688 4420 18694 4472
rect 18725 4463 18783 4469
rect 18725 4429 18737 4463
rect 18771 4429 18783 4463
rect 18725 4423 18783 4429
rect 17207 4364 18584 4392
rect 17207 4361 17219 4364
rect 17161 4355 17219 4361
rect 16330 4324 16336 4336
rect 15520 4296 16336 4324
rect 16330 4284 16336 4296
rect 16388 4284 16394 4336
rect 17805 4327 17863 4333
rect 17805 4293 17817 4327
rect 17851 4324 17863 4327
rect 18740 4324 18768 4423
rect 28014 4420 28020 4472
rect 28072 4460 28078 4472
rect 29121 4463 29179 4469
rect 29121 4460 29133 4463
rect 28072 4432 29133 4460
rect 28072 4420 28078 4432
rect 29121 4429 29133 4432
rect 29167 4429 29179 4463
rect 29121 4423 29179 4429
rect 20562 4352 20568 4404
rect 20620 4392 20626 4404
rect 28750 4392 28756 4404
rect 20620 4364 28756 4392
rect 20620 4352 20626 4364
rect 28750 4352 28756 4364
rect 28808 4352 28814 4404
rect 21022 4324 21028 4336
rect 17851 4296 21028 4324
rect 17851 4293 17863 4296
rect 17805 4287 17863 4293
rect 21022 4284 21028 4296
rect 21080 4284 21086 4336
rect 21485 4327 21543 4333
rect 21485 4293 21497 4327
rect 21531 4324 21543 4327
rect 21574 4324 21580 4336
rect 21531 4296 21580 4324
rect 21531 4293 21543 4296
rect 21485 4287 21543 4293
rect 21574 4284 21580 4296
rect 21632 4284 21638 4336
rect 24058 4284 24064 4336
rect 24116 4324 24122 4336
rect 24426 4324 24432 4336
rect 24116 4296 24432 4324
rect 24116 4284 24122 4296
rect 24426 4284 24432 4296
rect 24484 4284 24490 4336
rect 27278 4324 27284 4336
rect 27239 4296 27284 4324
rect 27278 4284 27284 4296
rect 27336 4284 27342 4336
rect 28658 4324 28664 4336
rect 28619 4296 28664 4324
rect 28658 4284 28664 4296
rect 28716 4284 28722 4336
rect 400 4234 31680 4256
rect 400 4182 18870 4234
rect 18922 4182 18934 4234
rect 18986 4182 18998 4234
rect 19050 4182 19062 4234
rect 19114 4182 19126 4234
rect 19178 4182 31680 4234
rect 400 4160 31680 4182
rect 1242 4120 1248 4132
rect 1203 4092 1248 4120
rect 1242 4080 1248 4092
rect 1300 4080 1306 4132
rect 6394 4080 6400 4132
rect 6452 4120 6458 4132
rect 9430 4120 9436 4132
rect 6452 4092 9436 4120
rect 6452 4080 6458 4092
rect 9430 4080 9436 4092
rect 9488 4120 9494 4132
rect 10994 4120 11000 4132
rect 9488 4092 11000 4120
rect 9488 4080 9494 4092
rect 10994 4080 11000 4092
rect 11052 4080 11058 4132
rect 13846 4120 13852 4132
rect 13807 4092 13852 4120
rect 13846 4080 13852 4092
rect 13904 4080 13910 4132
rect 15410 4080 15416 4132
rect 15468 4120 15474 4132
rect 15597 4123 15655 4129
rect 15597 4120 15609 4123
rect 15468 4092 15609 4120
rect 15468 4080 15474 4092
rect 15597 4089 15609 4092
rect 15643 4089 15655 4123
rect 15597 4083 15655 4089
rect 18170 4080 18176 4132
rect 18228 4120 18234 4132
rect 18725 4123 18783 4129
rect 18725 4120 18737 4123
rect 18228 4092 18737 4120
rect 18228 4080 18234 4092
rect 18725 4089 18737 4092
rect 18771 4089 18783 4123
rect 18725 4083 18783 4089
rect 24794 4080 24800 4132
rect 24852 4120 24858 4132
rect 24889 4123 24947 4129
rect 24889 4120 24901 4123
rect 24852 4092 24901 4120
rect 24852 4080 24858 4092
rect 24889 4089 24901 4092
rect 24935 4089 24947 4123
rect 25162 4120 25168 4132
rect 25123 4092 25168 4120
rect 24889 4083 24947 4089
rect 4646 4012 4652 4064
rect 4704 4052 4710 4064
rect 5474 4052 5480 4064
rect 4704 4024 5480 4052
rect 4704 4012 4710 4024
rect 5474 4012 5480 4024
rect 5532 4052 5538 4064
rect 7501 4055 7559 4061
rect 5532 4024 5796 4052
rect 5532 4012 5538 4024
rect 3453 3987 3511 3993
rect 3453 3953 3465 3987
rect 3499 3984 3511 3987
rect 3910 3984 3916 3996
rect 3499 3956 3916 3984
rect 3499 3953 3511 3956
rect 3453 3947 3511 3953
rect 3910 3944 3916 3956
rect 3968 3944 3974 3996
rect 5569 3987 5627 3993
rect 5569 3953 5581 3987
rect 5615 3984 5627 3987
rect 5658 3984 5664 3996
rect 5615 3956 5664 3984
rect 5615 3953 5627 3956
rect 5569 3947 5627 3953
rect 5658 3944 5664 3956
rect 5716 3944 5722 3996
rect 5768 3993 5796 4024
rect 7501 4021 7513 4055
rect 7547 4052 7559 4055
rect 7590 4052 7596 4064
rect 7547 4024 7596 4052
rect 7547 4021 7559 4024
rect 7501 4015 7559 4021
rect 7590 4012 7596 4024
rect 7648 4012 7654 4064
rect 12285 4055 12343 4061
rect 12285 4052 12297 4055
rect 11656 4024 12297 4052
rect 5753 3987 5811 3993
rect 5753 3953 5765 3987
rect 5799 3953 5811 3987
rect 5934 3984 5940 3996
rect 5895 3956 5940 3984
rect 5753 3947 5811 3953
rect 5934 3944 5940 3956
rect 5992 3944 5998 3996
rect 6946 3984 6952 3996
rect 6907 3956 6952 3984
rect 6946 3944 6952 3956
rect 7004 3944 7010 3996
rect 7130 3984 7136 3996
rect 7091 3956 7136 3984
rect 7130 3944 7136 3956
rect 7188 3944 7194 3996
rect 11656 3993 11684 4024
rect 12285 4021 12297 4024
rect 12331 4052 12343 4055
rect 12374 4052 12380 4064
rect 12331 4024 12380 4052
rect 12331 4021 12343 4024
rect 12285 4015 12343 4021
rect 12374 4012 12380 4024
rect 12432 4012 12438 4064
rect 16790 4012 16796 4064
rect 16848 4052 16854 4064
rect 17253 4055 17311 4061
rect 17253 4052 17265 4055
rect 16848 4024 17265 4052
rect 16848 4012 16854 4024
rect 17253 4021 17265 4024
rect 17299 4021 17311 4055
rect 17253 4015 17311 4021
rect 17342 4012 17348 4064
rect 17400 4052 17406 4064
rect 17400 4024 18308 4052
rect 17400 4012 17406 4024
rect 10905 3987 10963 3993
rect 10905 3953 10917 3987
rect 10951 3984 10963 3987
rect 11641 3987 11699 3993
rect 11641 3984 11653 3987
rect 10951 3956 11653 3984
rect 10951 3953 10963 3956
rect 10905 3947 10963 3953
rect 11641 3953 11653 3956
rect 11687 3953 11699 3987
rect 12006 3984 12012 3996
rect 11967 3956 12012 3984
rect 11641 3947 11699 3953
rect 12006 3944 12012 3956
rect 12064 3944 12070 3996
rect 14585 3987 14643 3993
rect 14585 3953 14597 3987
rect 14631 3984 14643 3987
rect 14950 3984 14956 3996
rect 14631 3956 14956 3984
rect 14631 3953 14643 3956
rect 14585 3947 14643 3953
rect 14950 3944 14956 3956
rect 15008 3984 15014 3996
rect 15873 3987 15931 3993
rect 15873 3984 15885 3987
rect 15008 3956 15885 3984
rect 15008 3944 15014 3956
rect 15873 3953 15885 3956
rect 15919 3953 15931 3987
rect 17894 3984 17900 3996
rect 17855 3956 17900 3984
rect 15873 3947 15931 3953
rect 17894 3944 17900 3956
rect 17952 3944 17958 3996
rect 18280 3993 18308 4024
rect 18354 4012 18360 4064
rect 18412 4052 18418 4064
rect 18541 4055 18599 4061
rect 18541 4052 18553 4055
rect 18412 4024 18553 4052
rect 18412 4012 18418 4024
rect 18541 4021 18553 4024
rect 18587 4021 18599 4055
rect 24904 4052 24932 4083
rect 25162 4080 25168 4092
rect 25220 4080 25226 4132
rect 28014 4080 28020 4132
rect 28072 4120 28078 4132
rect 28201 4123 28259 4129
rect 28201 4120 28213 4123
rect 28072 4092 28213 4120
rect 28072 4080 28078 4092
rect 28201 4089 28213 4092
rect 28247 4089 28259 4123
rect 28201 4083 28259 4089
rect 24904 4024 25944 4052
rect 18541 4015 18599 4021
rect 18265 3987 18323 3993
rect 18265 3953 18277 3987
rect 18311 3953 18323 3987
rect 21666 3984 21672 3996
rect 21627 3956 21672 3984
rect 18265 3947 18323 3953
rect 21666 3944 21672 3956
rect 21724 3944 21730 3996
rect 21850 3944 21856 3996
rect 21908 3984 21914 3996
rect 22037 3987 22095 3993
rect 22037 3984 22049 3987
rect 21908 3956 22049 3984
rect 21908 3944 21914 3956
rect 22037 3953 22049 3956
rect 22083 3953 22095 3987
rect 22037 3947 22095 3953
rect 23693 3987 23751 3993
rect 23693 3953 23705 3987
rect 23739 3984 23751 3987
rect 23874 3984 23880 3996
rect 23739 3956 23880 3984
rect 23739 3953 23751 3956
rect 23693 3947 23751 3953
rect 23874 3944 23880 3956
rect 23932 3944 23938 3996
rect 24058 3984 24064 3996
rect 24019 3956 24064 3984
rect 24058 3944 24064 3956
rect 24116 3944 24122 3996
rect 25916 3993 25944 4024
rect 26174 4012 26180 4064
rect 26232 4052 26238 4064
rect 26361 4055 26419 4061
rect 26361 4052 26373 4055
rect 26232 4024 26373 4052
rect 26232 4012 26238 4024
rect 26361 4021 26373 4024
rect 26407 4021 26419 4055
rect 26361 4015 26419 4021
rect 24245 3987 24303 3993
rect 24245 3953 24257 3987
rect 24291 3984 24303 3987
rect 25809 3987 25867 3993
rect 25809 3984 25821 3987
rect 24291 3956 25821 3984
rect 24291 3953 24303 3956
rect 24245 3947 24303 3953
rect 25809 3953 25821 3956
rect 25855 3953 25867 3987
rect 25809 3947 25867 3953
rect 25901 3987 25959 3993
rect 25901 3953 25913 3987
rect 25947 3984 25959 3987
rect 26082 3984 26088 3996
rect 25947 3956 26088 3984
rect 25947 3953 25959 3956
rect 25901 3947 25959 3953
rect 3266 3876 3272 3928
rect 3324 3916 3330 3928
rect 3361 3919 3419 3925
rect 3361 3916 3373 3919
rect 3324 3888 3373 3916
rect 3324 3876 3330 3888
rect 3361 3885 3373 3888
rect 3407 3885 3419 3919
rect 11730 3916 11736 3928
rect 11691 3888 11736 3916
rect 3361 3879 3419 3885
rect 11730 3876 11736 3888
rect 11788 3876 11794 3928
rect 11917 3919 11975 3925
rect 11917 3885 11929 3919
rect 11963 3885 11975 3919
rect 11917 3879 11975 3885
rect 5382 3848 5388 3860
rect 5343 3820 5388 3848
rect 5382 3808 5388 3820
rect 5440 3808 5446 3860
rect 9154 3808 9160 3860
rect 9212 3848 9218 3860
rect 9433 3851 9491 3857
rect 9433 3848 9445 3851
rect 9212 3820 9445 3848
rect 9212 3808 9218 3820
rect 9433 3817 9445 3820
rect 9479 3848 9491 3851
rect 10166 3848 10172 3860
rect 9479 3820 10172 3848
rect 9479 3817 9491 3820
rect 9433 3811 9491 3817
rect 10166 3808 10172 3820
rect 10224 3808 10230 3860
rect 10626 3808 10632 3860
rect 10684 3848 10690 3860
rect 11638 3848 11644 3860
rect 10684 3820 11644 3848
rect 10684 3808 10690 3820
rect 11638 3808 11644 3820
rect 11696 3848 11702 3860
rect 11932 3848 11960 3879
rect 14398 3876 14404 3928
rect 14456 3916 14462 3928
rect 14769 3919 14827 3925
rect 14769 3916 14781 3919
rect 14456 3888 14781 3916
rect 14456 3876 14462 3888
rect 14769 3885 14781 3888
rect 14815 3916 14827 3919
rect 15413 3919 15471 3925
rect 15413 3916 15425 3919
rect 14815 3888 15425 3916
rect 14815 3885 14827 3888
rect 14769 3879 14827 3885
rect 15413 3885 15425 3888
rect 15459 3916 15471 3919
rect 15686 3916 15692 3928
rect 15459 3888 15692 3916
rect 15459 3885 15471 3888
rect 15413 3879 15471 3885
rect 15686 3876 15692 3888
rect 15744 3876 15750 3928
rect 17802 3916 17808 3928
rect 17763 3888 17808 3916
rect 17802 3876 17808 3888
rect 17860 3876 17866 3928
rect 18357 3919 18415 3925
rect 18357 3885 18369 3919
rect 18403 3885 18415 3919
rect 18357 3879 18415 3885
rect 11696 3820 11960 3848
rect 11696 3808 11702 3820
rect 14490 3808 14496 3860
rect 14548 3848 14554 3860
rect 15965 3851 16023 3857
rect 15965 3848 15977 3851
rect 14548 3820 15977 3848
rect 14548 3808 14554 3820
rect 15965 3817 15977 3820
rect 16011 3848 16023 3851
rect 16054 3848 16060 3860
rect 16011 3820 16060 3848
rect 16011 3817 16023 3820
rect 15965 3811 16023 3817
rect 16054 3808 16060 3820
rect 16112 3808 16118 3860
rect 17526 3808 17532 3860
rect 17584 3848 17590 3860
rect 18372 3848 18400 3879
rect 20470 3876 20476 3928
rect 20528 3916 20534 3928
rect 21482 3916 21488 3928
rect 20528 3888 21488 3916
rect 20528 3876 20534 3888
rect 21482 3876 21488 3888
rect 21540 3876 21546 3928
rect 21945 3919 22003 3925
rect 21945 3885 21957 3919
rect 21991 3916 22003 3919
rect 22218 3916 22224 3928
rect 21991 3888 22224 3916
rect 21991 3885 22003 3888
rect 21945 3879 22003 3885
rect 19182 3848 19188 3860
rect 17584 3820 19188 3848
rect 17584 3808 17590 3820
rect 19182 3808 19188 3820
rect 19240 3808 19246 3860
rect 21022 3808 21028 3860
rect 21080 3848 21086 3860
rect 21960 3848 21988 3879
rect 22218 3876 22224 3888
rect 22276 3876 22282 3928
rect 23782 3916 23788 3928
rect 23743 3888 23788 3916
rect 23782 3876 23788 3888
rect 23840 3876 23846 3928
rect 21080 3820 21988 3848
rect 21080 3808 21086 3820
rect 23138 3808 23144 3860
rect 23196 3848 23202 3860
rect 24260 3848 24288 3947
rect 26082 3944 26088 3956
rect 26140 3944 26146 3996
rect 28216 3984 28244 4083
rect 28658 4080 28664 4132
rect 28716 4120 28722 4132
rect 28716 4092 29164 4120
rect 28716 4080 28722 4092
rect 29136 4064 29164 4092
rect 29118 4012 29124 4064
rect 29176 4012 29182 4064
rect 28385 3987 28443 3993
rect 28385 3984 28397 3987
rect 28216 3956 28397 3984
rect 28385 3953 28397 3956
rect 28431 3953 28443 3987
rect 28385 3947 28443 3953
rect 28750 3916 28756 3928
rect 28711 3888 28756 3916
rect 28750 3876 28756 3888
rect 28808 3876 28814 3928
rect 23196 3820 24288 3848
rect 23196 3808 23202 3820
rect 2346 3780 2352 3792
rect 2259 3752 2352 3780
rect 2346 3740 2352 3752
rect 2404 3780 2410 3792
rect 2898 3780 2904 3792
rect 2404 3752 2904 3780
rect 2404 3740 2410 3752
rect 2898 3740 2904 3752
rect 2956 3740 2962 3792
rect 3358 3740 3364 3792
rect 3416 3780 3422 3792
rect 3637 3783 3695 3789
rect 3637 3780 3649 3783
rect 3416 3752 3649 3780
rect 3416 3740 3422 3752
rect 3637 3749 3649 3752
rect 3683 3749 3695 3783
rect 11270 3780 11276 3792
rect 11231 3752 11276 3780
rect 3637 3743 3695 3749
rect 11270 3740 11276 3752
rect 11328 3740 11334 3792
rect 18906 3780 18912 3792
rect 18867 3752 18912 3780
rect 18906 3740 18912 3752
rect 18964 3740 18970 3792
rect 21298 3780 21304 3792
rect 21259 3752 21304 3780
rect 21298 3740 21304 3752
rect 21356 3740 21362 3792
rect 23322 3780 23328 3792
rect 23283 3752 23328 3780
rect 23322 3740 23328 3752
rect 23380 3740 23386 3792
rect 30498 3780 30504 3792
rect 30459 3752 30504 3780
rect 30498 3740 30504 3752
rect 30556 3740 30562 3792
rect 400 3690 31680 3712
rect 400 3638 3510 3690
rect 3562 3638 3574 3690
rect 3626 3638 3638 3690
rect 3690 3638 3702 3690
rect 3754 3638 3766 3690
rect 3818 3638 31680 3690
rect 400 3616 31680 3638
rect 1242 3576 1248 3588
rect 1203 3548 1248 3576
rect 1242 3536 1248 3548
rect 1300 3536 1306 3588
rect 3637 3579 3695 3585
rect 3637 3545 3649 3579
rect 3683 3576 3695 3579
rect 3910 3576 3916 3588
rect 3683 3548 3916 3576
rect 3683 3545 3695 3548
rect 3637 3539 3695 3545
rect 3910 3536 3916 3548
rect 3968 3576 3974 3588
rect 4005 3579 4063 3585
rect 4005 3576 4017 3579
rect 3968 3548 4017 3576
rect 3968 3536 3974 3548
rect 4005 3545 4017 3548
rect 4051 3576 4063 3579
rect 4370 3576 4376 3588
rect 4051 3548 4376 3576
rect 4051 3545 4063 3548
rect 4005 3539 4063 3545
rect 4370 3536 4376 3548
rect 4428 3536 4434 3588
rect 5382 3576 5388 3588
rect 5343 3548 5388 3576
rect 5382 3536 5388 3548
rect 5440 3536 5446 3588
rect 5474 3536 5480 3588
rect 5532 3576 5538 3588
rect 5532 3548 5577 3576
rect 5532 3536 5538 3548
rect 5658 3536 5664 3588
rect 5716 3576 5722 3588
rect 6397 3579 6455 3585
rect 6397 3576 6409 3579
rect 5716 3548 6409 3576
rect 5716 3536 5722 3548
rect 6397 3545 6409 3548
rect 6443 3545 6455 3579
rect 6946 3576 6952 3588
rect 6907 3548 6952 3576
rect 6397 3539 6455 3545
rect 6946 3536 6952 3548
rect 7004 3536 7010 3588
rect 7130 3576 7136 3588
rect 7091 3548 7136 3576
rect 7130 3536 7136 3548
rect 7188 3536 7194 3588
rect 7409 3579 7467 3585
rect 7409 3545 7421 3579
rect 7455 3576 7467 3579
rect 7590 3576 7596 3588
rect 7455 3548 7596 3576
rect 7455 3545 7467 3548
rect 7409 3539 7467 3545
rect 7590 3536 7596 3548
rect 7648 3536 7654 3588
rect 11270 3576 11276 3588
rect 11231 3548 11276 3576
rect 11270 3536 11276 3548
rect 11328 3536 11334 3588
rect 14950 3536 14956 3588
rect 15008 3576 15014 3588
rect 15045 3579 15103 3585
rect 15045 3576 15057 3579
rect 15008 3548 15057 3576
rect 15008 3536 15014 3548
rect 15045 3545 15057 3548
rect 15091 3576 15103 3579
rect 15502 3576 15508 3588
rect 15091 3548 15508 3576
rect 15091 3545 15103 3548
rect 15045 3539 15103 3545
rect 15502 3536 15508 3548
rect 15560 3576 15566 3588
rect 15873 3579 15931 3585
rect 15873 3576 15885 3579
rect 15560 3548 15885 3576
rect 15560 3536 15566 3548
rect 15873 3545 15885 3548
rect 15919 3545 15931 3579
rect 16054 3576 16060 3588
rect 16015 3548 16060 3576
rect 15873 3539 15931 3545
rect 16054 3536 16060 3548
rect 16112 3536 16118 3588
rect 16790 3576 16796 3588
rect 16751 3548 16796 3576
rect 16790 3536 16796 3548
rect 16848 3536 16854 3588
rect 18173 3579 18231 3585
rect 18173 3545 18185 3579
rect 18219 3576 18231 3579
rect 18446 3576 18452 3588
rect 18219 3548 18452 3576
rect 18219 3545 18231 3548
rect 18173 3539 18231 3545
rect 18446 3536 18452 3548
rect 18504 3576 18510 3588
rect 18906 3576 18912 3588
rect 18504 3548 18912 3576
rect 18504 3536 18510 3548
rect 18906 3536 18912 3548
rect 18964 3536 18970 3588
rect 19829 3579 19887 3585
rect 19829 3545 19841 3579
rect 19875 3576 19887 3579
rect 20194 3576 20200 3588
rect 19875 3548 20200 3576
rect 19875 3545 19887 3548
rect 19829 3539 19887 3545
rect 20194 3536 20200 3548
rect 20252 3576 20258 3588
rect 20381 3579 20439 3585
rect 20381 3576 20393 3579
rect 20252 3548 20393 3576
rect 20252 3536 20258 3548
rect 20381 3545 20393 3548
rect 20427 3545 20439 3579
rect 21022 3576 21028 3588
rect 20983 3548 21028 3576
rect 20381 3539 20439 3545
rect 21022 3536 21028 3548
rect 21080 3536 21086 3588
rect 21298 3576 21304 3588
rect 21259 3548 21304 3576
rect 21298 3536 21304 3548
rect 21356 3536 21362 3588
rect 21669 3579 21727 3585
rect 21669 3545 21681 3579
rect 21715 3576 21727 3579
rect 21850 3576 21856 3588
rect 21715 3548 21856 3576
rect 21715 3545 21727 3548
rect 21669 3539 21727 3545
rect 21850 3536 21856 3548
rect 21908 3536 21914 3588
rect 23322 3576 23328 3588
rect 23283 3548 23328 3576
rect 23322 3536 23328 3548
rect 23380 3536 23386 3588
rect 27649 3579 27707 3585
rect 27649 3545 27661 3579
rect 27695 3576 27707 3579
rect 27833 3579 27891 3585
rect 27833 3576 27845 3579
rect 27695 3548 27845 3576
rect 27695 3545 27707 3548
rect 27649 3539 27707 3545
rect 27833 3545 27845 3548
rect 27879 3576 27891 3579
rect 28750 3576 28756 3588
rect 27879 3548 28756 3576
rect 27879 3545 27891 3548
rect 27833 3539 27891 3545
rect 28750 3536 28756 3548
rect 28808 3576 28814 3588
rect 28845 3579 28903 3585
rect 28845 3576 28857 3579
rect 28808 3548 28857 3576
rect 28808 3536 28814 3548
rect 28845 3545 28857 3548
rect 28891 3545 28903 3579
rect 28845 3539 28903 3545
rect 5201 3511 5259 3517
rect 5201 3477 5213 3511
rect 5247 3508 5259 3511
rect 5934 3508 5940 3520
rect 5247 3480 5940 3508
rect 5247 3477 5259 3480
rect 5201 3471 5259 3477
rect 5934 3468 5940 3480
rect 5992 3468 5998 3520
rect 3358 3440 3364 3452
rect 2732 3412 3364 3440
rect 2732 3381 2760 3412
rect 3358 3400 3364 3412
rect 3416 3400 3422 3452
rect 4189 3443 4247 3449
rect 4189 3409 4201 3443
rect 4235 3440 4247 3443
rect 4925 3443 4983 3449
rect 4925 3440 4937 3443
rect 4235 3412 4937 3440
rect 4235 3409 4247 3412
rect 4189 3403 4247 3409
rect 4925 3409 4937 3412
rect 4971 3440 4983 3443
rect 5842 3440 5848 3452
rect 4971 3412 5848 3440
rect 4971 3409 4983 3412
rect 4925 3403 4983 3409
rect 2717 3375 2775 3381
rect 2717 3341 2729 3375
rect 2763 3341 2775 3375
rect 2898 3372 2904 3384
rect 2859 3344 2904 3372
rect 2717 3335 2775 3341
rect 2898 3332 2904 3344
rect 2956 3332 2962 3384
rect 3085 3375 3143 3381
rect 3085 3341 3097 3375
rect 3131 3372 3143 3375
rect 4204 3372 4232 3403
rect 5842 3400 5848 3412
rect 5900 3440 5906 3452
rect 6964 3440 6992 3536
rect 10721 3511 10779 3517
rect 10721 3477 10733 3511
rect 10767 3508 10779 3511
rect 12006 3508 12012 3520
rect 10767 3480 12012 3508
rect 10767 3477 10779 3480
rect 10721 3471 10779 3477
rect 12006 3468 12012 3480
rect 12064 3468 12070 3520
rect 12374 3468 12380 3520
rect 12432 3508 12438 3520
rect 13110 3508 13116 3520
rect 12432 3480 13116 3508
rect 12432 3468 12438 3480
rect 13110 3468 13116 3480
rect 13168 3508 13174 3520
rect 13205 3511 13263 3517
rect 13205 3508 13217 3511
rect 13168 3480 13217 3508
rect 13168 3468 13174 3480
rect 13205 3477 13217 3480
rect 13251 3477 13263 3511
rect 13205 3471 13263 3477
rect 5900 3412 6992 3440
rect 8881 3443 8939 3449
rect 5900 3400 5906 3412
rect 8881 3409 8893 3443
rect 8927 3440 8939 3443
rect 9890 3440 9896 3452
rect 8927 3412 9896 3440
rect 8927 3409 8939 3412
rect 8881 3403 8939 3409
rect 9890 3400 9896 3412
rect 9948 3440 9954 3452
rect 10077 3443 10135 3449
rect 9948 3412 10028 3440
rect 9948 3400 9954 3412
rect 4370 3381 4376 3384
rect 3131 3344 4232 3372
rect 4322 3375 4376 3381
rect 3131 3341 3143 3344
rect 3085 3335 3143 3341
rect 4322 3341 4334 3375
rect 4368 3341 4376 3375
rect 4322 3335 4376 3341
rect 1058 3264 1064 3316
rect 1116 3304 1122 3316
rect 1981 3307 2039 3313
rect 1981 3304 1993 3307
rect 1116 3276 1993 3304
rect 1116 3264 1122 3276
rect 1981 3273 1993 3276
rect 2027 3304 2039 3307
rect 2257 3307 2315 3313
rect 2257 3304 2269 3307
rect 2027 3276 2269 3304
rect 2027 3273 2039 3276
rect 1981 3267 2039 3273
rect 2257 3273 2269 3276
rect 2303 3273 2315 3307
rect 2257 3267 2315 3273
rect 2165 3239 2223 3245
rect 2165 3205 2177 3239
rect 2211 3236 2223 3239
rect 3100 3236 3128 3335
rect 4370 3332 4376 3335
rect 4428 3372 4434 3384
rect 5937 3375 5995 3381
rect 5937 3372 5949 3375
rect 4428 3344 5949 3372
rect 4428 3332 4434 3344
rect 5937 3341 5949 3344
rect 5983 3341 5995 3375
rect 5937 3335 5995 3341
rect 4741 3307 4799 3313
rect 4741 3304 4753 3307
rect 4526 3276 4753 3304
rect 2211 3208 3128 3236
rect 2211 3205 2223 3208
rect 2165 3199 2223 3205
rect 3266 3196 3272 3248
rect 3324 3236 3330 3248
rect 3361 3239 3419 3245
rect 3361 3236 3373 3239
rect 3324 3208 3373 3236
rect 3324 3196 3330 3208
rect 3361 3205 3373 3208
rect 3407 3205 3419 3239
rect 3910 3236 3916 3248
rect 3871 3208 3916 3236
rect 3361 3199 3419 3205
rect 3910 3196 3916 3208
rect 3968 3236 3974 3248
rect 4526 3236 4554 3276
rect 4741 3273 4753 3276
rect 4787 3273 4799 3307
rect 5952 3304 5980 3335
rect 6026 3332 6032 3384
rect 6084 3372 6090 3384
rect 10000 3381 10028 3412
rect 10077 3409 10089 3443
rect 10123 3440 10135 3443
rect 10166 3440 10172 3452
rect 10123 3412 10172 3440
rect 10123 3409 10135 3412
rect 10077 3403 10135 3409
rect 10166 3400 10172 3412
rect 10224 3400 10230 3452
rect 10905 3443 10963 3449
rect 10905 3409 10917 3443
rect 10951 3440 10963 3443
rect 11730 3440 11736 3452
rect 10951 3412 11736 3440
rect 10951 3409 10963 3412
rect 10905 3403 10963 3409
rect 11730 3400 11736 3412
rect 11788 3400 11794 3452
rect 12024 3440 12052 3468
rect 13220 3440 13248 3471
rect 13846 3468 13852 3520
rect 13904 3508 13910 3520
rect 13904 3480 14444 3508
rect 13904 3468 13910 3480
rect 14416 3440 14444 3480
rect 15410 3468 15416 3520
rect 15468 3508 15474 3520
rect 17069 3511 17127 3517
rect 17069 3508 17081 3511
rect 15468 3480 17081 3508
rect 15468 3468 15474 3480
rect 17069 3477 17081 3480
rect 17115 3508 17127 3511
rect 17802 3508 17808 3520
rect 17115 3480 17808 3508
rect 17115 3477 17127 3480
rect 17069 3471 17127 3477
rect 17802 3468 17808 3480
rect 17860 3468 17866 3520
rect 17989 3511 18047 3517
rect 17989 3477 18001 3511
rect 18035 3508 18047 3511
rect 18035 3480 18952 3508
rect 18035 3477 18047 3480
rect 17989 3471 18047 3477
rect 14493 3443 14551 3449
rect 14493 3440 14505 3443
rect 12024 3412 12788 3440
rect 13220 3412 14260 3440
rect 14416 3412 14505 3440
rect 6121 3375 6179 3381
rect 6121 3372 6133 3375
rect 6084 3344 6133 3372
rect 6084 3332 6090 3344
rect 6121 3341 6133 3344
rect 6167 3341 6179 3375
rect 6121 3335 6179 3341
rect 6213 3375 6271 3381
rect 6213 3341 6225 3375
rect 6259 3341 6271 3375
rect 6213 3335 6271 3341
rect 9985 3375 10043 3381
rect 9985 3341 9997 3375
rect 10031 3341 10043 3375
rect 10350 3372 10356 3384
rect 10311 3344 10356 3372
rect 9985 3335 10043 3341
rect 6228 3304 6256 3335
rect 10350 3332 10356 3344
rect 10408 3332 10414 3384
rect 10445 3375 10503 3381
rect 10445 3341 10457 3375
rect 10491 3372 10503 3375
rect 10534 3372 10540 3384
rect 10491 3344 10540 3372
rect 10491 3341 10503 3344
rect 10445 3335 10503 3341
rect 5952 3276 6256 3304
rect 4741 3267 4799 3273
rect 8142 3264 8148 3316
rect 8200 3304 8206 3316
rect 9065 3307 9123 3313
rect 9065 3304 9077 3307
rect 8200 3276 9077 3304
rect 8200 3264 8206 3276
rect 9065 3273 9077 3276
rect 9111 3304 9123 3307
rect 9341 3307 9399 3313
rect 9341 3304 9353 3307
rect 9111 3276 9353 3304
rect 9111 3273 9123 3276
rect 9065 3267 9123 3273
rect 9341 3273 9353 3276
rect 9387 3273 9399 3307
rect 9341 3267 9399 3273
rect 5658 3236 5664 3248
rect 3968 3208 4554 3236
rect 5619 3208 5664 3236
rect 3968 3196 3974 3208
rect 5658 3196 5664 3208
rect 5716 3196 5722 3248
rect 6026 3196 6032 3248
rect 6084 3236 6090 3248
rect 6765 3239 6823 3245
rect 6765 3236 6777 3239
rect 6084 3208 6777 3236
rect 6084 3196 6090 3208
rect 6765 3205 6777 3208
rect 6811 3236 6823 3239
rect 7498 3236 7504 3248
rect 6811 3208 7504 3236
rect 6811 3205 6823 3208
rect 6765 3199 6823 3205
rect 7498 3196 7504 3208
rect 7556 3196 7562 3248
rect 9246 3236 9252 3248
rect 9207 3208 9252 3236
rect 9246 3196 9252 3208
rect 9304 3236 9310 3248
rect 10460 3236 10488 3335
rect 10534 3332 10540 3344
rect 10592 3332 10598 3384
rect 12098 3332 12104 3384
rect 12156 3372 12162 3384
rect 12193 3375 12251 3381
rect 12193 3372 12205 3375
rect 12156 3344 12205 3372
rect 12156 3332 12162 3344
rect 12193 3341 12205 3344
rect 12239 3372 12251 3375
rect 12282 3372 12288 3384
rect 12239 3344 12288 3372
rect 12239 3341 12251 3344
rect 12193 3335 12251 3341
rect 12282 3332 12288 3344
rect 12340 3332 12346 3384
rect 12374 3332 12380 3384
rect 12432 3372 12438 3384
rect 12760 3381 12788 3412
rect 12745 3375 12803 3381
rect 12432 3344 12477 3372
rect 12432 3332 12438 3344
rect 12745 3341 12757 3375
rect 12791 3341 12803 3375
rect 12926 3372 12932 3384
rect 12887 3344 12932 3372
rect 12745 3335 12803 3341
rect 12926 3332 12932 3344
rect 12984 3332 12990 3384
rect 11549 3307 11607 3313
rect 11549 3273 11561 3307
rect 11595 3304 11607 3307
rect 11730 3304 11736 3316
rect 11595 3276 11736 3304
rect 11595 3273 11607 3276
rect 11549 3267 11607 3273
rect 11730 3264 11736 3276
rect 11788 3304 11794 3316
rect 12944 3304 12972 3332
rect 13478 3304 13484 3316
rect 11788 3276 12972 3304
rect 13391 3276 13484 3304
rect 11788 3264 11794 3276
rect 13478 3264 13484 3276
rect 13536 3304 13542 3316
rect 13757 3307 13815 3313
rect 13757 3304 13769 3307
rect 13536 3276 13769 3304
rect 13536 3264 13542 3276
rect 13757 3273 13769 3276
rect 13803 3273 13815 3307
rect 14232 3304 14260 3412
rect 14493 3409 14505 3412
rect 14539 3409 14551 3443
rect 15229 3443 15287 3449
rect 15229 3440 15241 3443
rect 14493 3403 14551 3409
rect 14600 3412 15241 3440
rect 14398 3332 14404 3384
rect 14456 3372 14462 3384
rect 14600 3372 14628 3412
rect 15229 3409 15241 3412
rect 15275 3409 15287 3443
rect 17820 3440 17848 3468
rect 18630 3440 18636 3452
rect 17820 3412 18636 3440
rect 15229 3403 15287 3409
rect 18630 3400 18636 3412
rect 18688 3400 18694 3452
rect 14766 3372 14772 3384
rect 14456 3344 14628 3372
rect 14727 3344 14772 3372
rect 14456 3332 14462 3344
rect 14766 3332 14772 3344
rect 14824 3332 14830 3384
rect 14953 3375 15011 3381
rect 14953 3341 14965 3375
rect 14999 3372 15011 3375
rect 15686 3372 15692 3384
rect 14999 3344 15692 3372
rect 14999 3341 15011 3344
rect 14953 3335 15011 3341
rect 14416 3304 14444 3332
rect 14232 3276 14444 3304
rect 13757 3267 13815 3273
rect 9304 3208 10488 3236
rect 11089 3239 11147 3245
rect 9304 3196 9310 3208
rect 11089 3205 11101 3239
rect 11135 3236 11147 3239
rect 11638 3236 11644 3248
rect 11135 3208 11644 3236
rect 11135 3205 11147 3208
rect 11089 3199 11147 3205
rect 11638 3196 11644 3208
rect 11696 3196 11702 3248
rect 11822 3236 11828 3248
rect 11783 3208 11828 3236
rect 11822 3196 11828 3208
rect 11880 3196 11886 3248
rect 13570 3236 13576 3248
rect 13531 3208 13576 3236
rect 13570 3196 13576 3208
rect 13628 3236 13634 3248
rect 14968 3236 14996 3335
rect 15686 3332 15692 3344
rect 15744 3332 15750 3384
rect 16974 3372 16980 3384
rect 16887 3344 16980 3372
rect 16974 3332 16980 3344
rect 17032 3372 17038 3384
rect 17894 3372 17900 3384
rect 17032 3344 17900 3372
rect 17032 3332 17038 3344
rect 17894 3332 17900 3344
rect 17952 3332 17958 3384
rect 18747 3375 18805 3381
rect 18747 3372 18759 3375
rect 18648 3344 18759 3372
rect 18648 3316 18676 3344
rect 18747 3341 18759 3344
rect 18793 3341 18805 3375
rect 18924 3372 18952 3480
rect 21206 3468 21212 3520
rect 21264 3508 21270 3520
rect 24429 3511 24487 3517
rect 24429 3508 24441 3511
rect 21264 3480 24441 3508
rect 21264 3468 21270 3480
rect 24429 3477 24441 3480
rect 24475 3508 24487 3511
rect 24886 3508 24892 3520
rect 24475 3480 24892 3508
rect 24475 3477 24487 3480
rect 24429 3471 24487 3477
rect 24886 3468 24892 3480
rect 24944 3468 24950 3520
rect 25162 3468 25168 3520
rect 25220 3508 25226 3520
rect 25257 3511 25315 3517
rect 25257 3508 25269 3511
rect 25220 3480 25269 3508
rect 25220 3468 25226 3480
rect 25257 3477 25269 3480
rect 25303 3477 25315 3511
rect 25257 3471 25315 3477
rect 27278 3468 27284 3520
rect 27336 3508 27342 3520
rect 29210 3508 29216 3520
rect 27336 3480 29216 3508
rect 27336 3468 27342 3480
rect 29210 3468 29216 3480
rect 29268 3508 29274 3520
rect 30225 3511 30283 3517
rect 30225 3508 30237 3511
rect 29268 3480 30237 3508
rect 29268 3468 29274 3480
rect 30225 3477 30237 3480
rect 30271 3477 30283 3511
rect 30225 3471 30283 3477
rect 19182 3440 19188 3452
rect 19143 3412 19188 3440
rect 19182 3400 19188 3412
rect 19240 3440 19246 3452
rect 19921 3443 19979 3449
rect 19921 3440 19933 3443
rect 19240 3412 19933 3440
rect 19240 3400 19246 3412
rect 19921 3409 19933 3412
rect 19967 3440 19979 3443
rect 21482 3440 21488 3452
rect 19967 3412 20240 3440
rect 21443 3412 21488 3440
rect 19967 3409 19979 3412
rect 19921 3403 19979 3409
rect 19093 3375 19151 3381
rect 19093 3372 19105 3375
rect 18924 3344 19105 3372
rect 18747 3335 18805 3341
rect 19093 3341 19105 3344
rect 19139 3372 19151 3375
rect 19274 3372 19280 3384
rect 19139 3344 19280 3372
rect 19139 3341 19151 3344
rect 19093 3335 19151 3341
rect 19274 3332 19280 3344
rect 19332 3332 19338 3384
rect 20212 3381 20240 3412
rect 21482 3400 21488 3412
rect 21540 3400 21546 3452
rect 21850 3400 21856 3452
rect 21908 3440 21914 3452
rect 23601 3443 23659 3449
rect 23601 3440 23613 3443
rect 21908 3412 23613 3440
rect 21908 3400 21914 3412
rect 23601 3409 23613 3412
rect 23647 3409 23659 3443
rect 23601 3403 23659 3409
rect 20105 3375 20163 3381
rect 20105 3341 20117 3375
rect 20151 3341 20163 3375
rect 20105 3335 20163 3341
rect 20197 3375 20255 3381
rect 20197 3341 20209 3375
rect 20243 3341 20255 3375
rect 23616 3372 23644 3403
rect 23782 3400 23788 3452
rect 23840 3440 23846 3452
rect 29029 3443 29087 3449
rect 29029 3440 29041 3443
rect 23840 3412 29041 3440
rect 23840 3400 23846 3412
rect 29029 3409 29041 3412
rect 29075 3440 29087 3443
rect 29857 3443 29915 3449
rect 29857 3440 29869 3443
rect 29075 3412 29869 3440
rect 29075 3409 29087 3412
rect 29029 3403 29087 3409
rect 29857 3409 29869 3412
rect 29903 3409 29915 3443
rect 29857 3403 29915 3409
rect 24058 3372 24064 3384
rect 23616 3344 24064 3372
rect 20197 3335 20255 3341
rect 15042 3264 15048 3316
rect 15100 3304 15106 3316
rect 15100 3276 18032 3304
rect 15100 3264 15106 3276
rect 17342 3236 17348 3248
rect 13628 3208 14996 3236
rect 17303 3208 17348 3236
rect 13628 3196 13634 3208
rect 17342 3196 17348 3208
rect 17400 3196 17406 3248
rect 17526 3236 17532 3248
rect 17487 3208 17532 3236
rect 17526 3196 17532 3208
rect 17584 3236 17590 3248
rect 17713 3239 17771 3245
rect 17713 3236 17725 3239
rect 17584 3208 17725 3236
rect 17584 3196 17590 3208
rect 17713 3205 17725 3208
rect 17759 3205 17771 3239
rect 18004 3236 18032 3276
rect 18630 3264 18636 3316
rect 18688 3304 18694 3316
rect 19369 3307 19427 3313
rect 19369 3304 19381 3307
rect 18688 3276 19381 3304
rect 18688 3264 18694 3276
rect 19369 3273 19381 3276
rect 19415 3273 19427 3307
rect 19369 3267 19427 3273
rect 20120 3304 20148 3335
rect 24058 3332 24064 3344
rect 24116 3332 24122 3384
rect 24613 3375 24671 3381
rect 24613 3341 24625 3375
rect 24659 3372 24671 3375
rect 25530 3372 25536 3384
rect 24659 3344 25536 3372
rect 24659 3341 24671 3344
rect 24613 3335 24671 3341
rect 25530 3332 25536 3344
rect 25588 3332 25594 3384
rect 25625 3375 25683 3381
rect 25625 3341 25637 3375
rect 25671 3341 25683 3375
rect 26082 3372 26088 3384
rect 26043 3344 26088 3372
rect 25625 3335 25683 3341
rect 20749 3307 20807 3313
rect 20749 3304 20761 3307
rect 20120 3276 20761 3304
rect 20120 3236 20148 3276
rect 20749 3273 20761 3276
rect 20795 3273 20807 3307
rect 20749 3267 20807 3273
rect 21666 3264 21672 3316
rect 21724 3304 21730 3316
rect 21853 3307 21911 3313
rect 21853 3304 21865 3307
rect 21724 3276 21865 3304
rect 21724 3264 21730 3276
rect 21853 3273 21865 3276
rect 21899 3304 21911 3307
rect 21899 3276 23874 3304
rect 21899 3273 21911 3276
rect 21853 3267 21911 3273
rect 23846 3248 23874 3276
rect 23138 3236 23144 3248
rect 18004 3208 20148 3236
rect 23099 3208 23144 3236
rect 17713 3199 17771 3205
rect 23138 3196 23144 3208
rect 23196 3196 23202 3248
rect 23414 3236 23420 3248
rect 23375 3208 23420 3236
rect 23414 3196 23420 3208
rect 23472 3196 23478 3248
rect 23846 3208 23880 3248
rect 23874 3196 23880 3208
rect 23932 3236 23938 3248
rect 24794 3236 24800 3248
rect 23932 3208 23977 3236
rect 24707 3208 24800 3236
rect 23932 3196 23938 3208
rect 24794 3196 24800 3208
rect 24852 3236 24858 3248
rect 25640 3236 25668 3335
rect 26082 3332 26088 3344
rect 26140 3332 26146 3384
rect 26542 3372 26548 3384
rect 26503 3344 26548 3372
rect 26542 3332 26548 3344
rect 26600 3332 26606 3384
rect 28290 3332 28296 3384
rect 28348 3332 28354 3384
rect 29210 3372 29216 3384
rect 29171 3344 29216 3372
rect 29210 3332 29216 3344
rect 29268 3332 29274 3384
rect 29302 3332 29308 3384
rect 29360 3372 29366 3384
rect 29578 3372 29584 3384
rect 29360 3344 29584 3372
rect 29360 3332 29366 3344
rect 29578 3332 29584 3344
rect 29636 3332 29642 3384
rect 29765 3375 29823 3381
rect 29765 3341 29777 3375
rect 29811 3372 29823 3375
rect 30498 3372 30504 3384
rect 29811 3344 30504 3372
rect 29811 3341 29823 3344
rect 29765 3335 29823 3341
rect 28017 3307 28075 3313
rect 28017 3273 28029 3307
rect 28063 3304 28075 3307
rect 28201 3307 28259 3313
rect 28201 3304 28213 3307
rect 28063 3276 28213 3304
rect 28063 3273 28075 3276
rect 28017 3267 28075 3273
rect 28201 3273 28213 3276
rect 28247 3304 28259 3307
rect 28308 3304 28336 3332
rect 29780 3304 29808 3335
rect 30498 3332 30504 3344
rect 30556 3332 30562 3384
rect 28247 3276 29808 3304
rect 28247 3273 28259 3276
rect 28201 3267 28259 3273
rect 28290 3236 28296 3248
rect 24852 3208 25668 3236
rect 28251 3208 28296 3236
rect 24852 3196 24858 3208
rect 28290 3196 28296 3208
rect 28348 3236 28354 3248
rect 28750 3236 28756 3248
rect 28348 3208 28756 3236
rect 28348 3196 28354 3208
rect 28750 3196 28756 3208
rect 28808 3196 28814 3248
rect 29578 3196 29584 3248
rect 29636 3236 29642 3248
rect 30041 3239 30099 3245
rect 30041 3236 30053 3239
rect 29636 3208 30053 3236
rect 29636 3196 29642 3208
rect 30041 3205 30053 3208
rect 30087 3205 30099 3239
rect 30041 3199 30099 3205
rect 400 3146 31680 3168
rect 400 3094 18870 3146
rect 18922 3094 18934 3146
rect 18986 3094 18998 3146
rect 19050 3094 19062 3146
rect 19114 3094 19126 3146
rect 19178 3094 31680 3146
rect 400 3072 31680 3094
rect 1058 3032 1064 3044
rect 1019 3004 1064 3032
rect 1058 2992 1064 3004
rect 1116 2992 1122 3044
rect 2349 3035 2407 3041
rect 2349 3001 2361 3035
rect 2395 3032 2407 3035
rect 3358 3032 3364 3044
rect 2395 3004 3364 3032
rect 2395 3001 2407 3004
rect 2349 2995 2407 3001
rect 3358 2992 3364 3004
rect 3416 2992 3422 3044
rect 5201 3035 5259 3041
rect 5201 3001 5213 3035
rect 5247 3032 5259 3035
rect 5658 3032 5664 3044
rect 5247 3004 5664 3032
rect 5247 3001 5259 3004
rect 5201 2995 5259 3001
rect 5658 2992 5664 3004
rect 5716 2992 5722 3044
rect 8142 3032 8148 3044
rect 8103 3004 8148 3032
rect 8142 2992 8148 3004
rect 8200 2992 8206 3044
rect 9433 3035 9491 3041
rect 9433 3001 9445 3035
rect 9479 3032 9491 3035
rect 10350 3032 10356 3044
rect 9479 3004 10356 3032
rect 9479 3001 9491 3004
rect 9433 2995 9491 3001
rect 10350 2992 10356 3004
rect 10408 2992 10414 3044
rect 11822 3032 11828 3044
rect 11783 3004 11828 3032
rect 11822 2992 11828 3004
rect 11880 2992 11886 3044
rect 12006 2992 12012 3044
rect 12064 3032 12070 3044
rect 12193 3035 12251 3041
rect 12193 3032 12205 3035
rect 12064 3004 12205 3032
rect 12064 2992 12070 3004
rect 12193 3001 12205 3004
rect 12239 3032 12251 3035
rect 13386 3032 13392 3044
rect 12239 3004 13392 3032
rect 12239 3001 12251 3004
rect 12193 2995 12251 3001
rect 13386 2992 13392 3004
rect 13444 3032 13450 3044
rect 13757 3035 13815 3041
rect 13757 3032 13769 3035
rect 13444 3004 13769 3032
rect 13444 2992 13450 3004
rect 13757 3001 13769 3004
rect 13803 3032 13815 3035
rect 14766 3032 14772 3044
rect 13803 3004 14772 3032
rect 13803 3001 13815 3004
rect 13757 2995 13815 3001
rect 14766 2992 14772 3004
rect 14824 2992 14830 3044
rect 17802 2992 17808 3044
rect 17860 3032 17866 3044
rect 18081 3035 18139 3041
rect 18081 3032 18093 3035
rect 17860 3004 18093 3032
rect 17860 2992 17866 3004
rect 18081 3001 18093 3004
rect 18127 3001 18139 3035
rect 18081 2995 18139 3001
rect 18170 2992 18176 3044
rect 18228 3032 18234 3044
rect 18265 3035 18323 3041
rect 18265 3032 18277 3035
rect 18228 3004 18277 3032
rect 18228 2992 18234 3004
rect 18265 3001 18277 3004
rect 18311 3032 18323 3035
rect 18311 3004 18676 3032
rect 18311 3001 18323 3004
rect 18265 2995 18323 3001
rect 5382 2924 5388 2976
rect 5440 2964 5446 2976
rect 5753 2967 5811 2973
rect 5753 2964 5765 2967
rect 5440 2936 5765 2964
rect 5440 2924 5446 2936
rect 5753 2933 5765 2936
rect 5799 2933 5811 2967
rect 7498 2964 7504 2976
rect 7459 2936 7504 2964
rect 5753 2927 5811 2933
rect 7498 2924 7504 2936
rect 7556 2924 7562 2976
rect 11730 2964 11736 2976
rect 11691 2936 11736 2964
rect 11730 2924 11736 2936
rect 11788 2924 11794 2976
rect 12098 2964 12104 2976
rect 12059 2936 12104 2964
rect 12098 2924 12104 2936
rect 12156 2924 12162 2976
rect 13110 2964 13116 2976
rect 13071 2936 13116 2964
rect 13110 2924 13116 2936
rect 13168 2924 13174 2976
rect 15502 2964 15508 2976
rect 15463 2936 15508 2964
rect 15502 2924 15508 2936
rect 15560 2924 15566 2976
rect 17066 2964 17072 2976
rect 17027 2936 17072 2964
rect 17066 2924 17072 2936
rect 17124 2924 17130 2976
rect 17621 2967 17679 2973
rect 17621 2933 17633 2967
rect 17667 2964 17679 2967
rect 17894 2964 17900 2976
rect 17667 2936 17900 2964
rect 17667 2933 17679 2936
rect 17621 2927 17679 2933
rect 17894 2924 17900 2936
rect 17952 2924 17958 2976
rect 18648 2973 18676 3004
rect 21206 2992 21212 3044
rect 21264 3032 21270 3044
rect 21574 3032 21580 3044
rect 21264 3004 21580 3032
rect 21264 2992 21270 3004
rect 21574 2992 21580 3004
rect 21632 3032 21638 3044
rect 21632 3004 21896 3032
rect 21632 2992 21638 3004
rect 18633 2967 18691 2973
rect 18633 2933 18645 2967
rect 18679 2933 18691 2967
rect 18633 2927 18691 2933
rect 21298 2924 21304 2976
rect 21356 2964 21362 2976
rect 21393 2967 21451 2973
rect 21393 2964 21405 2967
rect 21356 2936 21405 2964
rect 21356 2924 21362 2936
rect 21393 2933 21405 2936
rect 21439 2933 21451 2967
rect 21868 2936 21896 3004
rect 22218 2992 22224 3044
rect 22276 3032 22282 3044
rect 22276 3004 23184 3032
rect 22276 2992 22282 3004
rect 23156 2973 23184 3004
rect 23322 2992 23328 3044
rect 23380 3032 23386 3044
rect 23509 3035 23567 3041
rect 23509 3032 23521 3035
rect 23380 3004 23521 3032
rect 23380 2992 23386 3004
rect 23509 3001 23521 3004
rect 23555 3001 23567 3035
rect 26174 3032 26180 3044
rect 26135 3004 26180 3032
rect 23509 2995 23567 3001
rect 26174 2992 26180 3004
rect 26232 2992 26238 3044
rect 23141 2967 23199 2973
rect 21393 2927 21451 2933
rect 23141 2933 23153 2967
rect 23187 2933 23199 2967
rect 26082 2964 26088 2976
rect 26043 2936 26088 2964
rect 23141 2927 23199 2933
rect 26082 2924 26088 2936
rect 26140 2924 26146 2976
rect 28750 2924 28756 2976
rect 28808 2924 28814 2976
rect 3358 2856 3364 2908
rect 3416 2896 3422 2908
rect 3910 2896 3916 2908
rect 3416 2868 3916 2896
rect 3416 2856 3422 2868
rect 3910 2856 3916 2868
rect 3968 2896 3974 2908
rect 4097 2899 4155 2905
rect 4097 2896 4109 2899
rect 3968 2868 4109 2896
rect 3968 2856 3974 2868
rect 4097 2865 4109 2868
rect 4143 2865 4155 2899
rect 4462 2896 4468 2908
rect 4423 2868 4468 2896
rect 4097 2859 4155 2865
rect 4462 2856 4468 2868
rect 4520 2856 4526 2908
rect 4557 2899 4615 2905
rect 4557 2865 4569 2899
rect 4603 2896 4615 2899
rect 4646 2896 4652 2908
rect 4603 2868 4652 2896
rect 4603 2865 4615 2868
rect 4557 2859 4615 2865
rect 4646 2856 4652 2868
rect 4704 2856 4710 2908
rect 6854 2856 6860 2908
rect 6912 2856 6918 2908
rect 11086 2856 11092 2908
rect 11144 2856 11150 2908
rect 11638 2856 11644 2908
rect 11696 2896 11702 2908
rect 13297 2899 13355 2905
rect 13297 2896 13309 2899
rect 11696 2868 13309 2896
rect 11696 2856 11702 2868
rect 13297 2865 13309 2868
rect 13343 2865 13355 2899
rect 15686 2896 15692 2908
rect 15647 2868 15692 2896
rect 13297 2859 13355 2865
rect 15686 2856 15692 2868
rect 15744 2856 15750 2908
rect 16238 2856 16244 2908
rect 16296 2896 16302 2908
rect 16882 2896 16888 2908
rect 16296 2868 16888 2896
rect 16296 2856 16302 2868
rect 16882 2856 16888 2868
rect 16940 2856 16946 2908
rect 17158 2896 17164 2908
rect 17119 2868 17164 2896
rect 17158 2856 17164 2868
rect 17216 2856 17222 2908
rect 18725 2899 18783 2905
rect 18725 2865 18737 2899
rect 18771 2865 18783 2899
rect 21114 2896 21120 2908
rect 21075 2868 21120 2896
rect 18725 2859 18783 2865
rect 4002 2788 4008 2840
rect 4060 2828 4066 2840
rect 5477 2831 5535 2837
rect 4060 2800 4554 2828
rect 4060 2788 4066 2800
rect 3910 2760 3916 2772
rect 3871 2732 3916 2760
rect 3910 2720 3916 2732
rect 3968 2720 3974 2772
rect 4526 2760 4554 2800
rect 5477 2797 5489 2831
rect 5523 2828 5535 2831
rect 6118 2828 6124 2840
rect 5523 2800 6124 2828
rect 5523 2797 5535 2800
rect 5477 2791 5535 2797
rect 5492 2760 5520 2791
rect 6118 2788 6124 2800
rect 6176 2788 6182 2840
rect 9706 2828 9712 2840
rect 9667 2800 9712 2828
rect 9706 2788 9712 2800
rect 9764 2788 9770 2840
rect 9982 2828 9988 2840
rect 9943 2800 9988 2828
rect 9982 2788 9988 2800
rect 10040 2788 10046 2840
rect 16054 2828 16060 2840
rect 16015 2800 16060 2828
rect 16054 2788 16060 2800
rect 16112 2788 16118 2840
rect 18740 2828 18768 2859
rect 21114 2856 21120 2868
rect 21172 2856 21178 2908
rect 24981 2899 25039 2905
rect 24981 2865 24993 2899
rect 25027 2896 25039 2899
rect 26542 2896 26548 2908
rect 25027 2868 26548 2896
rect 25027 2865 25039 2868
rect 24981 2859 25039 2865
rect 26542 2856 26548 2868
rect 26600 2856 26606 2908
rect 28014 2896 28020 2908
rect 27975 2868 28020 2896
rect 28014 2856 28020 2868
rect 28072 2856 28078 2908
rect 17912 2800 18768 2828
rect 17912 2769 17940 2800
rect 23690 2788 23696 2840
rect 23748 2828 23754 2840
rect 26361 2831 26419 2837
rect 26361 2828 26373 2831
rect 23748 2800 26373 2828
rect 23748 2788 23754 2800
rect 26361 2797 26373 2800
rect 26407 2828 26419 2831
rect 26818 2828 26824 2840
rect 26407 2800 26824 2828
rect 26407 2797 26419 2800
rect 26361 2791 26419 2797
rect 26818 2788 26824 2800
rect 26876 2788 26882 2840
rect 28385 2831 28443 2837
rect 28385 2797 28397 2831
rect 28431 2828 28443 2831
rect 28842 2828 28848 2840
rect 28431 2800 28848 2828
rect 28431 2797 28443 2800
rect 28385 2791 28443 2797
rect 28842 2788 28848 2800
rect 28900 2788 28906 2840
rect 29302 2788 29308 2840
rect 29360 2828 29366 2840
rect 29765 2831 29823 2837
rect 29765 2828 29777 2831
rect 29360 2800 29777 2828
rect 29360 2788 29366 2800
rect 29765 2797 29777 2800
rect 29811 2797 29823 2831
rect 29765 2791 29823 2797
rect 17897 2763 17955 2769
rect 17897 2760 17909 2763
rect 4526 2732 5520 2760
rect 13404 2732 17909 2760
rect 4572 2704 4600 2732
rect 13404 2704 13432 2732
rect 17897 2729 17909 2732
rect 17943 2729 17955 2763
rect 19277 2763 19335 2769
rect 19277 2760 19289 2763
rect 17897 2723 17955 2729
rect 18464 2732 19289 2760
rect 18464 2704 18492 2732
rect 19277 2729 19289 2732
rect 19323 2729 19335 2763
rect 19277 2723 19335 2729
rect 1245 2695 1303 2701
rect 1245 2661 1257 2695
rect 1291 2692 1303 2695
rect 1702 2692 1708 2704
rect 1291 2664 1708 2692
rect 1291 2661 1303 2664
rect 1245 2655 1303 2661
rect 1702 2652 1708 2664
rect 1760 2652 1766 2704
rect 4554 2652 4560 2704
rect 4612 2652 4618 2704
rect 13386 2692 13392 2704
rect 13347 2664 13392 2692
rect 13386 2652 13392 2664
rect 13444 2652 13450 2704
rect 18446 2692 18452 2704
rect 18407 2664 18452 2692
rect 18446 2652 18452 2664
rect 18504 2652 18510 2704
rect 18630 2652 18636 2704
rect 18688 2692 18694 2704
rect 18909 2695 18967 2701
rect 18909 2692 18921 2695
rect 18688 2664 18921 2692
rect 18688 2652 18694 2664
rect 18909 2661 18921 2664
rect 18955 2661 18967 2695
rect 18909 2655 18967 2661
rect 19090 2652 19096 2704
rect 19148 2692 19154 2704
rect 19461 2695 19519 2701
rect 19461 2692 19473 2695
rect 19148 2664 19473 2692
rect 19148 2652 19154 2664
rect 19461 2661 19473 2664
rect 19507 2661 19519 2695
rect 19461 2655 19519 2661
rect 19734 2652 19740 2704
rect 19792 2692 19798 2704
rect 23598 2692 23604 2704
rect 19792 2664 23604 2692
rect 19792 2652 19798 2664
rect 23598 2652 23604 2664
rect 23656 2652 23662 2704
rect 25806 2692 25812 2704
rect 25767 2664 25812 2692
rect 25806 2652 25812 2664
rect 25864 2652 25870 2704
rect 400 2602 31680 2624
rect 400 2550 3510 2602
rect 3562 2550 3574 2602
rect 3626 2550 3638 2602
rect 3690 2550 3702 2602
rect 3754 2550 3766 2602
rect 3818 2550 31680 2602
rect 400 2528 31680 2550
rect 1058 2448 1064 2500
rect 1116 2448 1122 2500
rect 3358 2488 3364 2500
rect 3319 2460 3364 2488
rect 3358 2448 3364 2460
rect 3416 2448 3422 2500
rect 3910 2448 3916 2500
rect 3968 2488 3974 2500
rect 4373 2491 4431 2497
rect 4373 2488 4385 2491
rect 3968 2460 4385 2488
rect 3968 2448 3974 2460
rect 4373 2457 4385 2460
rect 4419 2457 4431 2491
rect 4373 2451 4431 2457
rect 5382 2448 5388 2500
rect 5440 2488 5446 2500
rect 5661 2491 5719 2497
rect 5661 2488 5673 2491
rect 5440 2460 5673 2488
rect 5440 2448 5446 2460
rect 5661 2457 5673 2460
rect 5707 2457 5719 2491
rect 6118 2488 6124 2500
rect 6079 2460 6124 2488
rect 5661 2451 5719 2457
rect 6118 2448 6124 2460
rect 6176 2448 6182 2500
rect 6854 2488 6860 2500
rect 6688 2460 6860 2488
rect 1076 2352 1104 2448
rect 3729 2423 3787 2429
rect 3729 2389 3741 2423
rect 3775 2420 3787 2423
rect 4462 2420 4468 2432
rect 3775 2392 4468 2420
rect 3775 2389 3787 2392
rect 3729 2383 3787 2389
rect 4462 2380 4468 2392
rect 4520 2420 4526 2432
rect 5477 2423 5535 2429
rect 5477 2420 5489 2423
rect 4520 2392 5489 2420
rect 4520 2380 4526 2392
rect 5477 2389 5489 2392
rect 5523 2420 5535 2423
rect 6026 2420 6032 2432
rect 5523 2392 6032 2420
rect 5523 2389 5535 2392
rect 5477 2383 5535 2389
rect 6026 2380 6032 2392
rect 6084 2380 6090 2432
rect 1245 2355 1303 2361
rect 1245 2352 1257 2355
rect 1076 2324 1257 2352
rect 1245 2321 1257 2324
rect 1291 2321 1303 2355
rect 1245 2315 1303 2321
rect 1702 2312 1708 2364
rect 1760 2352 1766 2364
rect 3545 2355 3603 2361
rect 1760 2324 2760 2352
rect 1760 2312 1766 2324
rect 966 2284 972 2296
rect 927 2256 972 2284
rect 966 2244 972 2256
rect 1024 2244 1030 2296
rect 2732 2284 2760 2324
rect 3545 2321 3557 2355
rect 3591 2352 3603 2355
rect 3591 2324 4140 2352
rect 3591 2321 3603 2324
rect 3545 2315 3603 2321
rect 3177 2287 3235 2293
rect 2732 2256 3128 2284
rect 1702 2176 1708 2228
rect 1760 2176 1766 2228
rect 2993 2219 3051 2225
rect 2993 2185 3005 2219
rect 3039 2185 3051 2219
rect 3100 2216 3128 2256
rect 3177 2253 3189 2287
rect 3223 2284 3235 2287
rect 3821 2287 3879 2293
rect 3821 2284 3833 2287
rect 3223 2256 3833 2284
rect 3223 2253 3235 2256
rect 3177 2247 3235 2253
rect 3821 2253 3833 2256
rect 3867 2284 3879 2287
rect 4002 2284 4008 2296
rect 3867 2256 4008 2284
rect 3867 2253 3879 2256
rect 3821 2247 3879 2253
rect 4002 2244 4008 2256
rect 4060 2244 4066 2296
rect 4112 2284 4140 2324
rect 4186 2312 4192 2364
rect 4244 2352 4250 2364
rect 6688 2361 6716 2460
rect 6854 2448 6860 2460
rect 6912 2488 6918 2500
rect 6949 2491 7007 2497
rect 6949 2488 6961 2491
rect 6912 2460 6961 2488
rect 6912 2448 6918 2460
rect 6949 2457 6961 2460
rect 6995 2457 7007 2491
rect 6949 2451 7007 2457
rect 9982 2448 9988 2500
rect 10040 2488 10046 2500
rect 10721 2491 10779 2497
rect 10721 2488 10733 2491
rect 10040 2460 10733 2488
rect 10040 2448 10046 2460
rect 10721 2457 10733 2460
rect 10767 2488 10779 2491
rect 11822 2488 11828 2500
rect 10767 2460 11828 2488
rect 10767 2457 10779 2460
rect 10721 2451 10779 2457
rect 11822 2448 11828 2460
rect 11880 2448 11886 2500
rect 12469 2491 12527 2497
rect 12469 2457 12481 2491
rect 12515 2488 12527 2491
rect 13386 2488 13392 2500
rect 12515 2460 13392 2488
rect 12515 2457 12527 2460
rect 12469 2451 12527 2457
rect 13386 2448 13392 2460
rect 13444 2448 13450 2500
rect 15502 2448 15508 2500
rect 15560 2488 15566 2500
rect 15689 2491 15747 2497
rect 15689 2488 15701 2491
rect 15560 2460 15701 2488
rect 15560 2448 15566 2460
rect 15689 2457 15701 2460
rect 15735 2457 15747 2491
rect 15689 2451 15747 2457
rect 15965 2491 16023 2497
rect 15965 2457 15977 2491
rect 16011 2488 16023 2491
rect 16054 2488 16060 2500
rect 16011 2460 16060 2488
rect 16011 2457 16023 2460
rect 15965 2451 16023 2457
rect 16054 2448 16060 2460
rect 16112 2488 16118 2500
rect 16609 2491 16667 2497
rect 16609 2488 16621 2491
rect 16112 2460 16621 2488
rect 16112 2448 16118 2460
rect 16609 2457 16621 2460
rect 16655 2488 16667 2491
rect 17158 2488 17164 2500
rect 16655 2460 17164 2488
rect 16655 2457 16667 2460
rect 16609 2451 16667 2457
rect 17158 2448 17164 2460
rect 17216 2448 17222 2500
rect 19366 2488 19372 2500
rect 18464 2460 19372 2488
rect 10537 2423 10595 2429
rect 10537 2389 10549 2423
rect 10583 2420 10595 2423
rect 11730 2420 11736 2432
rect 10583 2392 11736 2420
rect 10583 2389 10595 2392
rect 10537 2383 10595 2389
rect 11730 2380 11736 2392
rect 11788 2380 11794 2432
rect 16793 2423 16851 2429
rect 16793 2389 16805 2423
rect 16839 2420 16851 2423
rect 17066 2420 17072 2432
rect 16839 2392 17072 2420
rect 16839 2389 16851 2392
rect 16793 2383 16851 2389
rect 17066 2380 17072 2392
rect 17124 2380 17130 2432
rect 18464 2429 18492 2460
rect 19366 2448 19372 2460
rect 19424 2488 19430 2500
rect 21206 2488 21212 2500
rect 19424 2460 21212 2488
rect 19424 2448 19430 2460
rect 21206 2448 21212 2460
rect 21264 2448 21270 2500
rect 21298 2448 21304 2500
rect 21356 2488 21362 2500
rect 21485 2491 21543 2497
rect 21485 2488 21497 2491
rect 21356 2460 21497 2488
rect 21356 2448 21362 2460
rect 21485 2457 21497 2460
rect 21531 2457 21543 2491
rect 21485 2451 21543 2457
rect 23230 2448 23236 2500
rect 23288 2488 23294 2500
rect 24426 2488 24432 2500
rect 23288 2460 24432 2488
rect 23288 2448 23294 2460
rect 24426 2448 24432 2460
rect 24484 2448 24490 2500
rect 25438 2448 25444 2500
rect 25496 2488 25502 2500
rect 25809 2491 25867 2497
rect 25809 2488 25821 2491
rect 25496 2460 25821 2488
rect 25496 2448 25502 2460
rect 25809 2457 25821 2460
rect 25855 2488 25867 2491
rect 27278 2488 27284 2500
rect 25855 2460 27284 2488
rect 25855 2457 25867 2460
rect 25809 2451 25867 2457
rect 17345 2423 17403 2429
rect 17345 2389 17357 2423
rect 17391 2420 17403 2423
rect 18449 2423 18507 2429
rect 18449 2420 18461 2423
rect 17391 2392 18461 2420
rect 17391 2389 17403 2392
rect 17345 2383 17403 2389
rect 18449 2389 18461 2392
rect 18495 2389 18507 2423
rect 18449 2383 18507 2389
rect 21114 2380 21120 2432
rect 21172 2420 21178 2432
rect 21669 2423 21727 2429
rect 21669 2420 21681 2423
rect 21172 2392 21681 2420
rect 21172 2380 21178 2392
rect 21669 2389 21681 2392
rect 21715 2420 21727 2423
rect 22957 2423 23015 2429
rect 22957 2420 22969 2423
rect 21715 2392 22969 2420
rect 21715 2389 21727 2392
rect 21669 2383 21727 2389
rect 22957 2389 22969 2392
rect 23003 2389 23015 2423
rect 22957 2383 23015 2389
rect 4557 2355 4615 2361
rect 4557 2352 4569 2355
rect 4244 2324 4569 2352
rect 4244 2312 4250 2324
rect 4557 2321 4569 2324
rect 4603 2321 4615 2355
rect 4557 2315 4615 2321
rect 5937 2355 5995 2361
rect 5937 2321 5949 2355
rect 5983 2352 5995 2355
rect 6673 2355 6731 2361
rect 6673 2352 6685 2355
rect 5983 2324 6685 2352
rect 5983 2321 5995 2324
rect 5937 2315 5995 2321
rect 6673 2321 6685 2324
rect 6719 2321 6731 2355
rect 9246 2352 9252 2364
rect 6673 2315 6731 2321
rect 7700 2324 9252 2352
rect 4112 2256 4232 2284
rect 4094 2216 4100 2228
rect 3100 2188 4100 2216
rect 2993 2179 3051 2185
rect 877 2151 935 2157
rect 877 2117 889 2151
rect 923 2148 935 2151
rect 3008 2148 3036 2179
rect 4094 2176 4100 2188
rect 4152 2176 4158 2228
rect 4204 2216 4232 2256
rect 4278 2244 4284 2296
rect 4336 2284 4342 2296
rect 6397 2287 6455 2293
rect 6397 2284 6409 2287
rect 4336 2256 6409 2284
rect 4336 2244 4342 2256
rect 6397 2253 6409 2256
rect 6443 2284 6455 2287
rect 6762 2284 6768 2296
rect 6443 2256 6768 2284
rect 6443 2253 6455 2256
rect 6397 2247 6455 2253
rect 6762 2244 6768 2256
rect 6820 2284 6826 2296
rect 7133 2287 7191 2293
rect 7133 2284 7145 2287
rect 6820 2256 7145 2284
rect 6820 2244 6826 2256
rect 7133 2253 7145 2256
rect 7179 2253 7191 2287
rect 7133 2247 7191 2253
rect 4646 2216 4652 2228
rect 4204 2188 4652 2216
rect 4646 2176 4652 2188
rect 4704 2176 4710 2228
rect 3266 2148 3272 2160
rect 923 2120 3272 2148
rect 923 2117 935 2120
rect 877 2111 935 2117
rect 3266 2108 3272 2120
rect 3324 2108 3330 2160
rect 7222 2108 7228 2160
rect 7280 2148 7286 2160
rect 7700 2157 7728 2324
rect 9246 2312 9252 2324
rect 9304 2352 9310 2364
rect 9801 2355 9859 2361
rect 9801 2352 9813 2355
rect 9304 2324 9813 2352
rect 9304 2312 9310 2324
rect 9801 2321 9813 2324
rect 9847 2321 9859 2355
rect 9801 2315 9859 2321
rect 12653 2355 12711 2361
rect 12653 2321 12665 2355
rect 12699 2352 12711 2355
rect 13389 2355 13447 2361
rect 13389 2352 13401 2355
rect 12699 2324 13401 2352
rect 12699 2321 12711 2324
rect 12653 2315 12711 2321
rect 13389 2321 13401 2324
rect 13435 2352 13447 2355
rect 13478 2352 13484 2364
rect 13435 2324 13484 2352
rect 13435 2321 13447 2324
rect 13389 2315 13447 2321
rect 13478 2312 13484 2324
rect 13536 2312 13542 2364
rect 16882 2352 16888 2364
rect 16843 2324 16888 2352
rect 16882 2312 16888 2324
rect 16940 2352 16946 2364
rect 18173 2355 18231 2361
rect 16940 2324 17480 2352
rect 16940 2312 16946 2324
rect 8050 2284 8056 2296
rect 8011 2256 8056 2284
rect 8050 2244 8056 2256
rect 8108 2244 8114 2296
rect 8142 2244 8148 2296
rect 8200 2284 8206 2296
rect 8421 2287 8479 2293
rect 8421 2284 8433 2287
rect 8200 2256 8433 2284
rect 8200 2244 8206 2256
rect 8421 2253 8433 2256
rect 8467 2253 8479 2287
rect 8421 2247 8479 2253
rect 10350 2244 10356 2296
rect 10408 2284 10414 2296
rect 10905 2287 10963 2293
rect 10905 2284 10917 2287
rect 10408 2256 10917 2284
rect 10408 2244 10414 2256
rect 10905 2253 10917 2256
rect 10951 2284 10963 2287
rect 11178 2284 11184 2296
rect 10951 2256 11184 2284
rect 10951 2253 10963 2256
rect 10905 2247 10963 2253
rect 11178 2244 11184 2256
rect 11236 2284 11242 2296
rect 17452 2293 17480 2324
rect 18173 2321 18185 2355
rect 18219 2352 18231 2355
rect 18354 2352 18360 2364
rect 18219 2324 18360 2352
rect 18219 2321 18231 2324
rect 18173 2315 18231 2321
rect 18354 2312 18360 2324
rect 18412 2352 18418 2364
rect 19001 2355 19059 2361
rect 19001 2352 19013 2355
rect 18412 2324 19013 2352
rect 18412 2312 18418 2324
rect 19001 2321 19013 2324
rect 19047 2321 19059 2355
rect 19001 2315 19059 2321
rect 21022 2312 21028 2364
rect 21080 2352 21086 2364
rect 21301 2355 21359 2361
rect 21301 2352 21313 2355
rect 21080 2324 21313 2352
rect 21080 2312 21086 2324
rect 21301 2321 21313 2324
rect 21347 2321 21359 2355
rect 21301 2315 21359 2321
rect 13113 2287 13171 2293
rect 13113 2284 13125 2287
rect 11236 2256 13125 2284
rect 11236 2244 11242 2256
rect 13113 2253 13125 2256
rect 13159 2253 13171 2287
rect 17345 2287 17403 2293
rect 17345 2284 17357 2287
rect 13113 2247 13171 2253
rect 15060 2256 17357 2284
rect 9798 2216 9804 2228
rect 9448 2188 9804 2216
rect 7685 2151 7743 2157
rect 7685 2148 7697 2151
rect 7280 2120 7697 2148
rect 7280 2108 7286 2120
rect 7685 2117 7697 2120
rect 7731 2117 7743 2151
rect 7685 2111 7743 2117
rect 7961 2151 8019 2157
rect 7961 2117 7973 2151
rect 8007 2148 8019 2151
rect 9448 2148 9476 2188
rect 9798 2176 9804 2188
rect 9856 2216 9862 2228
rect 10261 2219 10319 2225
rect 10261 2216 10273 2219
rect 9856 2188 10273 2216
rect 9856 2176 9862 2188
rect 10261 2185 10273 2188
rect 10307 2216 10319 2219
rect 11086 2216 11092 2228
rect 10307 2188 11092 2216
rect 10307 2185 10319 2188
rect 10261 2179 10319 2185
rect 11086 2176 11092 2188
rect 11144 2216 11150 2228
rect 13128 2216 13156 2247
rect 13478 2216 13484 2228
rect 11144 2188 13064 2216
rect 13128 2188 13484 2216
rect 11144 2176 11150 2188
rect 8007 2120 9476 2148
rect 8007 2117 8019 2120
rect 7961 2111 8019 2117
rect 11730 2108 11736 2160
rect 11788 2148 11794 2160
rect 13036 2157 13064 2188
rect 13478 2176 13484 2188
rect 13536 2176 13542 2228
rect 12745 2151 12803 2157
rect 12745 2148 12757 2151
rect 11788 2120 12757 2148
rect 11788 2108 11794 2120
rect 12745 2117 12757 2120
rect 12791 2117 12803 2151
rect 12745 2111 12803 2117
rect 13021 2151 13079 2157
rect 13021 2117 13033 2151
rect 13067 2148 13079 2151
rect 14416 2148 14444 2216
rect 15060 2148 15088 2256
rect 17345 2253 17357 2256
rect 17391 2253 17403 2287
rect 17345 2247 17403 2253
rect 17437 2287 17495 2293
rect 17437 2253 17449 2287
rect 17483 2284 17495 2287
rect 17897 2287 17955 2293
rect 17897 2284 17909 2287
rect 17483 2256 17909 2284
rect 17483 2253 17495 2256
rect 17437 2247 17495 2253
rect 17897 2253 17909 2256
rect 17943 2284 17955 2287
rect 18446 2284 18452 2296
rect 17943 2256 18452 2284
rect 17943 2253 17955 2256
rect 17897 2247 17955 2253
rect 18446 2244 18452 2256
rect 18504 2244 18510 2296
rect 18538 2244 18544 2296
rect 18596 2284 18602 2296
rect 18633 2287 18691 2293
rect 18633 2284 18645 2287
rect 18596 2256 18645 2284
rect 18596 2244 18602 2256
rect 18633 2253 18645 2256
rect 18679 2284 18691 2287
rect 19090 2284 19096 2296
rect 18679 2256 19096 2284
rect 18679 2253 18691 2256
rect 18633 2247 18691 2253
rect 19090 2244 19096 2256
rect 19148 2244 19154 2296
rect 22972 2284 23000 2383
rect 23322 2312 23328 2364
rect 23380 2352 23386 2364
rect 23785 2355 23843 2361
rect 23785 2352 23797 2355
rect 23380 2324 23797 2352
rect 23380 2312 23386 2324
rect 23785 2321 23797 2324
rect 23831 2321 23843 2355
rect 23785 2315 23843 2321
rect 25533 2355 25591 2361
rect 25533 2321 25545 2355
rect 25579 2352 25591 2355
rect 25806 2352 25812 2364
rect 25579 2324 25812 2352
rect 25579 2321 25591 2324
rect 25533 2315 25591 2321
rect 23414 2284 23420 2296
rect 22972 2256 23420 2284
rect 23414 2244 23420 2256
rect 23472 2284 23478 2296
rect 23509 2287 23567 2293
rect 23509 2284 23521 2287
rect 23472 2256 23521 2284
rect 23472 2244 23478 2256
rect 23509 2253 23521 2256
rect 23555 2253 23567 2287
rect 23509 2247 23567 2253
rect 15137 2219 15195 2225
rect 15137 2185 15149 2219
rect 15183 2216 15195 2219
rect 15597 2219 15655 2225
rect 15597 2216 15609 2219
rect 15183 2188 15609 2216
rect 15183 2185 15195 2188
rect 15137 2179 15195 2185
rect 15597 2185 15609 2188
rect 15643 2216 15655 2219
rect 15686 2216 15692 2228
rect 15643 2188 15692 2216
rect 15643 2185 15655 2188
rect 15597 2179 15655 2185
rect 15686 2176 15692 2188
rect 15744 2216 15750 2228
rect 18170 2216 18176 2228
rect 15744 2188 18176 2216
rect 15744 2176 15750 2188
rect 18170 2176 18176 2188
rect 18228 2176 18234 2228
rect 18357 2219 18415 2225
rect 18357 2185 18369 2219
rect 18403 2216 18415 2219
rect 18403 2188 18768 2216
rect 18403 2185 18415 2188
rect 18357 2179 18415 2185
rect 13067 2120 15088 2148
rect 17161 2151 17219 2157
rect 13067 2117 13079 2120
rect 13021 2111 13079 2117
rect 17161 2117 17173 2151
rect 17207 2148 17219 2151
rect 17526 2148 17532 2160
rect 17207 2120 17532 2148
rect 17207 2117 17219 2120
rect 17161 2111 17219 2117
rect 17526 2108 17532 2120
rect 17584 2108 17590 2160
rect 18740 2148 18768 2188
rect 19366 2176 19372 2228
rect 19424 2176 19430 2228
rect 22494 2176 22500 2228
rect 22552 2216 22558 2228
rect 23138 2216 23144 2228
rect 22552 2188 23144 2216
rect 22552 2176 22558 2188
rect 23138 2176 23144 2188
rect 23196 2216 23202 2228
rect 23196 2188 23874 2216
rect 23196 2176 23202 2188
rect 19458 2148 19464 2160
rect 18740 2120 19464 2148
rect 19458 2108 19464 2120
rect 19516 2148 19522 2160
rect 20746 2148 20752 2160
rect 19516 2120 20752 2148
rect 19516 2108 19522 2120
rect 20746 2108 20752 2120
rect 20804 2108 20810 2160
rect 23322 2148 23328 2160
rect 23283 2120 23328 2148
rect 23322 2108 23328 2120
rect 23380 2108 23386 2160
rect 23846 2148 23874 2188
rect 24426 2176 24432 2228
rect 24484 2176 24490 2228
rect 25548 2148 25576 2315
rect 25806 2312 25812 2324
rect 25864 2312 25870 2364
rect 26818 2352 26824 2364
rect 26779 2324 26824 2352
rect 26818 2312 26824 2324
rect 26876 2312 26882 2364
rect 27020 2293 27048 2460
rect 27278 2448 27284 2460
rect 27336 2448 27342 2500
rect 28661 2491 28719 2497
rect 28661 2457 28673 2491
rect 28707 2488 28719 2491
rect 28842 2488 28848 2500
rect 28707 2460 28848 2488
rect 28707 2457 28719 2460
rect 28661 2451 28719 2457
rect 28842 2448 28848 2460
rect 28900 2448 28906 2500
rect 27462 2380 27468 2432
rect 27520 2420 27526 2432
rect 28017 2423 28075 2429
rect 28017 2420 28029 2423
rect 27520 2392 28029 2420
rect 27520 2380 27526 2392
rect 28017 2389 28029 2392
rect 28063 2420 28075 2423
rect 28198 2420 28204 2432
rect 28063 2392 28204 2420
rect 28063 2389 28075 2392
rect 28017 2383 28075 2389
rect 28198 2380 28204 2392
rect 28256 2380 28262 2432
rect 29578 2352 29584 2364
rect 27388 2324 29584 2352
rect 27388 2296 27416 2324
rect 29578 2312 29584 2324
rect 29636 2312 29642 2364
rect 27005 2287 27063 2293
rect 27005 2253 27017 2287
rect 27051 2253 27063 2287
rect 27370 2284 27376 2296
rect 27331 2256 27376 2284
rect 27005 2247 27063 2253
rect 27370 2244 27376 2256
rect 27428 2244 27434 2296
rect 27557 2287 27615 2293
rect 27557 2253 27569 2287
rect 27603 2284 27615 2287
rect 27738 2284 27744 2296
rect 27603 2256 27744 2284
rect 27603 2253 27615 2256
rect 27557 2247 27615 2253
rect 27738 2244 27744 2256
rect 27796 2244 27802 2296
rect 28014 2244 28020 2296
rect 28072 2284 28078 2296
rect 28753 2287 28811 2293
rect 28753 2284 28765 2287
rect 28072 2256 28765 2284
rect 28072 2244 28078 2256
rect 28753 2253 28765 2256
rect 28799 2253 28811 2287
rect 28753 2247 28811 2253
rect 25622 2176 25628 2228
rect 25680 2216 25686 2228
rect 26085 2219 26143 2225
rect 25680 2188 25944 2216
rect 25680 2176 25686 2188
rect 23846 2120 25576 2148
rect 25916 2148 25944 2188
rect 26085 2185 26097 2219
rect 26131 2216 26143 2219
rect 26361 2219 26419 2225
rect 26361 2216 26373 2219
rect 26131 2188 26373 2216
rect 26131 2185 26143 2188
rect 26085 2179 26143 2185
rect 26361 2185 26373 2188
rect 26407 2216 26419 2219
rect 27830 2216 27836 2228
rect 26407 2188 27836 2216
rect 26407 2185 26419 2188
rect 26361 2179 26419 2185
rect 27830 2176 27836 2188
rect 27888 2176 27894 2228
rect 28293 2219 28351 2225
rect 28293 2185 28305 2219
rect 28339 2216 28351 2219
rect 28382 2216 28388 2228
rect 28339 2188 28388 2216
rect 28339 2185 28351 2188
rect 28293 2179 28351 2185
rect 28382 2176 28388 2188
rect 28440 2216 28446 2228
rect 29302 2216 29308 2228
rect 28440 2188 29308 2216
rect 28440 2176 28446 2188
rect 29302 2176 29308 2188
rect 29360 2176 29366 2228
rect 26269 2151 26327 2157
rect 26269 2148 26281 2151
rect 25916 2120 26281 2148
rect 26269 2117 26281 2120
rect 26315 2148 26327 2151
rect 27738 2148 27744 2160
rect 26315 2120 27744 2148
rect 26315 2117 26327 2120
rect 26269 2111 26327 2117
rect 27738 2108 27744 2120
rect 27796 2108 27802 2160
rect 400 2058 31680 2080
rect 400 2006 18870 2058
rect 18922 2006 18934 2058
rect 18986 2006 18998 2058
rect 19050 2006 19062 2058
rect 19114 2006 19126 2058
rect 19178 2006 31680 2058
rect 400 1984 31680 2006
rect 966 1904 972 1956
rect 1024 1944 1030 1956
rect 1245 1947 1303 1953
rect 1245 1944 1257 1947
rect 1024 1916 1257 1944
rect 1024 1904 1030 1916
rect 1245 1913 1257 1916
rect 1291 1913 1303 1947
rect 1245 1907 1303 1913
rect 1150 1808 1156 1820
rect 1111 1780 1156 1808
rect 1150 1768 1156 1780
rect 1208 1768 1214 1820
rect 1260 1740 1288 1907
rect 1702 1904 1708 1956
rect 1760 1944 1766 1956
rect 5566 1944 5572 1956
rect 1760 1916 5572 1944
rect 1760 1904 1766 1916
rect 5566 1904 5572 1916
rect 5624 1904 5630 1956
rect 8050 1904 8056 1956
rect 8108 1944 8114 1956
rect 8145 1947 8203 1953
rect 8145 1944 8157 1947
rect 8108 1916 8157 1944
rect 8108 1904 8114 1916
rect 8145 1913 8157 1916
rect 8191 1944 8203 1947
rect 9706 1944 9712 1956
rect 8191 1916 9712 1944
rect 8191 1913 8203 1916
rect 8145 1907 8203 1913
rect 9706 1904 9712 1916
rect 9764 1944 9770 1956
rect 10350 1944 10356 1956
rect 9764 1916 10356 1944
rect 9764 1904 9770 1916
rect 10350 1904 10356 1916
rect 10408 1904 10414 1956
rect 13205 1947 13263 1953
rect 13205 1913 13217 1947
rect 13251 1944 13263 1947
rect 13570 1944 13576 1956
rect 13251 1916 13576 1944
rect 13251 1913 13263 1916
rect 13205 1907 13263 1913
rect 13570 1904 13576 1916
rect 13628 1904 13634 1956
rect 16974 1944 16980 1956
rect 16935 1916 16980 1944
rect 16974 1904 16980 1916
rect 17032 1904 17038 1956
rect 18354 1944 18360 1956
rect 18315 1916 18360 1944
rect 18354 1904 18360 1916
rect 18412 1904 18418 1956
rect 18446 1904 18452 1956
rect 18504 1944 18510 1956
rect 19369 1947 19427 1953
rect 19369 1944 19381 1947
rect 18504 1916 19381 1944
rect 18504 1904 18510 1916
rect 3910 1836 3916 1888
rect 3968 1876 3974 1888
rect 4189 1879 4247 1885
rect 4189 1876 4201 1879
rect 3968 1848 4201 1876
rect 3968 1836 3974 1848
rect 4189 1845 4201 1848
rect 4235 1845 4247 1879
rect 4189 1839 4247 1845
rect 4646 1836 4652 1888
rect 4704 1836 4710 1888
rect 5842 1836 5848 1888
rect 5900 1876 5906 1888
rect 5937 1879 5995 1885
rect 5937 1876 5949 1879
rect 5900 1848 5949 1876
rect 5900 1836 5906 1848
rect 5937 1845 5949 1848
rect 5983 1845 5995 1879
rect 5937 1839 5995 1845
rect 6762 1808 6768 1820
rect 6723 1780 6768 1808
rect 6762 1768 6768 1780
rect 6820 1768 6826 1820
rect 9724 1817 9752 1904
rect 13110 1836 13116 1888
rect 13168 1876 13174 1888
rect 13297 1879 13355 1885
rect 13297 1876 13309 1879
rect 13168 1848 13309 1876
rect 13168 1836 13174 1848
rect 13297 1845 13309 1848
rect 13343 1845 13355 1879
rect 13478 1876 13484 1888
rect 13391 1848 13484 1876
rect 13297 1839 13355 1845
rect 13478 1836 13484 1848
rect 13536 1876 13542 1888
rect 17805 1879 17863 1885
rect 17805 1876 17817 1879
rect 13536 1848 17817 1876
rect 13536 1836 13542 1848
rect 17805 1845 17817 1848
rect 17851 1845 17863 1879
rect 17805 1839 17863 1845
rect 17989 1879 18047 1885
rect 17989 1845 18001 1879
rect 18035 1876 18047 1879
rect 18630 1876 18636 1888
rect 18035 1848 18636 1876
rect 18035 1845 18047 1848
rect 17989 1839 18047 1845
rect 18630 1836 18636 1848
rect 18688 1836 18694 1888
rect 18740 1820 18768 1916
rect 19369 1913 19381 1916
rect 19415 1913 19427 1947
rect 19369 1907 19427 1913
rect 20197 1947 20255 1953
rect 20197 1913 20209 1947
rect 20243 1944 20255 1947
rect 26453 1947 26511 1953
rect 20243 1916 21804 1944
rect 20243 1913 20255 1916
rect 20197 1907 20255 1913
rect 9709 1811 9767 1817
rect 9709 1777 9721 1811
rect 9755 1777 9767 1811
rect 9709 1771 9767 1777
rect 11086 1768 11092 1820
rect 11144 1768 11150 1820
rect 18446 1808 18452 1820
rect 14186 1780 18452 1808
rect 3913 1743 3971 1749
rect 3913 1740 3925 1743
rect 1260 1712 3925 1740
rect 3913 1709 3925 1712
rect 3959 1740 3971 1743
rect 4554 1740 4560 1752
rect 3959 1712 4560 1740
rect 3959 1709 3971 1712
rect 3913 1703 3971 1709
rect 4554 1700 4560 1712
rect 4612 1700 4618 1752
rect 6946 1740 6952 1752
rect 6907 1712 6952 1740
rect 6946 1700 6952 1712
rect 7004 1700 7010 1752
rect 9985 1743 10043 1749
rect 9985 1709 9997 1743
rect 10031 1740 10043 1743
rect 10074 1740 10080 1752
rect 10031 1712 10080 1740
rect 10031 1709 10043 1712
rect 9985 1703 10043 1709
rect 10074 1700 10080 1712
rect 10132 1740 10138 1752
rect 11270 1740 11276 1752
rect 10132 1712 11276 1740
rect 10132 1700 10138 1712
rect 11270 1700 11276 1712
rect 11328 1700 11334 1752
rect 11730 1740 11736 1752
rect 11691 1712 11736 1740
rect 11730 1700 11736 1712
rect 11788 1700 11794 1752
rect 13938 1700 13944 1752
rect 13996 1740 14002 1752
rect 14186 1740 14214 1780
rect 18446 1768 18452 1780
rect 18504 1808 18510 1820
rect 18541 1811 18599 1817
rect 18541 1808 18553 1811
rect 18504 1780 18553 1808
rect 18504 1768 18510 1780
rect 18541 1777 18553 1780
rect 18587 1777 18599 1811
rect 18722 1808 18728 1820
rect 18635 1780 18728 1808
rect 18541 1771 18599 1777
rect 18722 1768 18728 1780
rect 18780 1768 18786 1820
rect 19090 1808 19096 1820
rect 19003 1780 19096 1808
rect 19090 1768 19096 1780
rect 19148 1808 19154 1820
rect 20194 1808 20200 1820
rect 19148 1780 20200 1808
rect 19148 1768 19154 1780
rect 20194 1768 20200 1780
rect 20252 1768 20258 1820
rect 20304 1817 20332 1916
rect 21776 1888 21804 1916
rect 26453 1913 26465 1947
rect 26499 1944 26511 1947
rect 27370 1944 27376 1956
rect 26499 1916 27376 1944
rect 26499 1913 26511 1916
rect 26453 1907 26511 1913
rect 27370 1904 27376 1916
rect 27428 1904 27434 1956
rect 21206 1836 21212 1888
rect 21264 1836 21270 1888
rect 21758 1836 21764 1888
rect 21816 1876 21822 1888
rect 21816 1848 27508 1876
rect 21816 1836 21822 1848
rect 20289 1811 20347 1817
rect 20289 1777 20301 1811
rect 20335 1777 20347 1811
rect 20289 1771 20347 1777
rect 23046 1768 23052 1820
rect 23104 1808 23110 1820
rect 23104 1780 23828 1808
rect 23104 1768 23110 1780
rect 13996 1712 14214 1740
rect 13996 1700 14002 1712
rect 17342 1700 17348 1752
rect 17400 1740 17406 1752
rect 18170 1740 18176 1752
rect 17400 1712 18176 1740
rect 17400 1700 17406 1712
rect 18170 1700 18176 1712
rect 18228 1740 18234 1752
rect 19001 1743 19059 1749
rect 19001 1740 19013 1743
rect 18228 1712 19013 1740
rect 18228 1700 18234 1712
rect 19001 1709 19013 1712
rect 19047 1740 19059 1743
rect 19458 1740 19464 1752
rect 19047 1712 19464 1740
rect 19047 1709 19059 1712
rect 19001 1703 19059 1709
rect 19458 1700 19464 1712
rect 19516 1700 19522 1752
rect 20654 1740 20660 1752
rect 20615 1712 20660 1740
rect 20654 1700 20660 1712
rect 20712 1700 20718 1752
rect 22034 1740 22040 1752
rect 21995 1712 22040 1740
rect 22034 1700 22040 1712
rect 22092 1700 22098 1752
rect 22586 1700 22592 1752
rect 22644 1740 22650 1752
rect 23690 1740 23696 1752
rect 22644 1712 23696 1740
rect 22644 1700 22650 1712
rect 23690 1700 23696 1712
rect 23748 1700 23754 1752
rect 23800 1740 23828 1780
rect 23874 1768 23880 1820
rect 23932 1808 23938 1820
rect 23932 1780 23977 1808
rect 23932 1768 23938 1780
rect 24058 1768 24064 1820
rect 24116 1808 24122 1820
rect 24245 1811 24303 1817
rect 24245 1808 24257 1811
rect 24116 1780 24257 1808
rect 24116 1768 24122 1780
rect 24245 1777 24257 1780
rect 24291 1777 24303 1811
rect 24245 1771 24303 1777
rect 24429 1811 24487 1817
rect 24429 1777 24441 1811
rect 24475 1808 24487 1811
rect 24794 1808 24800 1820
rect 24475 1780 24800 1808
rect 24475 1777 24487 1780
rect 24429 1771 24487 1777
rect 24444 1740 24472 1771
rect 24794 1768 24800 1780
rect 24852 1768 24858 1820
rect 27480 1749 27508 1848
rect 28198 1836 28204 1888
rect 28256 1836 28262 1888
rect 27830 1808 27836 1820
rect 27791 1780 27836 1808
rect 27830 1768 27836 1780
rect 27888 1768 27894 1820
rect 23800 1712 24472 1740
rect 27465 1743 27523 1749
rect 27465 1709 27477 1743
rect 27511 1740 27523 1743
rect 28014 1740 28020 1752
rect 27511 1712 28020 1740
rect 27511 1709 27523 1712
rect 27465 1703 27523 1709
rect 28014 1700 28020 1712
rect 28072 1700 28078 1752
rect 17805 1675 17863 1681
rect 17805 1641 17817 1675
rect 17851 1672 17863 1675
rect 18538 1672 18544 1684
rect 17851 1644 18544 1672
rect 17851 1641 17863 1644
rect 17805 1635 17863 1641
rect 18538 1632 18544 1644
rect 18596 1672 18602 1684
rect 20197 1675 20255 1681
rect 20197 1672 20209 1675
rect 18596 1644 20209 1672
rect 18596 1632 18602 1644
rect 20197 1641 20209 1644
rect 20243 1641 20255 1675
rect 22052 1672 22080 1700
rect 26542 1672 26548 1684
rect 22052 1644 26548 1672
rect 20197 1635 20255 1641
rect 26542 1632 26548 1644
rect 26600 1632 26606 1684
rect 2162 1604 2168 1616
rect 2123 1576 2168 1604
rect 2162 1564 2168 1576
rect 2220 1564 2226 1616
rect 12742 1604 12748 1616
rect 12703 1576 12748 1604
rect 12742 1564 12748 1576
rect 12800 1564 12806 1616
rect 15134 1604 15140 1616
rect 15095 1576 15140 1604
rect 15134 1564 15140 1576
rect 15192 1564 15198 1616
rect 16606 1564 16612 1616
rect 16664 1604 16670 1616
rect 16701 1607 16759 1613
rect 16701 1604 16713 1607
rect 16664 1576 16713 1604
rect 16664 1564 16670 1576
rect 16701 1573 16713 1576
rect 16747 1573 16759 1607
rect 16701 1567 16759 1573
rect 23509 1607 23567 1613
rect 23509 1573 23521 1607
rect 23555 1604 23567 1607
rect 23690 1604 23696 1616
rect 23555 1576 23696 1604
rect 23555 1573 23567 1576
rect 23509 1567 23567 1573
rect 23690 1564 23696 1576
rect 23748 1564 23754 1616
rect 25990 1604 25996 1616
rect 25951 1576 25996 1604
rect 25990 1564 25996 1576
rect 26048 1564 26054 1616
rect 27738 1564 27744 1616
rect 27796 1604 27802 1616
rect 29581 1607 29639 1613
rect 29581 1604 29593 1607
rect 27796 1576 29593 1604
rect 27796 1564 27802 1576
rect 29581 1573 29593 1576
rect 29627 1604 29639 1607
rect 30774 1604 30780 1616
rect 29627 1576 30780 1604
rect 29627 1573 29639 1576
rect 29581 1567 29639 1573
rect 30774 1564 30780 1576
rect 30832 1564 30838 1616
rect 400 1514 31680 1536
rect 400 1462 3510 1514
rect 3562 1462 3574 1514
rect 3626 1462 3638 1514
rect 3690 1462 3702 1514
rect 3754 1462 3766 1514
rect 3818 1462 31680 1514
rect 400 1440 31680 1462
rect 1061 1403 1119 1409
rect 1061 1369 1073 1403
rect 1107 1400 1119 1403
rect 1150 1400 1156 1412
rect 1107 1372 1156 1400
rect 1107 1369 1119 1372
rect 1061 1363 1119 1369
rect 1150 1360 1156 1372
rect 1208 1360 1214 1412
rect 3910 1360 3916 1412
rect 3968 1400 3974 1412
rect 4097 1403 4155 1409
rect 4097 1400 4109 1403
rect 3968 1372 4109 1400
rect 3968 1360 3974 1372
rect 4097 1369 4109 1372
rect 4143 1369 4155 1403
rect 4097 1363 4155 1369
rect 4373 1403 4431 1409
rect 4373 1369 4385 1403
rect 4419 1400 4431 1403
rect 4646 1400 4652 1412
rect 4419 1372 4652 1400
rect 4419 1369 4431 1372
rect 4373 1363 4431 1369
rect 4646 1360 4652 1372
rect 4704 1400 4710 1412
rect 6765 1403 6823 1409
rect 6765 1400 6777 1403
rect 4704 1372 6777 1400
rect 4704 1360 4710 1372
rect 6765 1369 6777 1372
rect 6811 1400 6823 1403
rect 6946 1400 6952 1412
rect 6811 1372 6952 1400
rect 6811 1369 6823 1372
rect 6765 1363 6823 1369
rect 6946 1360 6952 1372
rect 7004 1360 7010 1412
rect 9798 1400 9804 1412
rect 9759 1372 9804 1400
rect 9798 1360 9804 1372
rect 9856 1360 9862 1412
rect 10074 1400 10080 1412
rect 10035 1372 10080 1400
rect 10074 1360 10080 1372
rect 10132 1360 10138 1412
rect 10350 1400 10356 1412
rect 10311 1372 10356 1400
rect 10350 1360 10356 1372
rect 10408 1360 10414 1412
rect 18170 1400 18176 1412
rect 18131 1372 18176 1400
rect 18170 1360 18176 1372
rect 18228 1360 18234 1412
rect 18446 1400 18452 1412
rect 18407 1372 18452 1400
rect 18446 1360 18452 1372
rect 18504 1360 18510 1412
rect 18722 1400 18728 1412
rect 18683 1372 18728 1400
rect 18722 1360 18728 1372
rect 18780 1360 18786 1412
rect 18909 1403 18967 1409
rect 18909 1369 18921 1403
rect 18955 1400 18967 1403
rect 19461 1403 19519 1409
rect 19461 1400 19473 1403
rect 18955 1372 19473 1400
rect 18955 1369 18967 1372
rect 18909 1363 18967 1369
rect 19461 1369 19473 1372
rect 19507 1400 19519 1403
rect 20654 1400 20660 1412
rect 19507 1372 20660 1400
rect 19507 1369 19519 1372
rect 19461 1363 19519 1369
rect 20654 1360 20660 1372
rect 20712 1400 20718 1412
rect 20841 1403 20899 1409
rect 20841 1400 20853 1403
rect 20712 1372 20853 1400
rect 20712 1360 20718 1372
rect 20841 1369 20853 1372
rect 20887 1369 20899 1403
rect 20841 1363 20899 1369
rect 21117 1403 21175 1409
rect 21117 1369 21129 1403
rect 21163 1400 21175 1403
rect 21758 1400 21764 1412
rect 21163 1372 21764 1400
rect 21163 1369 21175 1372
rect 21117 1363 21175 1369
rect 21758 1360 21764 1372
rect 21816 1360 21822 1412
rect 22405 1403 22463 1409
rect 22405 1369 22417 1403
rect 22451 1400 22463 1403
rect 24058 1400 24064 1412
rect 22451 1372 24064 1400
rect 22451 1369 22463 1372
rect 22405 1363 22463 1369
rect 24058 1360 24064 1372
rect 24116 1360 24122 1412
rect 24426 1360 24432 1412
rect 24484 1400 24490 1412
rect 27462 1400 27468 1412
rect 24484 1372 27468 1400
rect 24484 1360 24490 1372
rect 27462 1360 27468 1372
rect 27520 1360 27526 1412
rect 27830 1400 27836 1412
rect 27791 1372 27836 1400
rect 27830 1360 27836 1372
rect 27888 1360 27894 1412
rect 28014 1400 28020 1412
rect 27975 1372 28020 1400
rect 28014 1360 28020 1372
rect 28072 1360 28078 1412
rect 4005 1335 4063 1341
rect 4005 1301 4017 1335
rect 4051 1332 4063 1335
rect 5842 1332 5848 1344
rect 4051 1304 5848 1332
rect 4051 1301 4063 1304
rect 4005 1295 4063 1301
rect 5842 1292 5848 1304
rect 5900 1292 5906 1344
rect 9985 1335 10043 1341
rect 9985 1301 9997 1335
rect 10031 1332 10043 1335
rect 11730 1332 11736 1344
rect 10031 1304 11736 1332
rect 10031 1301 10043 1304
rect 9985 1295 10043 1301
rect 11730 1292 11736 1304
rect 11788 1292 11794 1344
rect 18354 1332 18360 1344
rect 18315 1304 18360 1332
rect 18354 1292 18360 1304
rect 18412 1292 18418 1344
rect 18740 1332 18768 1360
rect 22586 1332 22592 1344
rect 18740 1304 19872 1332
rect 22547 1304 22592 1332
rect 4554 1224 4560 1276
rect 4612 1264 4618 1276
rect 4612 1236 4657 1264
rect 4612 1224 4618 1236
rect 6762 1224 6768 1276
rect 6820 1264 6826 1276
rect 6949 1267 7007 1273
rect 6949 1264 6961 1267
rect 6820 1236 6961 1264
rect 6820 1224 6826 1236
rect 6949 1233 6961 1236
rect 6995 1233 7007 1267
rect 6949 1227 7007 1233
rect 17989 1267 18047 1273
rect 17989 1233 18001 1267
rect 18035 1264 18047 1267
rect 19090 1264 19096 1276
rect 18035 1236 19096 1264
rect 18035 1233 18047 1236
rect 17989 1227 18047 1233
rect 19090 1224 19096 1236
rect 19148 1224 19154 1276
rect 19642 1264 19648 1276
rect 19603 1236 19648 1264
rect 19642 1224 19648 1236
rect 19700 1224 19706 1276
rect 19844 1205 19872 1304
rect 22586 1292 22592 1304
rect 22644 1292 22650 1344
rect 23233 1335 23291 1341
rect 23233 1332 23245 1335
rect 22696 1304 23245 1332
rect 20565 1267 20623 1273
rect 20565 1233 20577 1267
rect 20611 1264 20623 1267
rect 21206 1264 21212 1276
rect 20611 1236 21212 1264
rect 20611 1233 20623 1236
rect 20565 1227 20623 1233
rect 21206 1224 21212 1236
rect 21264 1264 21270 1276
rect 22696 1264 22724 1304
rect 23233 1301 23245 1304
rect 23279 1332 23291 1335
rect 23322 1332 23328 1344
rect 23279 1304 23328 1332
rect 23279 1301 23291 1304
rect 23233 1295 23291 1301
rect 23322 1292 23328 1304
rect 23380 1292 23386 1344
rect 24794 1292 24800 1344
rect 24852 1332 24858 1344
rect 27738 1332 27744 1344
rect 24852 1304 25484 1332
rect 27699 1304 27744 1332
rect 24852 1292 24858 1304
rect 21264 1236 22724 1264
rect 22773 1267 22831 1273
rect 21264 1224 21270 1236
rect 22773 1233 22785 1267
rect 22819 1264 22831 1267
rect 23690 1264 23696 1276
rect 22819 1236 23696 1264
rect 22819 1233 22831 1236
rect 22773 1227 22831 1233
rect 23690 1224 23696 1236
rect 23748 1224 23754 1276
rect 25456 1273 25484 1304
rect 27738 1292 27744 1304
rect 27796 1292 27802 1344
rect 25441 1267 25499 1273
rect 25441 1233 25453 1267
rect 25487 1233 25499 1267
rect 25441 1227 25499 1233
rect 3545 1199 3603 1205
rect 3545 1165 3557 1199
rect 3591 1165 3603 1199
rect 3545 1159 3603 1165
rect 19829 1199 19887 1205
rect 19829 1165 19841 1199
rect 19875 1165 19887 1199
rect 20194 1196 20200 1208
rect 20155 1168 20200 1196
rect 19829 1159 19887 1165
rect 3560 1128 3588 1159
rect 20194 1156 20200 1168
rect 20252 1156 20258 1208
rect 20289 1199 20347 1205
rect 20289 1165 20301 1199
rect 20335 1196 20347 1199
rect 20657 1199 20715 1205
rect 20657 1196 20669 1199
rect 20335 1168 20669 1196
rect 20335 1165 20347 1168
rect 20289 1159 20347 1165
rect 20657 1165 20669 1168
rect 20703 1196 20715 1199
rect 22034 1196 22040 1208
rect 20703 1168 22040 1196
rect 20703 1165 20715 1168
rect 20657 1159 20715 1165
rect 3729 1131 3787 1137
rect 3729 1128 3741 1131
rect 3560 1100 3741 1128
rect 3729 1097 3741 1100
rect 3775 1128 3787 1131
rect 4462 1128 4468 1140
rect 3775 1100 4468 1128
rect 3775 1097 3787 1100
rect 3729 1091 3787 1097
rect 4462 1088 4468 1100
rect 4520 1088 4526 1140
rect 19093 1131 19151 1137
rect 19093 1097 19105 1131
rect 19139 1128 19151 1131
rect 19274 1128 19280 1140
rect 19139 1100 19280 1128
rect 19139 1097 19151 1100
rect 19093 1091 19151 1097
rect 19274 1088 19280 1100
rect 19332 1128 19338 1140
rect 20304 1128 20332 1159
rect 22034 1156 22040 1168
rect 22092 1156 22098 1208
rect 23414 1196 23420 1208
rect 23375 1168 23420 1196
rect 23414 1156 23420 1168
rect 23472 1156 23478 1208
rect 19332 1100 20332 1128
rect 19332 1088 19338 1100
rect 24426 1088 24432 1140
rect 24484 1088 24490 1140
rect 2073 1063 2131 1069
rect 2073 1029 2085 1063
rect 2119 1060 2131 1063
rect 2162 1060 2168 1072
rect 2119 1032 2168 1060
rect 2119 1029 2131 1032
rect 2073 1023 2131 1029
rect 2162 1020 2168 1032
rect 2220 1060 2226 1072
rect 3174 1060 3180 1072
rect 2220 1032 3180 1060
rect 2220 1020 2226 1032
rect 3174 1020 3180 1032
rect 3232 1020 3238 1072
rect 11454 1020 11460 1072
rect 11512 1060 11518 1072
rect 12561 1063 12619 1069
rect 12561 1060 12573 1063
rect 11512 1032 12573 1060
rect 11512 1020 11518 1032
rect 12561 1029 12573 1032
rect 12607 1060 12619 1063
rect 12742 1060 12748 1072
rect 12607 1032 12748 1060
rect 12607 1029 12619 1032
rect 12561 1023 12619 1029
rect 12742 1020 12748 1032
rect 12800 1020 12806 1072
rect 15045 1063 15103 1069
rect 15045 1029 15057 1063
rect 15091 1060 15103 1063
rect 15134 1060 15140 1072
rect 15091 1032 15140 1060
rect 15091 1029 15103 1032
rect 15045 1023 15103 1029
rect 15134 1020 15140 1032
rect 15192 1060 15198 1072
rect 15502 1060 15508 1072
rect 15192 1032 15508 1060
rect 15192 1020 15198 1032
rect 15502 1020 15508 1032
rect 15560 1020 15566 1072
rect 16606 1060 16612 1072
rect 16567 1032 16612 1060
rect 16606 1020 16612 1032
rect 16664 1020 16670 1072
rect 23046 1060 23052 1072
rect 23007 1032 23052 1060
rect 23046 1020 23052 1032
rect 23104 1020 23110 1072
rect 23782 1020 23788 1072
rect 23840 1060 23846 1072
rect 25809 1063 25867 1069
rect 25809 1060 25821 1063
rect 23840 1032 25821 1060
rect 23840 1020 23846 1032
rect 25809 1029 25821 1032
rect 25855 1060 25867 1063
rect 25990 1060 25996 1072
rect 25855 1032 25996 1060
rect 25855 1029 25867 1032
rect 25809 1023 25867 1029
rect 25990 1020 25996 1032
rect 26048 1020 26054 1072
rect 400 970 31680 992
rect 400 918 18870 970
rect 18922 918 18934 970
rect 18986 918 18998 970
rect 19050 918 19062 970
rect 19114 918 19126 970
rect 19178 918 31680 970
rect 400 896 31680 918
rect 19461 859 19519 865
rect 19461 825 19473 859
rect 19507 856 19519 859
rect 20194 856 20200 868
rect 19507 828 20200 856
rect 19507 825 19519 828
rect 19461 819 19519 825
rect 20194 816 20200 828
rect 20252 816 20258 868
rect 23690 856 23696 868
rect 23651 828 23696 856
rect 23690 816 23696 828
rect 23748 816 23754 868
rect 23874 816 23880 868
rect 23932 856 23938 868
rect 23932 828 23977 856
rect 23932 816 23938 828
rect 19277 791 19335 797
rect 19277 757 19289 791
rect 19323 788 19335 791
rect 19642 788 19648 800
rect 19323 760 19648 788
rect 19323 757 19335 760
rect 19277 751 19335 757
rect 19642 748 19648 760
rect 19700 748 19706 800
rect 23414 748 23420 800
rect 23472 788 23478 800
rect 23969 791 24027 797
rect 23969 788 23981 791
rect 23472 760 23981 788
rect 23472 748 23478 760
rect 23969 757 23981 760
rect 24015 757 24027 791
rect 23969 751 24027 757
rect 21022 476 21028 528
rect 21080 516 21086 528
rect 23046 516 23052 528
rect 21080 488 23052 516
rect 21080 476 21086 488
rect 23046 476 23052 488
rect 23104 516 23110 528
rect 23417 519 23475 525
rect 23417 516 23429 519
rect 23104 488 23429 516
rect 23104 476 23110 488
rect 23417 485 23429 488
rect 23463 485 23475 519
rect 23417 479 23475 485
rect 400 426 31680 448
rect 400 374 3510 426
rect 3562 374 3574 426
rect 3626 374 3638 426
rect 3690 374 3702 426
rect 3754 374 3766 426
rect 3818 374 31680 426
rect 400 352 31680 374
<< via1 >>
rect 18870 31382 18922 31434
rect 18934 31382 18986 31434
rect 18998 31382 19050 31434
rect 19062 31382 19114 31434
rect 19126 31382 19178 31434
rect 3510 30838 3562 30890
rect 3574 30838 3626 30890
rect 3638 30838 3690 30890
rect 3702 30838 3754 30890
rect 3766 30838 3818 30890
rect 2628 30668 2680 30720
rect 8608 30668 8660 30720
rect 1156 30600 1208 30652
rect 13392 30600 13444 30652
rect 19280 30600 19332 30652
rect 27468 30736 27520 30788
rect 4008 30532 4060 30584
rect 9988 30532 10040 30584
rect 5020 30507 5072 30516
rect 5020 30473 5029 30507
rect 5029 30473 5063 30507
rect 5063 30473 5072 30507
rect 5020 30464 5072 30473
rect 5388 30464 5440 30516
rect 9436 30464 9488 30516
rect 9896 30464 9948 30516
rect 16888 30464 16940 30516
rect 26916 30532 26968 30584
rect 28848 30507 28900 30516
rect 28848 30473 28857 30507
rect 28857 30473 28891 30507
rect 28891 30473 28900 30507
rect 28848 30464 28900 30473
rect 3916 30396 3968 30448
rect 10172 30396 10224 30448
rect 18360 30439 18412 30448
rect 18360 30405 18369 30439
rect 18369 30405 18403 30439
rect 18403 30405 18412 30439
rect 18360 30396 18412 30405
rect 18870 30294 18922 30346
rect 18934 30294 18986 30346
rect 18998 30294 19050 30346
rect 19062 30294 19114 30346
rect 19126 30294 19178 30346
rect 420 30192 472 30244
rect 6492 30192 6544 30244
rect 6676 30192 6728 30244
rect 7688 30192 7740 30244
rect 13668 30192 13720 30244
rect 14864 30192 14916 30244
rect 14956 30192 15008 30244
rect 18544 30192 18596 30244
rect 28848 30235 28900 30244
rect 28848 30201 28857 30235
rect 28857 30201 28891 30235
rect 28891 30201 28900 30235
rect 28848 30192 28900 30201
rect 4008 30167 4060 30176
rect 4008 30133 4017 30167
rect 4017 30133 4051 30167
rect 4051 30133 4060 30167
rect 4008 30124 4060 30133
rect 4468 30124 4520 30176
rect 5388 30124 5440 30176
rect 9160 30124 9212 30176
rect 10264 30124 10316 30176
rect 16888 30124 16940 30176
rect 6308 30056 6360 30108
rect 8976 30099 9028 30108
rect 8976 30065 8985 30099
rect 8985 30065 9019 30099
rect 9019 30065 9028 30099
rect 8976 30056 9028 30065
rect 12564 30099 12616 30108
rect 12564 30065 12573 30099
rect 12573 30065 12607 30099
rect 12607 30065 12616 30099
rect 12564 30056 12616 30065
rect 17716 30056 17768 30108
rect 19004 30056 19056 30108
rect 20476 30099 20528 30108
rect 20476 30065 20485 30099
rect 20485 30065 20519 30099
rect 20519 30065 20528 30099
rect 20476 30056 20528 30065
rect 23052 30099 23104 30108
rect 23052 30065 23061 30099
rect 23061 30065 23095 30099
rect 23095 30065 23104 30099
rect 23052 30056 23104 30065
rect 24524 30056 24576 30108
rect 24616 30056 24668 30108
rect 27836 30056 27888 30108
rect 29860 30056 29912 30108
rect 3180 29988 3232 30040
rect 4652 30031 4704 30040
rect 4652 29997 4661 30031
rect 4661 29997 4695 30031
rect 4695 29997 4704 30031
rect 4652 29988 4704 29997
rect 5388 29988 5440 30040
rect 6860 29988 6912 30040
rect 11000 30031 11052 30040
rect 11000 29997 11009 30031
rect 11009 29997 11043 30031
rect 11043 29997 11052 30031
rect 11000 29988 11052 29997
rect 12288 29988 12340 30040
rect 16152 30031 16204 30040
rect 16152 29997 16161 30031
rect 16161 29997 16195 30031
rect 16195 29997 16204 30031
rect 16152 29988 16204 29997
rect 16428 30031 16480 30040
rect 16428 29997 16437 30031
rect 16437 29997 16471 30031
rect 16471 29997 16480 30031
rect 16428 29988 16480 29997
rect 18268 29988 18320 30040
rect 23604 29988 23656 30040
rect 25996 30031 26048 30040
rect 25996 29997 26005 30031
rect 26005 29997 26039 30031
rect 26039 29997 26048 30031
rect 25996 29988 26048 29997
rect 27652 29988 27704 30040
rect 29400 29988 29452 30040
rect 1156 29920 1208 29972
rect 13024 29920 13076 29972
rect 1248 29895 1300 29904
rect 1248 29861 1257 29895
rect 1257 29861 1291 29895
rect 1291 29861 1300 29895
rect 1248 29852 1300 29861
rect 4652 29852 4704 29904
rect 13208 29895 13260 29904
rect 13208 29861 13217 29895
rect 13217 29861 13251 29895
rect 13251 29861 13260 29895
rect 13208 29852 13260 29861
rect 16244 29852 16296 29904
rect 23420 29920 23472 29972
rect 20660 29895 20712 29904
rect 20660 29861 20669 29895
rect 20669 29861 20703 29895
rect 20703 29861 20712 29895
rect 20660 29852 20712 29861
rect 23788 29852 23840 29904
rect 3510 29750 3562 29802
rect 3574 29750 3626 29802
rect 3638 29750 3690 29802
rect 3702 29750 3754 29802
rect 3766 29750 3818 29802
rect 2352 29648 2404 29700
rect 3180 29691 3232 29700
rect 3180 29657 3189 29691
rect 3189 29657 3223 29691
rect 3223 29657 3232 29691
rect 3180 29648 3232 29657
rect 3364 29691 3416 29700
rect 3364 29657 3373 29691
rect 3373 29657 3407 29691
rect 3407 29657 3416 29691
rect 3364 29648 3416 29657
rect 5020 29691 5072 29700
rect 5020 29657 5029 29691
rect 5029 29657 5063 29691
rect 5063 29657 5072 29691
rect 5020 29648 5072 29657
rect 7688 29691 7740 29700
rect 7688 29657 7697 29691
rect 7697 29657 7731 29691
rect 7731 29657 7740 29691
rect 7688 29648 7740 29657
rect 8976 29648 9028 29700
rect 10356 29648 10408 29700
rect 5388 29580 5440 29632
rect 5480 29580 5532 29632
rect 16244 29648 16296 29700
rect 16428 29648 16480 29700
rect 19004 29691 19056 29700
rect 1248 29512 1300 29564
rect 4560 29512 4612 29564
rect 10264 29555 10316 29564
rect 10264 29521 10273 29555
rect 10273 29521 10307 29555
rect 10307 29521 10316 29555
rect 10264 29512 10316 29521
rect 10908 29512 10960 29564
rect 12564 29555 12616 29564
rect 12564 29521 12573 29555
rect 12573 29521 12607 29555
rect 12607 29521 12616 29555
rect 12564 29512 12616 29521
rect 13668 29512 13720 29564
rect 15508 29512 15560 29564
rect 19004 29657 19013 29691
rect 19013 29657 19047 29691
rect 19047 29657 19056 29691
rect 19004 29648 19056 29657
rect 20476 29691 20528 29700
rect 20476 29657 20485 29691
rect 20485 29657 20519 29691
rect 20519 29657 20528 29691
rect 20476 29648 20528 29657
rect 23052 29691 23104 29700
rect 23052 29657 23061 29691
rect 23061 29657 23095 29691
rect 23095 29657 23104 29691
rect 23052 29648 23104 29657
rect 23236 29648 23288 29700
rect 23604 29691 23656 29700
rect 23604 29657 23613 29691
rect 23613 29657 23647 29691
rect 23647 29657 23656 29691
rect 23604 29648 23656 29657
rect 24156 29648 24208 29700
rect 26916 29691 26968 29700
rect 26916 29657 26925 29691
rect 26925 29657 26959 29691
rect 26959 29657 26968 29691
rect 26916 29648 26968 29657
rect 27836 29691 27888 29700
rect 27836 29657 27845 29691
rect 27845 29657 27879 29691
rect 27879 29657 27888 29691
rect 27836 29648 27888 29657
rect 2352 29444 2404 29496
rect 4100 29487 4152 29496
rect 4100 29453 4109 29487
rect 4109 29453 4143 29487
rect 4143 29453 4152 29487
rect 4100 29444 4152 29453
rect 6216 29444 6268 29496
rect 1156 29376 1208 29428
rect 2996 29385 3005 29406
rect 3005 29385 3039 29406
rect 3039 29385 3048 29406
rect 2996 29354 3048 29385
rect 3272 29308 3324 29360
rect 5296 29376 5348 29428
rect 7320 29444 7372 29496
rect 8976 29444 9028 29496
rect 9988 29487 10040 29496
rect 9988 29453 9997 29487
rect 9997 29453 10031 29487
rect 10031 29453 10040 29487
rect 9988 29444 10040 29453
rect 11828 29444 11880 29496
rect 12288 29487 12340 29496
rect 12288 29453 12297 29487
rect 12297 29453 12331 29487
rect 12331 29453 12340 29487
rect 12288 29444 12340 29453
rect 13024 29487 13076 29496
rect 8792 29376 8844 29428
rect 9068 29419 9120 29428
rect 9068 29385 9077 29419
rect 9077 29385 9111 29419
rect 9111 29385 9120 29419
rect 9068 29376 9120 29385
rect 10356 29376 10408 29428
rect 13024 29453 13033 29487
rect 13033 29453 13067 29487
rect 13067 29453 13076 29487
rect 13024 29444 13076 29453
rect 15968 29487 16020 29496
rect 15968 29453 15977 29487
rect 15977 29453 16011 29487
rect 16011 29453 16020 29487
rect 15968 29444 16020 29453
rect 16796 29444 16848 29496
rect 18268 29580 18320 29632
rect 17624 29512 17676 29564
rect 17900 29487 17952 29496
rect 17900 29453 17909 29487
rect 17909 29453 17943 29487
rect 17943 29453 17952 29487
rect 17900 29444 17952 29453
rect 24524 29512 24576 29564
rect 26456 29512 26508 29564
rect 18268 29444 18320 29496
rect 19556 29487 19608 29496
rect 19556 29453 19565 29487
rect 19565 29453 19599 29487
rect 19599 29453 19608 29487
rect 19556 29444 19608 29453
rect 20660 29444 20712 29496
rect 24156 29487 24208 29496
rect 24156 29453 24165 29487
rect 24165 29453 24199 29487
rect 24199 29453 24208 29487
rect 24156 29444 24208 29453
rect 28848 29512 28900 29564
rect 27836 29444 27888 29496
rect 13300 29419 13352 29428
rect 13300 29385 13309 29419
rect 13309 29385 13343 29419
rect 13343 29385 13352 29419
rect 13300 29376 13352 29385
rect 15048 29419 15100 29428
rect 4192 29308 4244 29360
rect 4560 29308 4612 29360
rect 4652 29308 4704 29360
rect 6308 29308 6360 29360
rect 9160 29351 9212 29360
rect 9160 29317 9169 29351
rect 9169 29317 9203 29351
rect 9203 29317 9212 29351
rect 9160 29308 9212 29317
rect 13116 29308 13168 29360
rect 13208 29308 13260 29360
rect 15048 29385 15057 29419
rect 15057 29385 15091 29419
rect 15091 29385 15100 29419
rect 15048 29376 15100 29385
rect 15416 29376 15468 29428
rect 17624 29376 17676 29428
rect 21120 29419 21172 29428
rect 16152 29308 16204 29360
rect 17348 29308 17400 29360
rect 18360 29308 18412 29360
rect 21120 29385 21129 29419
rect 21129 29385 21163 29419
rect 21163 29385 21172 29419
rect 21120 29376 21172 29385
rect 23880 29376 23932 29428
rect 24524 29376 24576 29428
rect 24892 29376 24944 29428
rect 26088 29376 26140 29428
rect 26916 29376 26968 29428
rect 27652 29376 27704 29428
rect 28204 29419 28256 29428
rect 28204 29385 28213 29419
rect 28213 29385 28247 29419
rect 28247 29385 28256 29419
rect 28204 29376 28256 29385
rect 29400 29376 29452 29428
rect 20108 29308 20160 29360
rect 23696 29308 23748 29360
rect 25996 29308 26048 29360
rect 27744 29308 27796 29360
rect 28480 29308 28532 29360
rect 18870 29206 18922 29258
rect 18934 29206 18986 29258
rect 18998 29206 19050 29258
rect 19062 29206 19114 29258
rect 19126 29206 19178 29258
rect 2352 29104 2404 29156
rect 4100 29104 4152 29156
rect 4468 29104 4520 29156
rect 5296 29104 5348 29156
rect 16888 29104 16940 29156
rect 13300 29036 13352 29088
rect 2996 28968 3048 29020
rect 4008 28968 4060 29020
rect 4284 28968 4336 29020
rect 5664 29011 5716 29020
rect 5664 28977 5673 29011
rect 5673 28977 5707 29011
rect 5707 28977 5716 29011
rect 5664 28968 5716 28977
rect 6860 29011 6912 29020
rect 6860 28977 6869 29011
rect 6869 28977 6903 29011
rect 6903 28977 6912 29011
rect 6860 28968 6912 28977
rect 8976 29011 9028 29020
rect 8976 28977 8985 29011
rect 8985 28977 9019 29011
rect 9019 28977 9028 29011
rect 8976 28968 9028 28977
rect 9068 28968 9120 29020
rect 11000 28968 11052 29020
rect 11828 29011 11880 29020
rect 11828 28977 11837 29011
rect 11837 28977 11871 29011
rect 11871 28977 11880 29011
rect 11828 28968 11880 28977
rect 13668 28968 13720 29020
rect 4928 28943 4980 28952
rect 4928 28909 4937 28943
rect 4937 28909 4971 28943
rect 4971 28909 4980 28943
rect 4928 28900 4980 28909
rect 5572 28943 5624 28952
rect 5572 28909 5581 28943
rect 5581 28909 5615 28943
rect 5615 28909 5624 28943
rect 5572 28900 5624 28909
rect 11920 28900 11972 28952
rect 13300 28943 13352 28952
rect 13300 28909 13309 28943
rect 13309 28909 13343 28943
rect 13343 28909 13352 28943
rect 13300 28900 13352 28909
rect 15232 29036 15284 29088
rect 15324 29011 15376 29020
rect 15324 28977 15333 29011
rect 15333 28977 15367 29011
rect 15367 28977 15376 29011
rect 15324 28968 15376 28977
rect 14588 28943 14640 28952
rect 14588 28909 14597 28943
rect 14597 28909 14631 28943
rect 14631 28909 14640 28943
rect 14588 28900 14640 28909
rect 14680 28900 14732 28952
rect 15508 28968 15560 29020
rect 16152 28968 16204 29020
rect 17900 29104 17952 29156
rect 24156 29147 24208 29156
rect 24156 29113 24165 29147
rect 24165 29113 24199 29147
rect 24199 29113 24208 29147
rect 24156 29104 24208 29113
rect 24892 29104 24944 29156
rect 29400 29147 29452 29156
rect 29400 29113 29409 29147
rect 29409 29113 29443 29147
rect 29443 29113 29452 29147
rect 29400 29104 29452 29113
rect 29952 29147 30004 29156
rect 29952 29113 29961 29147
rect 29961 29113 29995 29147
rect 29995 29113 30004 29147
rect 29952 29104 30004 29113
rect 17624 29036 17676 29088
rect 23420 29036 23472 29088
rect 27652 29036 27704 29088
rect 5296 28875 5348 28884
rect 5296 28841 5305 28875
rect 5305 28841 5339 28875
rect 5339 28841 5348 28875
rect 5296 28832 5348 28841
rect 1892 28807 1944 28816
rect 1892 28773 1901 28807
rect 1901 28773 1935 28807
rect 1935 28773 1944 28807
rect 1892 28764 1944 28773
rect 2076 28807 2128 28816
rect 2076 28773 2085 28807
rect 2085 28773 2119 28807
rect 2119 28773 2128 28807
rect 2076 28764 2128 28773
rect 3180 28764 3232 28816
rect 5020 28764 5072 28816
rect 7320 28832 7372 28884
rect 9528 28832 9580 28884
rect 15048 28832 15100 28884
rect 16980 28875 17032 28884
rect 16980 28841 16989 28875
rect 16989 28841 17023 28875
rect 17023 28841 17032 28875
rect 16980 28832 17032 28841
rect 17164 28832 17216 28884
rect 18728 28968 18780 29020
rect 20108 28968 20160 29020
rect 21120 28968 21172 29020
rect 23512 29011 23564 29020
rect 23512 28977 23521 29011
rect 23521 28977 23555 29011
rect 23555 28977 23564 29011
rect 23512 28968 23564 28977
rect 26916 29011 26968 29020
rect 26916 28977 26925 29011
rect 26925 28977 26959 29011
rect 26959 28977 26968 29011
rect 26916 28968 26968 28977
rect 29768 29011 29820 29020
rect 29768 28977 29777 29011
rect 29777 28977 29811 29011
rect 29811 28977 29820 29011
rect 29768 28968 29820 28977
rect 17532 28900 17584 28952
rect 20292 28900 20344 28952
rect 24616 28900 24668 28952
rect 27192 28943 27244 28952
rect 27192 28909 27201 28943
rect 27201 28909 27235 28943
rect 27235 28909 27244 28943
rect 27192 28900 27244 28909
rect 27284 28900 27336 28952
rect 6216 28807 6268 28816
rect 6216 28773 6225 28807
rect 6225 28773 6259 28807
rect 6259 28773 6268 28807
rect 6216 28764 6268 28773
rect 6952 28807 7004 28816
rect 6952 28773 6961 28807
rect 6961 28773 6995 28807
rect 6995 28773 7004 28807
rect 6952 28764 7004 28773
rect 8884 28764 8936 28816
rect 10448 28807 10500 28816
rect 10448 28773 10457 28807
rect 10457 28773 10491 28807
rect 10491 28773 10500 28807
rect 10448 28764 10500 28773
rect 18084 28764 18136 28816
rect 19280 28764 19332 28816
rect 26180 28764 26232 28816
rect 29860 28764 29912 28816
rect 3510 28662 3562 28714
rect 3574 28662 3626 28714
rect 3638 28662 3690 28714
rect 3702 28662 3754 28714
rect 3766 28662 3818 28714
rect 1156 28560 1208 28612
rect 4284 28603 4336 28612
rect 4284 28569 4293 28603
rect 4293 28569 4327 28603
rect 4327 28569 4336 28603
rect 4284 28560 4336 28569
rect 5296 28603 5348 28612
rect 5296 28569 5305 28603
rect 5305 28569 5339 28603
rect 5339 28569 5348 28603
rect 5296 28560 5348 28569
rect 5664 28603 5716 28612
rect 5664 28569 5673 28603
rect 5673 28569 5707 28603
rect 5707 28569 5716 28603
rect 5664 28560 5716 28569
rect 6216 28560 6268 28612
rect 6860 28603 6912 28612
rect 6860 28569 6869 28603
rect 6869 28569 6903 28603
rect 6903 28569 6912 28603
rect 6860 28560 6912 28569
rect 8976 28560 9028 28612
rect 10080 28560 10132 28612
rect 5572 28492 5624 28544
rect 9160 28492 9212 28544
rect 11000 28492 11052 28544
rect 11828 28492 11880 28544
rect 4744 28424 4796 28476
rect 4836 28424 4888 28476
rect 7688 28424 7740 28476
rect 9528 28424 9580 28476
rect 1892 28399 1944 28408
rect 1892 28365 1901 28399
rect 1901 28365 1935 28399
rect 1935 28365 1944 28399
rect 1892 28356 1944 28365
rect 2076 28356 2128 28408
rect 2260 28356 2312 28408
rect 3180 28356 3232 28408
rect 4192 28356 4244 28408
rect 5020 28399 5072 28408
rect 5020 28365 5029 28399
rect 5029 28365 5063 28399
rect 5063 28365 5072 28399
rect 5020 28356 5072 28365
rect 5664 28356 5716 28408
rect 6952 28356 7004 28408
rect 7596 28399 7648 28408
rect 7596 28365 7605 28399
rect 7605 28365 7639 28399
rect 7639 28365 7648 28399
rect 7596 28356 7648 28365
rect 9068 28399 9120 28408
rect 9068 28365 9077 28399
rect 9077 28365 9111 28399
rect 9111 28365 9120 28399
rect 9068 28356 9120 28365
rect 10448 28399 10500 28408
rect 10448 28365 10457 28399
rect 10457 28365 10491 28399
rect 10491 28365 10500 28399
rect 10448 28356 10500 28365
rect 13300 28560 13352 28612
rect 13668 28603 13720 28612
rect 13668 28569 13677 28603
rect 13677 28569 13711 28603
rect 13711 28569 13720 28603
rect 13668 28560 13720 28569
rect 14588 28560 14640 28612
rect 15416 28603 15468 28612
rect 15416 28569 15425 28603
rect 15425 28569 15459 28603
rect 15459 28569 15468 28603
rect 15416 28560 15468 28569
rect 16980 28603 17032 28612
rect 16980 28569 16989 28603
rect 16989 28569 17023 28603
rect 17023 28569 17032 28603
rect 16980 28560 17032 28569
rect 17164 28535 17216 28544
rect 17164 28501 17173 28535
rect 17173 28501 17207 28535
rect 17207 28501 17216 28535
rect 17164 28492 17216 28501
rect 17624 28535 17676 28544
rect 17624 28501 17633 28535
rect 17633 28501 17667 28535
rect 17667 28501 17676 28535
rect 17624 28492 17676 28501
rect 13208 28467 13260 28476
rect 13208 28433 13217 28467
rect 13217 28433 13251 28467
rect 13251 28433 13260 28467
rect 13208 28424 13260 28433
rect 16152 28467 16204 28476
rect 16152 28433 16161 28467
rect 16161 28433 16195 28467
rect 16195 28433 16204 28467
rect 16152 28424 16204 28433
rect 17532 28424 17584 28476
rect 23512 28560 23564 28612
rect 24524 28603 24576 28612
rect 24524 28569 24533 28603
rect 24533 28569 24567 28603
rect 24567 28569 24576 28603
rect 27192 28603 27244 28612
rect 24524 28560 24576 28569
rect 24616 28492 24668 28544
rect 18728 28424 18780 28476
rect 21856 28467 21908 28476
rect 21856 28433 21865 28467
rect 21865 28433 21899 28467
rect 21899 28433 21908 28467
rect 21856 28424 21908 28433
rect 13116 28356 13168 28408
rect 15048 28356 15100 28408
rect 1340 28263 1392 28272
rect 1340 28229 1349 28263
rect 1349 28229 1383 28263
rect 1383 28229 1392 28263
rect 1340 28220 1392 28229
rect 3456 28263 3508 28272
rect 3456 28229 3465 28263
rect 3465 28229 3499 28263
rect 3499 28229 3508 28263
rect 3456 28220 3508 28229
rect 4192 28220 4244 28272
rect 5756 28220 5808 28272
rect 9436 28288 9488 28340
rect 15416 28288 15468 28340
rect 15968 28288 16020 28340
rect 7688 28263 7740 28272
rect 7688 28229 7697 28263
rect 7697 28229 7731 28263
rect 7731 28229 7740 28263
rect 7688 28220 7740 28229
rect 10540 28263 10592 28272
rect 10540 28229 10549 28263
rect 10549 28229 10583 28263
rect 10583 28229 10592 28263
rect 10540 28220 10592 28229
rect 11000 28263 11052 28272
rect 11000 28229 11009 28263
rect 11009 28229 11043 28263
rect 11043 28229 11052 28263
rect 11000 28220 11052 28229
rect 11276 28220 11328 28272
rect 11920 28220 11972 28272
rect 14680 28263 14732 28272
rect 14680 28229 14689 28263
rect 14689 28229 14723 28263
rect 14723 28229 14732 28263
rect 14680 28220 14732 28229
rect 15232 28263 15284 28272
rect 15232 28229 15241 28263
rect 15241 28229 15275 28263
rect 15275 28229 15284 28263
rect 15232 28220 15284 28229
rect 17348 28356 17400 28408
rect 18084 28399 18136 28408
rect 18084 28365 18093 28399
rect 18093 28365 18127 28399
rect 18127 28365 18136 28399
rect 18084 28356 18136 28365
rect 23052 28424 23104 28476
rect 27192 28569 27201 28603
rect 27201 28569 27235 28603
rect 27235 28569 27244 28603
rect 27192 28560 27244 28569
rect 27652 28560 27704 28612
rect 28204 28603 28256 28612
rect 28204 28569 28213 28603
rect 28213 28569 28247 28603
rect 28247 28569 28256 28603
rect 29952 28603 30004 28612
rect 28204 28560 28256 28569
rect 26916 28492 26968 28544
rect 26180 28424 26232 28476
rect 28112 28424 28164 28476
rect 29952 28569 29961 28603
rect 29961 28569 29995 28603
rect 29995 28569 30004 28603
rect 29952 28560 30004 28569
rect 19372 28288 19424 28340
rect 20108 28288 20160 28340
rect 23696 28356 23748 28408
rect 24984 28399 25036 28408
rect 22500 28288 22552 28340
rect 23052 28288 23104 28340
rect 24984 28365 24993 28399
rect 24993 28365 25027 28399
rect 25027 28365 25036 28399
rect 24984 28356 25036 28365
rect 28020 28399 28072 28408
rect 28020 28365 28029 28399
rect 28029 28365 28063 28399
rect 28063 28365 28072 28399
rect 28020 28356 28072 28365
rect 26088 28288 26140 28340
rect 29584 28399 29636 28408
rect 29584 28365 29593 28399
rect 29593 28365 29627 28399
rect 29627 28365 29636 28399
rect 29584 28356 29636 28365
rect 16612 28220 16664 28272
rect 17992 28263 18044 28272
rect 17992 28229 18001 28263
rect 18001 28229 18035 28263
rect 18035 28229 18044 28263
rect 17992 28220 18044 28229
rect 20292 28220 20344 28272
rect 27284 28220 27336 28272
rect 28480 28220 28532 28272
rect 29032 28220 29084 28272
rect 29768 28263 29820 28272
rect 29768 28229 29777 28263
rect 29777 28229 29811 28263
rect 29811 28229 29820 28263
rect 29768 28220 29820 28229
rect 18870 28118 18922 28170
rect 18934 28118 18986 28170
rect 18998 28118 19050 28170
rect 19062 28118 19114 28170
rect 19126 28118 19178 28170
rect 3088 28016 3140 28068
rect 3364 28016 3416 28068
rect 4284 28059 4336 28068
rect 4284 28025 4293 28059
rect 4293 28025 4327 28059
rect 4327 28025 4336 28059
rect 4284 28016 4336 28025
rect 4928 28016 4980 28068
rect 7688 28016 7740 28068
rect 9068 28016 9120 28068
rect 9252 28059 9304 28068
rect 9252 28025 9261 28059
rect 9261 28025 9295 28059
rect 9295 28025 9304 28059
rect 9252 28016 9304 28025
rect 10540 28016 10592 28068
rect 16152 28016 16204 28068
rect 17992 28016 18044 28068
rect 18728 28016 18780 28068
rect 19280 28016 19332 28068
rect 23052 28059 23104 28068
rect 23052 28025 23061 28059
rect 23061 28025 23095 28059
rect 23095 28025 23104 28059
rect 23052 28016 23104 28025
rect 24984 28059 25036 28068
rect 24984 28025 24993 28059
rect 24993 28025 25027 28059
rect 25027 28025 25036 28059
rect 24984 28016 25036 28025
rect 1340 27948 1392 28000
rect 1984 27880 2036 27932
rect 4100 27948 4152 28000
rect 8792 27948 8844 28000
rect 11276 27948 11328 28000
rect 14956 27948 15008 28000
rect 17532 27948 17584 28000
rect 19372 27948 19424 28000
rect 20936 27948 20988 28000
rect 24616 27991 24668 28000
rect 24616 27957 24625 27991
rect 24625 27957 24659 27991
rect 24659 27957 24668 27991
rect 27836 28016 27888 28068
rect 27192 27991 27244 28000
rect 24616 27948 24668 27957
rect 27192 27957 27201 27991
rect 27201 27957 27235 27991
rect 27235 27957 27244 27991
rect 27192 27948 27244 27957
rect 2168 27880 2220 27932
rect 3364 27923 3416 27932
rect 3364 27889 3373 27923
rect 3373 27889 3407 27923
rect 3407 27889 3416 27923
rect 3364 27880 3416 27889
rect 3456 27880 3508 27932
rect 4008 27880 4060 27932
rect 5664 27923 5716 27932
rect 5664 27889 5673 27923
rect 5673 27889 5707 27923
rect 5707 27889 5716 27923
rect 5664 27880 5716 27889
rect 9344 27880 9396 27932
rect 9436 27923 9488 27932
rect 9436 27889 9445 27923
rect 9445 27889 9479 27923
rect 9479 27889 9488 27923
rect 9436 27880 9488 27889
rect 10356 27880 10408 27932
rect 15968 27880 16020 27932
rect 16796 27923 16848 27932
rect 16796 27889 16805 27923
rect 16805 27889 16839 27923
rect 16839 27889 16848 27923
rect 16796 27880 16848 27889
rect 20200 27923 20252 27932
rect 20200 27889 20209 27923
rect 20209 27889 20243 27923
rect 20243 27889 20252 27923
rect 20200 27880 20252 27889
rect 22408 27923 22460 27932
rect 22408 27889 22417 27923
rect 22417 27889 22451 27923
rect 22451 27889 22460 27923
rect 22408 27880 22460 27889
rect 22500 27880 22552 27932
rect 24340 27923 24392 27932
rect 24340 27889 24349 27923
rect 24349 27889 24383 27923
rect 24383 27889 24392 27923
rect 24340 27880 24392 27889
rect 27284 27880 27336 27932
rect 28112 27880 28164 27932
rect 29584 28016 29636 28068
rect 29676 27923 29728 27932
rect 29676 27889 29685 27923
rect 29685 27889 29719 27923
rect 29719 27889 29728 27923
rect 29676 27880 29728 27889
rect 2444 27855 2496 27864
rect 2444 27821 2453 27855
rect 2453 27821 2487 27855
rect 2487 27821 2496 27855
rect 2444 27812 2496 27821
rect 4836 27855 4888 27864
rect 4836 27821 4845 27855
rect 4845 27821 4879 27855
rect 4879 27821 4888 27855
rect 4836 27812 4888 27821
rect 5020 27812 5072 27864
rect 5756 27812 5808 27864
rect 5848 27855 5900 27864
rect 5848 27821 5857 27855
rect 5857 27821 5891 27855
rect 5891 27821 5900 27855
rect 10816 27855 10868 27864
rect 5848 27812 5900 27821
rect 10816 27821 10825 27855
rect 10825 27821 10859 27855
rect 10859 27821 10868 27855
rect 10816 27812 10868 27821
rect 12656 27812 12708 27864
rect 22224 27812 22276 27864
rect 27560 27812 27612 27864
rect 30044 27855 30096 27864
rect 30044 27821 30053 27855
rect 30053 27821 30087 27855
rect 30087 27821 30096 27855
rect 30044 27812 30096 27821
rect 8884 27744 8936 27796
rect 14864 27744 14916 27796
rect 23512 27744 23564 27796
rect 7872 27676 7924 27728
rect 15416 27719 15468 27728
rect 15416 27685 15425 27719
rect 15425 27685 15459 27719
rect 15459 27685 15468 27719
rect 15416 27676 15468 27685
rect 16612 27719 16664 27728
rect 16612 27685 16621 27719
rect 16621 27685 16655 27719
rect 16655 27685 16664 27719
rect 16612 27676 16664 27685
rect 3510 27574 3562 27626
rect 3574 27574 3626 27626
rect 3638 27574 3690 27626
rect 3702 27574 3754 27626
rect 3766 27574 3818 27626
rect 2168 27515 2220 27524
rect 2168 27481 2177 27515
rect 2177 27481 2211 27515
rect 2211 27481 2220 27515
rect 2168 27472 2220 27481
rect 4100 27472 4152 27524
rect 4836 27472 4888 27524
rect 6032 27472 6084 27524
rect 9436 27515 9488 27524
rect 2444 27404 2496 27456
rect 3272 27404 3324 27456
rect 5020 27447 5072 27456
rect 5020 27413 5029 27447
rect 5029 27413 5063 27447
rect 5063 27413 5072 27447
rect 5020 27404 5072 27413
rect 5664 27404 5716 27456
rect 6860 27404 6912 27456
rect 7596 27447 7648 27456
rect 7596 27413 7605 27447
rect 7605 27413 7639 27447
rect 7639 27413 7648 27447
rect 7596 27404 7648 27413
rect 1432 27336 1484 27388
rect 2076 27336 2128 27388
rect 2720 27336 2772 27388
rect 5848 27336 5900 27388
rect 2904 27311 2956 27320
rect 2904 27277 2913 27311
rect 2913 27277 2947 27311
rect 2947 27277 2956 27311
rect 2904 27268 2956 27277
rect 3088 27311 3140 27320
rect 3088 27277 3097 27311
rect 3097 27277 3131 27311
rect 3131 27277 3140 27311
rect 3088 27268 3140 27277
rect 7872 27311 7924 27320
rect 7872 27277 7881 27311
rect 7881 27277 7915 27311
rect 7915 27277 7924 27311
rect 7872 27268 7924 27277
rect 9436 27481 9445 27515
rect 9445 27481 9479 27515
rect 9479 27481 9488 27515
rect 9436 27472 9488 27481
rect 10356 27515 10408 27524
rect 10356 27481 10365 27515
rect 10365 27481 10399 27515
rect 10399 27481 10408 27515
rect 10356 27472 10408 27481
rect 10816 27515 10868 27524
rect 10816 27481 10825 27515
rect 10825 27481 10859 27515
rect 10859 27481 10868 27515
rect 10816 27472 10868 27481
rect 11276 27472 11328 27524
rect 15416 27472 15468 27524
rect 15968 27515 16020 27524
rect 15968 27481 15977 27515
rect 15977 27481 16011 27515
rect 16011 27481 16020 27515
rect 15968 27472 16020 27481
rect 16428 27472 16480 27524
rect 17164 27472 17216 27524
rect 20936 27515 20988 27524
rect 20936 27481 20945 27515
rect 20945 27481 20979 27515
rect 20979 27481 20988 27515
rect 20936 27472 20988 27481
rect 24340 27472 24392 27524
rect 27192 27515 27244 27524
rect 27192 27481 27201 27515
rect 27201 27481 27235 27515
rect 27235 27481 27244 27515
rect 27192 27472 27244 27481
rect 27560 27515 27612 27524
rect 27560 27481 27569 27515
rect 27569 27481 27603 27515
rect 27603 27481 27612 27515
rect 27560 27472 27612 27481
rect 30044 27472 30096 27524
rect 14956 27447 15008 27456
rect 14956 27413 14965 27447
rect 14965 27413 14999 27447
rect 14999 27413 15008 27447
rect 14956 27404 15008 27413
rect 15048 27404 15100 27456
rect 9344 27379 9396 27388
rect 9344 27345 9353 27379
rect 9353 27345 9387 27379
rect 9387 27345 9396 27379
rect 10632 27379 10684 27388
rect 9344 27336 9396 27345
rect 10632 27345 10641 27379
rect 10641 27345 10675 27379
rect 10675 27345 10684 27379
rect 10632 27336 10684 27345
rect 12656 27379 12708 27388
rect 12656 27345 12665 27379
rect 12665 27345 12699 27379
rect 12699 27345 12708 27379
rect 12656 27336 12708 27345
rect 8700 27311 8752 27320
rect 8700 27277 8709 27311
rect 8709 27277 8743 27311
rect 8743 27277 8752 27311
rect 8700 27268 8752 27277
rect 8884 27311 8936 27320
rect 8884 27277 8893 27311
rect 8893 27277 8927 27311
rect 8927 27277 8936 27311
rect 8884 27268 8936 27277
rect 9252 27268 9304 27320
rect 11000 27268 11052 27320
rect 12564 27311 12616 27320
rect 12564 27277 12573 27311
rect 12573 27277 12607 27311
rect 12607 27277 12616 27311
rect 12564 27268 12616 27277
rect 16796 27404 16848 27456
rect 28112 27404 28164 27456
rect 16888 27336 16940 27388
rect 20200 27336 20252 27388
rect 22960 27379 23012 27388
rect 22960 27345 22969 27379
rect 22969 27345 23003 27379
rect 23003 27345 23012 27379
rect 22960 27336 23012 27345
rect 1984 27243 2036 27252
rect 1984 27209 1993 27243
rect 1993 27209 2027 27243
rect 2027 27209 2036 27243
rect 1984 27200 2036 27209
rect 3272 27200 3324 27252
rect 3364 27200 3416 27252
rect 9988 27200 10040 27252
rect 15968 27200 16020 27252
rect 21120 27268 21172 27320
rect 1156 27132 1208 27184
rect 1524 27132 1576 27184
rect 4008 27132 4060 27184
rect 6952 27132 7004 27184
rect 12288 27132 12340 27184
rect 14956 27132 15008 27184
rect 15232 27132 15284 27184
rect 16612 27132 16664 27184
rect 22408 27200 22460 27252
rect 23328 27200 23380 27252
rect 23696 27200 23748 27252
rect 20660 27175 20712 27184
rect 20660 27141 20669 27175
rect 20669 27141 20703 27175
rect 20703 27141 20712 27175
rect 20660 27132 20712 27141
rect 22224 27175 22276 27184
rect 22224 27141 22233 27175
rect 22233 27141 22267 27175
rect 22267 27141 22276 27175
rect 22224 27132 22276 27141
rect 24524 27132 24576 27184
rect 27284 27132 27336 27184
rect 28296 27132 28348 27184
rect 29676 27175 29728 27184
rect 29676 27141 29685 27175
rect 29685 27141 29719 27175
rect 29719 27141 29728 27175
rect 29676 27132 29728 27141
rect 18870 27030 18922 27082
rect 18934 27030 18986 27082
rect 18998 27030 19050 27082
rect 19062 27030 19114 27082
rect 19126 27030 19178 27082
rect 2720 26971 2772 26980
rect 2720 26937 2729 26971
rect 2729 26937 2763 26971
rect 2763 26937 2772 26971
rect 2720 26928 2772 26937
rect 7596 26928 7648 26980
rect 8700 26971 8752 26980
rect 8700 26937 8709 26971
rect 8709 26937 8743 26971
rect 8743 26937 8752 26971
rect 8700 26928 8752 26937
rect 10540 26928 10592 26980
rect 12564 26928 12616 26980
rect 22224 26928 22276 26980
rect 23696 26928 23748 26980
rect 24616 26928 24668 26980
rect 10816 26860 10868 26912
rect 3272 26792 3324 26844
rect 6584 26835 6636 26844
rect 6584 26801 6593 26835
rect 6593 26801 6627 26835
rect 6627 26801 6636 26835
rect 6584 26792 6636 26801
rect 9804 26835 9856 26844
rect 9804 26801 9813 26835
rect 9813 26801 9847 26835
rect 9847 26801 9856 26835
rect 9804 26792 9856 26801
rect 9988 26835 10040 26844
rect 9988 26801 9997 26835
rect 9997 26801 10031 26835
rect 10031 26801 10040 26835
rect 9988 26792 10040 26801
rect 10632 26835 10684 26844
rect 6952 26767 7004 26776
rect 6952 26733 6961 26767
rect 6961 26733 6995 26767
rect 6995 26733 7004 26767
rect 6952 26724 7004 26733
rect 9620 26724 9672 26776
rect 10632 26801 10641 26835
rect 10641 26801 10675 26835
rect 10675 26801 10684 26835
rect 10632 26792 10684 26801
rect 14864 26835 14916 26844
rect 14864 26801 14873 26835
rect 14873 26801 14907 26835
rect 14907 26801 14916 26835
rect 14864 26792 14916 26801
rect 15232 26792 15284 26844
rect 16428 26835 16480 26844
rect 16428 26801 16437 26835
rect 16437 26801 16471 26835
rect 16471 26801 16480 26835
rect 16428 26792 16480 26801
rect 26180 26860 26232 26912
rect 16612 26792 16664 26844
rect 21856 26792 21908 26844
rect 25904 26792 25956 26844
rect 28572 26835 28624 26844
rect 28572 26801 28581 26835
rect 28581 26801 28615 26835
rect 28615 26801 28624 26835
rect 28572 26792 28624 26801
rect 10356 26767 10408 26776
rect 10356 26733 10365 26767
rect 10365 26733 10399 26767
rect 10399 26733 10408 26767
rect 10356 26724 10408 26733
rect 15324 26767 15376 26776
rect 15324 26733 15333 26767
rect 15333 26733 15367 26767
rect 15367 26733 15376 26767
rect 15324 26724 15376 26733
rect 2720 26656 2772 26708
rect 6860 26699 6912 26708
rect 6860 26665 6869 26699
rect 6869 26665 6903 26699
rect 6903 26665 6912 26699
rect 6860 26656 6912 26665
rect 15140 26656 15192 26708
rect 21396 26767 21448 26776
rect 21396 26733 21405 26767
rect 21405 26733 21439 26767
rect 21439 26733 21448 26767
rect 21396 26724 21448 26733
rect 1432 26588 1484 26640
rect 3364 26588 3416 26640
rect 6768 26631 6820 26640
rect 6768 26597 6792 26631
rect 6792 26597 6820 26631
rect 6768 26588 6820 26597
rect 7228 26631 7280 26640
rect 7228 26597 7237 26631
rect 7237 26597 7271 26631
rect 7271 26597 7280 26631
rect 7228 26588 7280 26597
rect 15048 26588 15100 26640
rect 16796 26588 16848 26640
rect 28756 26631 28808 26640
rect 28756 26597 28765 26631
rect 28765 26597 28799 26631
rect 28799 26597 28808 26631
rect 28756 26588 28808 26597
rect 3510 26486 3562 26538
rect 3574 26486 3626 26538
rect 3638 26486 3690 26538
rect 3702 26486 3754 26538
rect 3766 26486 3818 26538
rect 2904 26384 2956 26436
rect 6768 26384 6820 26436
rect 9804 26384 9856 26436
rect 11828 26384 11880 26436
rect 14956 26384 15008 26436
rect 15508 26384 15560 26436
rect 16428 26427 16480 26436
rect 16428 26393 16437 26427
rect 16437 26393 16471 26427
rect 16471 26393 16480 26427
rect 16428 26384 16480 26393
rect 16612 26427 16664 26436
rect 16612 26393 16621 26427
rect 16621 26393 16655 26427
rect 16655 26393 16664 26427
rect 16612 26384 16664 26393
rect 16796 26427 16848 26436
rect 16796 26393 16805 26427
rect 16805 26393 16839 26427
rect 16839 26393 16848 26427
rect 16796 26384 16848 26393
rect 21396 26427 21448 26436
rect 21396 26393 21405 26427
rect 21405 26393 21439 26427
rect 21439 26393 21448 26427
rect 21396 26384 21448 26393
rect 6952 26359 7004 26368
rect 6952 26325 6961 26359
rect 6961 26325 6995 26359
rect 6995 26325 7004 26359
rect 6952 26316 7004 26325
rect 10816 26316 10868 26368
rect 21856 26384 21908 26436
rect 24984 26427 25036 26436
rect 24984 26393 24993 26427
rect 24993 26393 25027 26427
rect 25027 26393 25036 26427
rect 24984 26384 25036 26393
rect 26180 26384 26232 26436
rect 28572 26427 28624 26436
rect 28572 26393 28581 26427
rect 28581 26393 28615 26427
rect 28615 26393 28624 26427
rect 28572 26384 28624 26393
rect 28756 26427 28808 26436
rect 28756 26393 28765 26427
rect 28765 26393 28799 26427
rect 28799 26393 28808 26427
rect 28756 26384 28808 26393
rect 2720 26291 2772 26300
rect 2720 26257 2729 26291
rect 2729 26257 2763 26291
rect 2763 26257 2772 26291
rect 2720 26248 2772 26257
rect 6860 26248 6912 26300
rect 696 26223 748 26232
rect 696 26189 705 26223
rect 705 26189 739 26223
rect 739 26189 748 26223
rect 696 26180 748 26189
rect 788 26044 840 26096
rect 1432 26112 1484 26164
rect 6124 26223 6176 26232
rect 6124 26189 6133 26223
rect 6133 26189 6167 26223
rect 6167 26189 6176 26223
rect 6124 26180 6176 26189
rect 8700 26180 8752 26232
rect 9252 26223 9304 26232
rect 9252 26189 9261 26223
rect 9261 26189 9295 26223
rect 9295 26189 9304 26223
rect 9252 26180 9304 26189
rect 10632 26248 10684 26300
rect 3272 26044 3324 26096
rect 3456 26044 3508 26096
rect 4560 26087 4612 26096
rect 4560 26053 4569 26087
rect 4569 26053 4603 26087
rect 4603 26053 4612 26087
rect 4560 26044 4612 26053
rect 7872 26044 7924 26096
rect 8240 26087 8292 26096
rect 8240 26053 8249 26087
rect 8249 26053 8283 26087
rect 8283 26053 8292 26087
rect 10540 26180 10592 26232
rect 11828 26180 11880 26232
rect 14680 26248 14732 26300
rect 15048 26223 15100 26232
rect 10724 26112 10776 26164
rect 15048 26189 15057 26223
rect 15057 26189 15091 26223
rect 15091 26189 15100 26223
rect 15048 26180 15100 26189
rect 16428 26248 16480 26300
rect 15508 26223 15560 26232
rect 15508 26189 15517 26223
rect 15517 26189 15551 26223
rect 15551 26189 15560 26223
rect 15508 26180 15560 26189
rect 17808 26180 17860 26232
rect 20108 26180 20160 26232
rect 20200 26180 20252 26232
rect 30044 26316 30096 26368
rect 28020 26248 28072 26300
rect 15232 26112 15284 26164
rect 14680 26087 14732 26096
rect 8240 26044 8292 26053
rect 14680 26053 14689 26087
rect 14689 26053 14723 26087
rect 14723 26053 14732 26087
rect 14680 26044 14732 26053
rect 17716 26044 17768 26096
rect 20936 26112 20988 26164
rect 24248 26112 24300 26164
rect 18268 26087 18320 26096
rect 18268 26053 18277 26087
rect 18277 26053 18311 26087
rect 18311 26053 18320 26087
rect 18268 26044 18320 26053
rect 27100 26180 27152 26232
rect 29860 26180 29912 26232
rect 25904 26087 25956 26096
rect 25904 26053 25913 26087
rect 25913 26053 25947 26087
rect 25947 26053 25956 26087
rect 25904 26044 25956 26053
rect 29308 26112 29360 26164
rect 27192 26044 27244 26096
rect 29860 26044 29912 26096
rect 18870 25942 18922 25994
rect 18934 25942 18986 25994
rect 18998 25942 19050 25994
rect 19062 25942 19114 25994
rect 19126 25942 19178 25994
rect 1892 25840 1944 25892
rect 2628 25840 2680 25892
rect 8700 25883 8752 25892
rect 8700 25849 8709 25883
rect 8709 25849 8743 25883
rect 8743 25849 8752 25883
rect 8700 25840 8752 25849
rect 3088 25772 3140 25824
rect 6032 25815 6084 25824
rect 3364 25704 3416 25756
rect 6032 25781 6041 25815
rect 6041 25781 6075 25815
rect 6075 25781 6084 25815
rect 6032 25772 6084 25781
rect 6584 25772 6636 25824
rect 9988 25840 10040 25892
rect 14680 25883 14732 25892
rect 14680 25849 14689 25883
rect 14689 25849 14723 25883
rect 14723 25849 14732 25883
rect 14680 25840 14732 25849
rect 14864 25840 14916 25892
rect 15324 25883 15376 25892
rect 15324 25849 15333 25883
rect 15333 25849 15367 25883
rect 15367 25849 15376 25883
rect 15324 25840 15376 25849
rect 24892 25840 24944 25892
rect 15048 25772 15100 25824
rect 5756 25747 5808 25756
rect 5756 25713 5765 25747
rect 5765 25713 5799 25747
rect 5799 25713 5808 25747
rect 5756 25704 5808 25713
rect 7688 25704 7740 25756
rect 9804 25704 9856 25756
rect 10356 25704 10408 25756
rect 15140 25704 15192 25756
rect 16796 25704 16848 25756
rect 22500 25772 22552 25824
rect 27560 25772 27612 25824
rect 18452 25704 18504 25756
rect 20200 25747 20252 25756
rect 20200 25713 20209 25747
rect 20209 25713 20243 25747
rect 20243 25713 20252 25747
rect 20200 25704 20252 25713
rect 21396 25704 21448 25756
rect 24524 25747 24576 25756
rect 24524 25713 24533 25747
rect 24533 25713 24567 25747
rect 24567 25713 24576 25747
rect 24524 25704 24576 25713
rect 26732 25747 26784 25756
rect 26732 25713 26741 25747
rect 26741 25713 26775 25747
rect 26775 25713 26784 25747
rect 26732 25704 26784 25713
rect 27100 25704 27152 25756
rect 27836 25704 27888 25756
rect 696 25636 748 25688
rect 2720 25636 2772 25688
rect 3916 25679 3968 25688
rect 788 25543 840 25552
rect 788 25509 797 25543
rect 797 25509 831 25543
rect 831 25509 840 25543
rect 788 25500 840 25509
rect 3916 25645 3925 25679
rect 3925 25645 3959 25679
rect 3959 25645 3968 25679
rect 3916 25636 3968 25645
rect 4284 25679 4336 25688
rect 4284 25645 4293 25679
rect 4293 25645 4327 25679
rect 4327 25645 4336 25679
rect 4284 25636 4336 25645
rect 7228 25636 7280 25688
rect 12748 25636 12800 25688
rect 15508 25636 15560 25688
rect 16336 25636 16388 25688
rect 17716 25679 17768 25688
rect 17716 25645 17725 25679
rect 17725 25645 17759 25679
rect 17759 25645 17768 25679
rect 17716 25636 17768 25645
rect 18176 25636 18228 25688
rect 20384 25679 20436 25688
rect 20384 25645 20393 25679
rect 20393 25645 20427 25679
rect 20427 25645 20436 25679
rect 20384 25636 20436 25645
rect 21856 25679 21908 25688
rect 21856 25645 21865 25679
rect 21865 25645 21899 25679
rect 21899 25645 21908 25679
rect 21856 25636 21908 25645
rect 22224 25636 22276 25688
rect 23236 25636 23288 25688
rect 28572 25636 28624 25688
rect 6492 25568 6544 25620
rect 10632 25568 10684 25620
rect 15600 25568 15652 25620
rect 18268 25568 18320 25620
rect 4928 25500 4980 25552
rect 9620 25543 9672 25552
rect 9620 25509 9629 25543
rect 9629 25509 9663 25543
rect 9663 25509 9672 25543
rect 9620 25500 9672 25509
rect 13024 25500 13076 25552
rect 14680 25500 14732 25552
rect 16244 25500 16296 25552
rect 16428 25543 16480 25552
rect 16428 25509 16437 25543
rect 16437 25509 16471 25543
rect 16471 25509 16480 25543
rect 16428 25500 16480 25509
rect 17348 25500 17400 25552
rect 24432 25500 24484 25552
rect 3510 25398 3562 25450
rect 3574 25398 3626 25450
rect 3638 25398 3690 25450
rect 3702 25398 3754 25450
rect 3766 25398 3818 25450
rect 4284 25296 4336 25348
rect 4928 25339 4980 25348
rect 788 25228 840 25280
rect 3272 25271 3324 25280
rect 3272 25237 3281 25271
rect 3281 25237 3315 25271
rect 3315 25237 3324 25271
rect 4928 25305 4937 25339
rect 4937 25305 4971 25339
rect 4971 25305 4980 25339
rect 4928 25296 4980 25305
rect 6032 25296 6084 25348
rect 12564 25296 12616 25348
rect 16428 25296 16480 25348
rect 20200 25339 20252 25348
rect 20200 25305 20209 25339
rect 20209 25305 20243 25339
rect 20243 25305 20252 25339
rect 20200 25296 20252 25305
rect 21396 25296 21448 25348
rect 22224 25339 22276 25348
rect 22224 25305 22233 25339
rect 22233 25305 22267 25339
rect 22267 25305 22276 25339
rect 22224 25296 22276 25305
rect 22500 25339 22552 25348
rect 22500 25305 22509 25339
rect 22509 25305 22543 25339
rect 22543 25305 22552 25339
rect 22500 25296 22552 25305
rect 23328 25339 23380 25348
rect 23328 25305 23337 25339
rect 23337 25305 23371 25339
rect 23371 25305 23380 25339
rect 23328 25296 23380 25305
rect 24524 25296 24576 25348
rect 3272 25228 3324 25237
rect 5756 25228 5808 25280
rect 2352 25135 2404 25144
rect 2352 25101 2361 25135
rect 2361 25101 2395 25135
rect 2395 25101 2404 25135
rect 2352 25092 2404 25101
rect 2628 25135 2680 25144
rect 2628 25101 2637 25135
rect 2637 25101 2671 25135
rect 2671 25101 2680 25135
rect 2628 25092 2680 25101
rect 2720 25135 2772 25144
rect 2720 25101 2729 25135
rect 2729 25101 2763 25135
rect 2763 25101 2772 25135
rect 2720 25092 2772 25101
rect 4560 25092 4612 25144
rect 4284 25024 4336 25076
rect 3088 24956 3140 25008
rect 3824 24999 3876 25008
rect 3824 24965 3833 24999
rect 3833 24965 3867 24999
rect 3867 24965 3876 24999
rect 3824 24956 3876 24965
rect 4560 24999 4612 25008
rect 4560 24965 4569 24999
rect 4569 24965 4603 24999
rect 4603 24965 4612 24999
rect 4560 24956 4612 24965
rect 14956 25228 15008 25280
rect 16336 25271 16388 25280
rect 16336 25237 16345 25271
rect 16345 25237 16379 25271
rect 16379 25237 16388 25271
rect 16336 25228 16388 25237
rect 16796 25271 16848 25280
rect 16796 25237 16805 25271
rect 16805 25237 16839 25271
rect 16839 25237 16848 25271
rect 16796 25228 16848 25237
rect 18636 25228 18688 25280
rect 20384 25228 20436 25280
rect 5940 25092 5992 25144
rect 10448 25160 10500 25212
rect 16244 25160 16296 25212
rect 18360 25160 18412 25212
rect 21672 25160 21724 25212
rect 24892 25228 24944 25280
rect 26180 25228 26232 25280
rect 17348 25135 17400 25144
rect 6400 25067 6452 25076
rect 6400 25033 6409 25067
rect 6409 25033 6443 25067
rect 6443 25033 6452 25067
rect 6400 25024 6452 25033
rect 8240 25024 8292 25076
rect 7044 24956 7096 25008
rect 17348 25101 17357 25135
rect 17357 25101 17391 25135
rect 17391 25101 17400 25135
rect 17348 25092 17400 25101
rect 20292 25135 20344 25144
rect 20292 25101 20301 25135
rect 20301 25101 20335 25135
rect 20335 25101 20344 25135
rect 20292 25092 20344 25101
rect 20660 25092 20712 25144
rect 11460 24956 11512 25008
rect 12656 24999 12708 25008
rect 12656 24965 12665 24999
rect 12665 24965 12699 24999
rect 12699 24965 12708 24999
rect 12656 24956 12708 24965
rect 13300 24999 13352 25008
rect 13300 24965 13309 24999
rect 13309 24965 13343 24999
rect 13343 24965 13352 24999
rect 16888 25024 16940 25076
rect 18268 25024 18320 25076
rect 19372 25067 19424 25076
rect 19372 25033 19381 25067
rect 19381 25033 19415 25067
rect 19415 25033 19424 25067
rect 19372 25024 19424 25033
rect 21856 25024 21908 25076
rect 14956 24999 15008 25008
rect 13300 24956 13352 24965
rect 14956 24965 14965 24999
rect 14965 24965 14999 24999
rect 14999 24965 15008 24999
rect 14956 24956 15008 24965
rect 15600 24956 15652 25008
rect 16980 24999 17032 25008
rect 16980 24965 16989 24999
rect 16989 24965 17023 24999
rect 17023 24965 17032 24999
rect 16980 24956 17032 24965
rect 17072 24956 17124 25008
rect 17900 24956 17952 25008
rect 22592 24956 22644 25008
rect 24524 25092 24576 25144
rect 24708 25135 24760 25144
rect 24708 25101 24717 25135
rect 24717 25101 24751 25135
rect 24751 25101 24760 25135
rect 24708 25092 24760 25101
rect 26180 25092 26232 25144
rect 27100 25296 27152 25348
rect 27560 25296 27612 25348
rect 28572 25203 28624 25212
rect 28572 25169 28581 25203
rect 28581 25169 28615 25203
rect 28615 25169 28624 25203
rect 28572 25160 28624 25169
rect 26732 25092 26784 25144
rect 24432 25024 24484 25076
rect 25904 25024 25956 25076
rect 28388 25024 28440 25076
rect 29308 25024 29360 25076
rect 30596 25067 30648 25076
rect 30596 25033 30605 25067
rect 30605 25033 30639 25067
rect 30639 25033 30648 25067
rect 30596 25024 30648 25033
rect 26548 24999 26600 25008
rect 26548 24965 26557 24999
rect 26557 24965 26591 24999
rect 26591 24965 26600 24999
rect 26548 24956 26600 24965
rect 27836 24999 27888 25008
rect 27836 24965 27845 24999
rect 27845 24965 27879 24999
rect 27879 24965 27888 24999
rect 27836 24956 27888 24965
rect 28480 24956 28532 25008
rect 18870 24854 18922 24906
rect 18934 24854 18986 24906
rect 18998 24854 19050 24906
rect 19062 24854 19114 24906
rect 19126 24854 19178 24906
rect 1892 24752 1944 24804
rect 2352 24752 2404 24804
rect 3364 24795 3416 24804
rect 3364 24761 3373 24795
rect 3373 24761 3407 24795
rect 3407 24761 3416 24795
rect 3364 24752 3416 24761
rect 18176 24795 18228 24804
rect 18176 24761 18185 24795
rect 18185 24761 18219 24795
rect 18219 24761 18228 24795
rect 18176 24752 18228 24761
rect 24708 24752 24760 24804
rect 29308 24752 29360 24804
rect 1156 24684 1208 24736
rect 3916 24548 3968 24600
rect 4284 24548 4336 24600
rect 4652 24659 4704 24668
rect 4652 24625 4661 24659
rect 4661 24625 4695 24659
rect 4695 24625 4704 24659
rect 4652 24616 4704 24625
rect 5388 24616 5440 24668
rect 5848 24616 5900 24668
rect 7780 24684 7832 24736
rect 16980 24684 17032 24736
rect 21672 24684 21724 24736
rect 26180 24727 26232 24736
rect 26180 24693 26189 24727
rect 26189 24693 26223 24727
rect 26223 24693 26232 24727
rect 26180 24684 26232 24693
rect 9252 24659 9304 24668
rect 9252 24625 9261 24659
rect 9261 24625 9295 24659
rect 9295 24625 9304 24659
rect 9252 24616 9304 24625
rect 15600 24659 15652 24668
rect 15600 24625 15609 24659
rect 15609 24625 15643 24659
rect 15643 24625 15652 24659
rect 15600 24616 15652 24625
rect 15784 24659 15836 24668
rect 15784 24625 15793 24659
rect 15793 24625 15827 24659
rect 15827 24625 15836 24659
rect 15784 24616 15836 24625
rect 17900 24659 17952 24668
rect 17900 24625 17909 24659
rect 17909 24625 17943 24659
rect 17943 24625 17952 24659
rect 17900 24616 17952 24625
rect 18728 24616 18780 24668
rect 19372 24616 19424 24668
rect 20936 24659 20988 24668
rect 20936 24625 20945 24659
rect 20945 24625 20979 24659
rect 20979 24625 20988 24659
rect 20936 24616 20988 24625
rect 25904 24659 25956 24668
rect 25904 24625 25913 24659
rect 25913 24625 25947 24659
rect 25947 24625 25956 24659
rect 25904 24616 25956 24625
rect 26272 24616 26324 24668
rect 27376 24616 27428 24668
rect 27560 24659 27612 24668
rect 27560 24625 27569 24659
rect 27569 24625 27603 24659
rect 27603 24625 27612 24659
rect 27560 24616 27612 24625
rect 28204 24659 28256 24668
rect 28204 24625 28213 24659
rect 28213 24625 28247 24659
rect 28247 24625 28256 24659
rect 28204 24616 28256 24625
rect 29860 24616 29912 24668
rect 4560 24548 4612 24600
rect 6216 24548 6268 24600
rect 7688 24548 7740 24600
rect 16060 24548 16112 24600
rect 17716 24548 17768 24600
rect 17992 24591 18044 24600
rect 17992 24557 18001 24591
rect 18001 24557 18035 24591
rect 18035 24557 18044 24591
rect 17992 24548 18044 24557
rect 21212 24591 21264 24600
rect 21212 24557 21221 24591
rect 21221 24557 21255 24591
rect 21255 24557 21264 24591
rect 21212 24548 21264 24557
rect 22960 24591 23012 24600
rect 22960 24557 22969 24591
rect 22969 24557 23003 24591
rect 23003 24557 23012 24591
rect 22960 24548 23012 24557
rect 29216 24548 29268 24600
rect 29768 24591 29820 24600
rect 29768 24557 29777 24591
rect 29777 24557 29811 24591
rect 29811 24557 29820 24591
rect 29768 24548 29820 24557
rect 28388 24523 28440 24532
rect 28388 24489 28397 24523
rect 28397 24489 28431 24523
rect 28431 24489 28440 24523
rect 28388 24480 28440 24489
rect 3088 24412 3140 24464
rect 9528 24455 9580 24464
rect 9528 24421 9537 24455
rect 9537 24421 9571 24455
rect 9571 24421 9580 24455
rect 9528 24412 9580 24421
rect 13944 24412 13996 24464
rect 18452 24455 18504 24464
rect 18452 24421 18461 24455
rect 18461 24421 18495 24455
rect 18495 24421 18504 24455
rect 18452 24412 18504 24421
rect 21580 24412 21632 24464
rect 23420 24412 23472 24464
rect 3510 24310 3562 24362
rect 3574 24310 3626 24362
rect 3638 24310 3690 24362
rect 3702 24310 3754 24362
rect 3766 24310 3818 24362
rect 3916 24208 3968 24260
rect 9068 24208 9120 24260
rect 9528 24251 9580 24260
rect 9528 24217 9537 24251
rect 9537 24217 9571 24251
rect 9571 24217 9580 24251
rect 9528 24208 9580 24217
rect 10448 24251 10500 24260
rect 10448 24217 10457 24251
rect 10457 24217 10491 24251
rect 10491 24217 10500 24251
rect 10448 24208 10500 24217
rect 972 24140 1024 24192
rect 4560 24140 4612 24192
rect 2720 24047 2772 24056
rect 2720 24013 2729 24047
rect 2729 24013 2763 24047
rect 2763 24013 2772 24047
rect 3088 24047 3140 24056
rect 2720 24004 2772 24013
rect 3088 24013 3097 24047
rect 3097 24013 3131 24047
rect 3131 24013 3140 24047
rect 3088 24004 3140 24013
rect 4652 24072 4704 24124
rect 9252 24115 9304 24124
rect 9252 24081 9261 24115
rect 9261 24081 9295 24115
rect 9295 24081 9304 24115
rect 9252 24072 9304 24081
rect 9620 24072 9672 24124
rect 4744 24004 4796 24056
rect 5756 24004 5808 24056
rect 6308 24004 6360 24056
rect 6952 24047 7004 24056
rect 6952 24013 6961 24047
rect 6961 24013 6995 24047
rect 6995 24013 7004 24047
rect 6952 24004 7004 24013
rect 10448 24004 10500 24056
rect 11276 24004 11328 24056
rect 11920 24004 11972 24056
rect 12564 24208 12616 24260
rect 15784 24208 15836 24260
rect 16060 24251 16112 24260
rect 16060 24217 16069 24251
rect 16069 24217 16103 24251
rect 16103 24217 16112 24251
rect 16060 24208 16112 24217
rect 16980 24208 17032 24260
rect 17716 24251 17768 24260
rect 17716 24217 17725 24251
rect 17725 24217 17759 24251
rect 17759 24217 17768 24251
rect 17716 24208 17768 24217
rect 20936 24208 20988 24260
rect 21672 24208 21724 24260
rect 25904 24251 25956 24260
rect 25904 24217 25913 24251
rect 25913 24217 25947 24251
rect 25947 24217 25956 24251
rect 25904 24208 25956 24217
rect 26180 24208 26232 24260
rect 27376 24251 27428 24260
rect 27376 24217 27385 24251
rect 27385 24217 27419 24251
rect 27419 24217 27428 24251
rect 27376 24208 27428 24217
rect 27928 24208 27980 24260
rect 28204 24208 28256 24260
rect 29308 24208 29360 24260
rect 29768 24251 29820 24260
rect 29768 24217 29777 24251
rect 29777 24217 29811 24251
rect 29811 24217 29820 24251
rect 29768 24208 29820 24217
rect 29860 24251 29912 24260
rect 29860 24217 29869 24251
rect 29869 24217 29903 24251
rect 29903 24217 29912 24251
rect 29860 24208 29912 24217
rect 17072 24183 17124 24192
rect 17072 24149 17081 24183
rect 17081 24149 17115 24183
rect 17115 24149 17124 24183
rect 17072 24140 17124 24149
rect 13944 24072 13996 24124
rect 13208 24047 13260 24056
rect 13208 24013 13217 24047
rect 13217 24013 13251 24047
rect 13251 24013 13260 24047
rect 13208 24004 13260 24013
rect 15600 24072 15652 24124
rect 17992 24140 18044 24192
rect 22960 24140 23012 24192
rect 28388 24140 28440 24192
rect 20292 24004 20344 24056
rect 27376 24004 27428 24056
rect 28480 24004 28532 24056
rect 30596 24140 30648 24192
rect 29768 24072 29820 24124
rect 31516 24072 31568 24124
rect 29216 24047 29268 24056
rect 29216 24013 29225 24047
rect 29225 24013 29259 24047
rect 29259 24013 29268 24047
rect 29216 24004 29268 24013
rect 3916 23936 3968 23988
rect 6584 23936 6636 23988
rect 7688 23936 7740 23988
rect 12012 23979 12064 23988
rect 12012 23945 12021 23979
rect 12021 23945 12055 23979
rect 12055 23945 12064 23979
rect 12012 23936 12064 23945
rect 12104 23936 12156 23988
rect 13944 23936 13996 23988
rect 4284 23868 4336 23920
rect 12564 23911 12616 23920
rect 12564 23877 12573 23911
rect 12573 23877 12607 23911
rect 12607 23877 12616 23911
rect 12564 23868 12616 23877
rect 12656 23868 12708 23920
rect 19372 23936 19424 23988
rect 21212 23979 21264 23988
rect 21212 23945 21221 23979
rect 21221 23945 21255 23979
rect 21255 23945 21264 23979
rect 21212 23936 21264 23945
rect 21948 23936 22000 23988
rect 25904 23936 25956 23988
rect 27560 23979 27612 23988
rect 27560 23945 27569 23979
rect 27569 23945 27603 23979
rect 27603 23945 27612 23979
rect 27560 23936 27612 23945
rect 20016 23911 20068 23920
rect 20016 23877 20025 23911
rect 20025 23877 20059 23911
rect 20059 23877 20068 23911
rect 20016 23868 20068 23877
rect 18870 23766 18922 23818
rect 18934 23766 18986 23818
rect 18998 23766 19050 23818
rect 19062 23766 19114 23818
rect 19126 23766 19178 23818
rect 2628 23664 2680 23716
rect 7688 23707 7740 23716
rect 7688 23673 7697 23707
rect 7697 23673 7731 23707
rect 7731 23673 7740 23707
rect 7688 23664 7740 23673
rect 7780 23707 7832 23716
rect 7780 23673 7789 23707
rect 7789 23673 7823 23707
rect 7823 23673 7832 23707
rect 7780 23664 7832 23673
rect 9988 23664 10040 23716
rect 13208 23707 13260 23716
rect 13208 23673 13217 23707
rect 13217 23673 13251 23707
rect 13251 23673 13260 23707
rect 13208 23664 13260 23673
rect 19372 23664 19424 23716
rect 20016 23664 20068 23716
rect 24248 23707 24300 23716
rect 24248 23673 24257 23707
rect 24257 23673 24291 23707
rect 24291 23673 24300 23707
rect 24248 23664 24300 23673
rect 30228 23596 30280 23648
rect 1156 23571 1208 23580
rect 1156 23537 1165 23571
rect 1165 23537 1199 23571
rect 1199 23537 1208 23571
rect 1156 23528 1208 23537
rect 1340 23528 1392 23580
rect 3364 23571 3416 23580
rect 3364 23537 3373 23571
rect 3373 23537 3407 23571
rect 3407 23537 3416 23571
rect 3364 23528 3416 23537
rect 7136 23528 7188 23580
rect 9068 23571 9120 23580
rect 9068 23537 9077 23571
rect 9077 23537 9111 23571
rect 9111 23537 9120 23571
rect 9068 23528 9120 23537
rect 11092 23571 11144 23580
rect 11092 23537 11101 23571
rect 11101 23537 11135 23571
rect 11135 23537 11144 23571
rect 11092 23528 11144 23537
rect 11184 23528 11236 23580
rect 18728 23528 18780 23580
rect 21580 23571 21632 23580
rect 21580 23537 21589 23571
rect 21589 23537 21623 23571
rect 21623 23537 21632 23571
rect 21580 23528 21632 23537
rect 22960 23571 23012 23580
rect 22960 23537 22969 23571
rect 22969 23537 23003 23571
rect 23003 23537 23012 23571
rect 22960 23528 23012 23537
rect 1432 23503 1484 23512
rect 1432 23469 1441 23503
rect 1441 23469 1475 23503
rect 1475 23469 1484 23503
rect 1432 23460 1484 23469
rect 7044 23503 7096 23512
rect 7044 23469 7053 23503
rect 7053 23469 7087 23503
rect 7087 23469 7096 23503
rect 7044 23460 7096 23469
rect 9528 23460 9580 23512
rect 10908 23503 10960 23512
rect 10908 23469 10917 23503
rect 10917 23469 10951 23503
rect 10951 23469 10960 23503
rect 10908 23460 10960 23469
rect 11460 23503 11512 23512
rect 11460 23469 11469 23503
rect 11469 23469 11503 23503
rect 11503 23469 11512 23503
rect 11460 23460 11512 23469
rect 18268 23460 18320 23512
rect 22868 23460 22920 23512
rect 26916 23528 26968 23580
rect 27284 23528 27336 23580
rect 27560 23571 27612 23580
rect 27560 23537 27569 23571
rect 27569 23537 27603 23571
rect 27603 23537 27612 23571
rect 27560 23528 27612 23537
rect 28480 23571 28532 23580
rect 27468 23460 27520 23512
rect 28480 23537 28489 23571
rect 28489 23537 28523 23571
rect 28523 23537 28532 23571
rect 28480 23528 28532 23537
rect 30044 23528 30096 23580
rect 30412 23460 30464 23512
rect 12104 23392 12156 23444
rect 12840 23392 12892 23444
rect 27008 23392 27060 23444
rect 27192 23435 27244 23444
rect 27192 23401 27201 23435
rect 27201 23401 27235 23435
rect 27235 23401 27244 23435
rect 27192 23392 27244 23401
rect 1984 23324 2036 23376
rect 3088 23324 3140 23376
rect 4008 23324 4060 23376
rect 7320 23324 7372 23376
rect 12380 23367 12432 23376
rect 12380 23333 12389 23367
rect 12389 23333 12423 23367
rect 12423 23333 12432 23367
rect 12380 23324 12432 23333
rect 17992 23324 18044 23376
rect 21488 23324 21540 23376
rect 21672 23367 21724 23376
rect 21672 23333 21681 23367
rect 21681 23333 21715 23367
rect 21715 23333 21724 23367
rect 21672 23324 21724 23333
rect 23144 23324 23196 23376
rect 24800 23324 24852 23376
rect 3510 23222 3562 23274
rect 3574 23222 3626 23274
rect 3638 23222 3690 23274
rect 3702 23222 3754 23274
rect 3766 23222 3818 23274
rect 4560 23120 4612 23172
rect 5756 23163 5808 23172
rect 5756 23129 5765 23163
rect 5765 23129 5799 23163
rect 5799 23129 5808 23163
rect 5756 23120 5808 23129
rect 6584 23052 6636 23104
rect 7136 23120 7188 23172
rect 7872 23120 7924 23172
rect 10264 23120 10316 23172
rect 12104 23120 12156 23172
rect 12380 23120 12432 23172
rect 13208 23120 13260 23172
rect 14956 23163 15008 23172
rect 972 23027 1024 23036
rect 972 22993 981 23027
rect 981 22993 1015 23027
rect 1015 22993 1024 23027
rect 972 22984 1024 22993
rect 1984 22984 2036 23036
rect 3364 23027 3416 23036
rect 3364 22993 3373 23027
rect 3373 22993 3407 23027
rect 3407 22993 3416 23027
rect 3364 22984 3416 22993
rect 696 22959 748 22968
rect 696 22925 705 22959
rect 705 22925 739 22959
rect 739 22925 748 22959
rect 696 22916 748 22925
rect 6308 23027 6360 23036
rect 6308 22993 6317 23027
rect 6317 22993 6351 23027
rect 6351 22993 6360 23027
rect 6308 22984 6360 22993
rect 11460 23052 11512 23104
rect 11092 23027 11144 23036
rect 11092 22993 11101 23027
rect 11101 22993 11135 23027
rect 11135 22993 11144 23027
rect 11092 22984 11144 22993
rect 11920 23027 11972 23036
rect 11920 22993 11929 23027
rect 11929 22993 11963 23027
rect 11963 22993 11972 23027
rect 11920 22984 11972 22993
rect 6492 22959 6544 22968
rect 6492 22925 6501 22959
rect 6501 22925 6535 22959
rect 6535 22925 6544 22959
rect 6492 22916 6544 22925
rect 7320 22959 7372 22968
rect 7320 22925 7329 22959
rect 7329 22925 7363 22959
rect 7363 22925 7372 22959
rect 7320 22916 7372 22925
rect 1432 22848 1484 22900
rect 2904 22848 2956 22900
rect 4376 22891 4428 22900
rect 4376 22857 4385 22891
rect 4385 22857 4419 22891
rect 4419 22857 4428 22891
rect 4376 22848 4428 22857
rect 4008 22780 4060 22832
rect 8148 22916 8200 22968
rect 12656 22959 12708 22968
rect 12656 22925 12665 22959
rect 12665 22925 12699 22959
rect 12699 22925 12708 22959
rect 12656 22916 12708 22925
rect 12840 22959 12892 22968
rect 12840 22925 12849 22959
rect 12849 22925 12883 22959
rect 12883 22925 12892 22959
rect 12840 22916 12892 22925
rect 13208 22959 13260 22968
rect 13208 22925 13217 22959
rect 13217 22925 13251 22959
rect 13251 22925 13260 22959
rect 13208 22916 13260 22925
rect 14956 23129 14965 23163
rect 14965 23129 14999 23163
rect 14999 23129 15008 23163
rect 14956 23120 15008 23129
rect 17992 23163 18044 23172
rect 17992 23129 18001 23163
rect 18001 23129 18035 23163
rect 18035 23129 18044 23163
rect 17992 23120 18044 23129
rect 18728 23120 18780 23172
rect 21672 23120 21724 23172
rect 24248 23163 24300 23172
rect 24248 23129 24257 23163
rect 24257 23129 24291 23163
rect 24291 23129 24300 23163
rect 24248 23120 24300 23129
rect 24524 23120 24576 23172
rect 26916 23163 26968 23172
rect 24156 23052 24208 23104
rect 18636 23027 18688 23036
rect 18636 22993 18645 23027
rect 18645 22993 18679 23027
rect 18679 22993 18688 23027
rect 18636 22984 18688 22993
rect 22960 22984 23012 23036
rect 24432 23027 24484 23036
rect 21580 22959 21632 22968
rect 21580 22925 21589 22959
rect 21589 22925 21623 22959
rect 21623 22925 21632 22959
rect 21580 22916 21632 22925
rect 22684 22916 22736 22968
rect 23144 22916 23196 22968
rect 24432 22993 24441 23027
rect 24441 22993 24475 23027
rect 24475 22993 24484 23027
rect 24432 22984 24484 22993
rect 26916 23129 26925 23163
rect 26925 23129 26959 23163
rect 26959 23129 26968 23163
rect 26916 23120 26968 23129
rect 27192 23120 27244 23172
rect 30412 23163 30464 23172
rect 30412 23129 30421 23163
rect 30421 23129 30455 23163
rect 30455 23129 30464 23163
rect 30412 23120 30464 23129
rect 27468 23095 27520 23104
rect 27468 23061 27477 23095
rect 27477 23061 27511 23095
rect 27511 23061 27520 23095
rect 27468 23052 27520 23061
rect 24616 22959 24668 22968
rect 24616 22925 24625 22959
rect 24625 22925 24659 22959
rect 24659 22925 24668 22959
rect 24616 22916 24668 22925
rect 24800 22916 24852 22968
rect 25996 22959 26048 22968
rect 25996 22925 26005 22959
rect 26005 22925 26039 22959
rect 26039 22925 26048 22959
rect 25996 22916 26048 22925
rect 27560 22984 27612 23036
rect 9068 22848 9120 22900
rect 14956 22848 15008 22900
rect 18084 22848 18136 22900
rect 19372 22848 19424 22900
rect 20660 22891 20712 22900
rect 20660 22857 20669 22891
rect 20669 22857 20703 22891
rect 20703 22857 20712 22891
rect 20660 22848 20712 22857
rect 23972 22848 24024 22900
rect 27192 22916 27244 22968
rect 27284 22916 27336 22968
rect 28480 23052 28532 23104
rect 30044 23052 30096 23104
rect 30136 23095 30188 23104
rect 30136 23061 30145 23095
rect 30145 23061 30179 23095
rect 30179 23061 30188 23095
rect 30136 23052 30188 23061
rect 27928 22848 27980 22900
rect 9528 22780 9580 22832
rect 10908 22780 10960 22832
rect 11184 22780 11236 22832
rect 11920 22780 11972 22832
rect 13024 22780 13076 22832
rect 18268 22823 18320 22832
rect 18268 22789 18277 22823
rect 18277 22789 18311 22823
rect 18311 22789 18320 22823
rect 18268 22780 18320 22789
rect 22868 22780 22920 22832
rect 27008 22780 27060 22832
rect 30228 22823 30280 22832
rect 30228 22789 30237 22823
rect 30237 22789 30271 22823
rect 30271 22789 30280 22823
rect 30228 22780 30280 22789
rect 18870 22678 18922 22730
rect 18934 22678 18986 22730
rect 18998 22678 19050 22730
rect 19062 22678 19114 22730
rect 19126 22678 19178 22730
rect 972 22576 1024 22628
rect 1432 22576 1484 22628
rect 2628 22576 2680 22628
rect 6308 22576 6360 22628
rect 6492 22619 6544 22628
rect 6492 22585 6501 22619
rect 6501 22585 6535 22619
rect 6535 22585 6544 22619
rect 6492 22576 6544 22585
rect 13208 22576 13260 22628
rect 15692 22576 15744 22628
rect 18636 22576 18688 22628
rect 19372 22576 19424 22628
rect 6952 22508 7004 22560
rect 10724 22508 10776 22560
rect 21856 22508 21908 22560
rect 23972 22576 24024 22628
rect 24432 22576 24484 22628
rect 3272 22440 3324 22492
rect 4100 22483 4152 22492
rect 4100 22449 4109 22483
rect 4109 22449 4143 22483
rect 4143 22449 4152 22483
rect 4100 22440 4152 22449
rect 4560 22483 4612 22492
rect 4560 22449 4569 22483
rect 4569 22449 4603 22483
rect 4603 22449 4612 22483
rect 4560 22440 4612 22449
rect 4928 22440 4980 22492
rect 6124 22440 6176 22492
rect 8148 22440 8200 22492
rect 9988 22483 10040 22492
rect 9988 22449 9997 22483
rect 9997 22449 10031 22483
rect 10031 22449 10040 22483
rect 9988 22440 10040 22449
rect 13024 22483 13076 22492
rect 13024 22449 13033 22483
rect 13033 22449 13067 22483
rect 13067 22449 13076 22483
rect 13024 22440 13076 22449
rect 15140 22440 15192 22492
rect 15968 22440 16020 22492
rect 16336 22483 16388 22492
rect 16336 22449 16345 22483
rect 16345 22449 16379 22483
rect 16379 22449 16388 22483
rect 16336 22440 16388 22449
rect 21764 22440 21816 22492
rect 22684 22483 22736 22492
rect 22684 22449 22693 22483
rect 22693 22449 22727 22483
rect 22727 22449 22736 22483
rect 22684 22440 22736 22449
rect 22960 22483 23012 22492
rect 22960 22449 22969 22483
rect 22969 22449 23003 22483
rect 23003 22449 23012 22483
rect 22960 22440 23012 22449
rect 23236 22508 23288 22560
rect 27100 22508 27152 22560
rect 26180 22440 26232 22492
rect 5940 22372 5992 22424
rect 7596 22415 7648 22424
rect 7596 22381 7605 22415
rect 7605 22381 7639 22415
rect 7639 22381 7648 22415
rect 7596 22372 7648 22381
rect 10724 22372 10776 22424
rect 10908 22372 10960 22424
rect 11552 22372 11604 22424
rect 14772 22372 14824 22424
rect 23236 22372 23288 22424
rect 25996 22372 26048 22424
rect 26916 22440 26968 22492
rect 28572 22483 28624 22492
rect 3180 22304 3232 22356
rect 3916 22304 3968 22356
rect 4192 22304 4244 22356
rect 5572 22304 5624 22356
rect 7044 22304 7096 22356
rect 15692 22304 15744 22356
rect 25812 22347 25864 22356
rect 25812 22313 25821 22347
rect 25821 22313 25855 22347
rect 25855 22313 25864 22347
rect 25812 22304 25864 22313
rect 25904 22347 25956 22356
rect 25904 22313 25913 22347
rect 25913 22313 25947 22347
rect 25947 22313 25956 22347
rect 25904 22304 25956 22313
rect 696 22236 748 22288
rect 1340 22279 1392 22288
rect 1340 22245 1349 22279
rect 1349 22245 1383 22279
rect 1383 22245 1392 22279
rect 1340 22236 1392 22245
rect 6308 22279 6360 22288
rect 6308 22245 6317 22279
rect 6317 22245 6351 22279
rect 6351 22245 6360 22279
rect 6308 22236 6360 22245
rect 12656 22236 12708 22288
rect 16520 22236 16572 22288
rect 16612 22279 16664 22288
rect 16612 22245 16621 22279
rect 16621 22245 16655 22279
rect 16655 22245 16664 22279
rect 16612 22236 16664 22245
rect 17624 22236 17676 22288
rect 20660 22236 20712 22288
rect 25536 22236 25588 22288
rect 26272 22236 26324 22288
rect 28572 22449 28581 22483
rect 28581 22449 28615 22483
rect 28615 22449 28624 22483
rect 28572 22440 28624 22449
rect 28756 22440 28808 22492
rect 28848 22279 28900 22288
rect 28848 22245 28857 22279
rect 28857 22245 28891 22279
rect 28891 22245 28900 22279
rect 28848 22236 28900 22245
rect 3510 22134 3562 22186
rect 3574 22134 3626 22186
rect 3638 22134 3690 22186
rect 3702 22134 3754 22186
rect 3766 22134 3818 22186
rect 2904 22075 2956 22084
rect 2904 22041 2913 22075
rect 2913 22041 2947 22075
rect 2947 22041 2956 22075
rect 2904 22032 2956 22041
rect 3272 22075 3324 22084
rect 3272 22041 3281 22075
rect 3281 22041 3315 22075
rect 3315 22041 3324 22075
rect 3272 22032 3324 22041
rect 4100 22032 4152 22084
rect 4192 22032 4244 22084
rect 5940 22075 5992 22084
rect 5940 22041 5949 22075
rect 5949 22041 5983 22075
rect 5983 22041 5992 22075
rect 8148 22075 8200 22084
rect 5940 22032 5992 22041
rect 4744 21964 4796 22016
rect 4928 22007 4980 22016
rect 4928 21973 4937 22007
rect 4937 21973 4971 22007
rect 4971 21973 4980 22007
rect 4928 21964 4980 21973
rect 6492 22007 6544 22016
rect 6492 21973 6501 22007
rect 6501 21973 6535 22007
rect 6535 21973 6544 22007
rect 6492 21964 6544 21973
rect 4284 21939 4336 21948
rect 4284 21905 4293 21939
rect 4293 21905 4327 21939
rect 4327 21905 4336 21939
rect 4284 21896 4336 21905
rect 8148 22041 8157 22075
rect 8157 22041 8191 22075
rect 8191 22041 8200 22075
rect 8148 22032 8200 22041
rect 10816 22032 10868 22084
rect 16520 22032 16572 22084
rect 21764 22075 21816 22084
rect 10908 21964 10960 22016
rect 11460 21964 11512 22016
rect 16612 22007 16664 22016
rect 4008 21871 4060 21880
rect 2720 21692 2772 21744
rect 3180 21692 3232 21744
rect 4008 21837 4017 21871
rect 4017 21837 4051 21871
rect 4051 21837 4060 21871
rect 4008 21828 4060 21837
rect 4100 21828 4152 21880
rect 4744 21828 4796 21880
rect 6124 21871 6176 21880
rect 6124 21837 6133 21871
rect 6133 21837 6167 21871
rect 6167 21837 6176 21871
rect 6124 21828 6176 21837
rect 6400 21828 6452 21880
rect 11000 21896 11052 21948
rect 13300 21896 13352 21948
rect 16612 21973 16621 22007
rect 16621 21973 16655 22007
rect 16655 21973 16664 22007
rect 16612 21964 16664 21973
rect 21764 22041 21773 22075
rect 21773 22041 21807 22075
rect 21807 22041 21816 22075
rect 21764 22032 21816 22041
rect 21856 22032 21908 22084
rect 25904 22032 25956 22084
rect 28572 22075 28624 22084
rect 28572 22041 28581 22075
rect 28581 22041 28615 22075
rect 28615 22041 28624 22075
rect 28572 22032 28624 22041
rect 28756 22075 28808 22084
rect 28756 22041 28765 22075
rect 28765 22041 28799 22075
rect 28799 22041 28808 22075
rect 28756 22032 28808 22041
rect 28848 22032 28900 22084
rect 22684 21964 22736 22016
rect 25536 22007 25588 22016
rect 25536 21973 25545 22007
rect 25545 21973 25579 22007
rect 25579 21973 25588 22007
rect 25536 21964 25588 21973
rect 26180 21964 26232 22016
rect 26364 21964 26416 22016
rect 28664 21964 28716 22016
rect 30228 21964 30280 22016
rect 18084 21939 18136 21948
rect 7780 21871 7832 21880
rect 4836 21692 4888 21744
rect 7780 21837 7789 21871
rect 7789 21837 7823 21871
rect 7823 21837 7832 21871
rect 7780 21828 7832 21837
rect 9988 21828 10040 21880
rect 12196 21828 12248 21880
rect 14772 21828 14824 21880
rect 18084 21905 18093 21939
rect 18093 21905 18127 21939
rect 18127 21905 18136 21939
rect 18084 21896 18136 21905
rect 22776 21896 22828 21948
rect 23144 21896 23196 21948
rect 26916 21939 26968 21948
rect 26916 21905 26925 21939
rect 26925 21905 26959 21939
rect 26959 21905 26968 21939
rect 26916 21896 26968 21905
rect 10724 21760 10776 21812
rect 12012 21760 12064 21812
rect 17624 21871 17676 21880
rect 17624 21837 17633 21871
rect 17633 21837 17667 21871
rect 17667 21837 17676 21871
rect 17624 21828 17676 21837
rect 18360 21828 18412 21880
rect 21488 21828 21540 21880
rect 22960 21828 23012 21880
rect 26364 21871 26416 21880
rect 26364 21837 26373 21871
rect 26373 21837 26407 21871
rect 26407 21837 26416 21871
rect 26364 21828 26416 21837
rect 26456 21828 26508 21880
rect 18268 21760 18320 21812
rect 24524 21760 24576 21812
rect 8700 21692 8752 21744
rect 12656 21735 12708 21744
rect 12656 21701 12665 21735
rect 12665 21701 12699 21735
rect 12699 21701 12708 21735
rect 12656 21692 12708 21701
rect 13024 21692 13076 21744
rect 15140 21692 15192 21744
rect 16336 21735 16388 21744
rect 16336 21701 16345 21735
rect 16345 21701 16379 21735
rect 16379 21701 16388 21735
rect 16336 21692 16388 21701
rect 18728 21735 18780 21744
rect 18728 21701 18737 21735
rect 18737 21701 18771 21735
rect 18771 21701 18780 21735
rect 18728 21692 18780 21701
rect 23236 21692 23288 21744
rect 25996 21735 26048 21744
rect 25996 21701 26005 21735
rect 26005 21701 26039 21735
rect 26039 21701 26048 21735
rect 25996 21692 26048 21701
rect 27100 21735 27152 21744
rect 27100 21701 27109 21735
rect 27109 21701 27143 21735
rect 27143 21701 27152 21735
rect 27100 21692 27152 21701
rect 18870 21590 18922 21642
rect 18934 21590 18986 21642
rect 18998 21590 19050 21642
rect 19062 21590 19114 21642
rect 19126 21590 19178 21642
rect 4560 21488 4612 21540
rect 7228 21488 7280 21540
rect 7596 21488 7648 21540
rect 13300 21488 13352 21540
rect 14772 21531 14824 21540
rect 14772 21497 14781 21531
rect 14781 21497 14815 21531
rect 14815 21497 14824 21531
rect 14772 21488 14824 21497
rect 17348 21488 17400 21540
rect 23420 21531 23472 21540
rect 23420 21497 23429 21531
rect 23429 21497 23463 21531
rect 23463 21497 23472 21531
rect 23420 21488 23472 21497
rect 27560 21488 27612 21540
rect 4284 21420 4336 21472
rect 7044 21420 7096 21472
rect 16428 21420 16480 21472
rect 1340 21352 1392 21404
rect 3916 21352 3968 21404
rect 4376 21395 4428 21404
rect 4376 21361 4385 21395
rect 4385 21361 4419 21395
rect 4419 21361 4428 21395
rect 4376 21352 4428 21361
rect 4744 21395 4796 21404
rect 4744 21361 4753 21395
rect 4753 21361 4787 21395
rect 4787 21361 4796 21395
rect 4744 21352 4796 21361
rect 5848 21352 5900 21404
rect 7596 21352 7648 21404
rect 10908 21352 10960 21404
rect 11092 21352 11144 21404
rect 11460 21395 11512 21404
rect 11460 21361 11469 21395
rect 11469 21361 11503 21395
rect 11503 21361 11512 21395
rect 11460 21352 11512 21361
rect 12840 21395 12892 21404
rect 12840 21361 12849 21395
rect 12849 21361 12883 21395
rect 12883 21361 12892 21395
rect 12840 21352 12892 21361
rect 15324 21352 15376 21404
rect 16520 21352 16572 21404
rect 18360 21395 18412 21404
rect 1432 21327 1484 21336
rect 1432 21293 1441 21327
rect 1441 21293 1475 21327
rect 1475 21293 1484 21327
rect 1432 21284 1484 21293
rect 3364 21284 3416 21336
rect 4192 21216 4244 21268
rect 4560 21284 4612 21336
rect 5572 21284 5624 21336
rect 5756 21327 5808 21336
rect 5756 21293 5765 21327
rect 5765 21293 5799 21327
rect 5799 21293 5808 21327
rect 5756 21284 5808 21293
rect 6308 21327 6360 21336
rect 6308 21293 6317 21327
rect 6317 21293 6351 21327
rect 6351 21293 6360 21327
rect 6308 21284 6360 21293
rect 6400 21284 6452 21336
rect 10724 21284 10776 21336
rect 10816 21284 10868 21336
rect 11828 21284 11880 21336
rect 13024 21327 13076 21336
rect 7780 21216 7832 21268
rect 11184 21216 11236 21268
rect 13024 21293 13033 21327
rect 13033 21293 13067 21327
rect 13067 21293 13076 21327
rect 13024 21284 13076 21293
rect 17072 21327 17124 21336
rect 17072 21293 17081 21327
rect 17081 21293 17115 21327
rect 17115 21293 17124 21327
rect 17072 21284 17124 21293
rect 17440 21284 17492 21336
rect 18360 21361 18369 21395
rect 18369 21361 18403 21395
rect 18403 21361 18412 21395
rect 18360 21352 18412 21361
rect 19372 21352 19424 21404
rect 21948 21420 22000 21472
rect 22132 21352 22184 21404
rect 22316 21395 22368 21404
rect 22316 21361 22325 21395
rect 22325 21361 22359 21395
rect 22359 21361 22368 21395
rect 22316 21352 22368 21361
rect 22592 21395 22644 21404
rect 22592 21361 22601 21395
rect 22601 21361 22635 21395
rect 22635 21361 22644 21395
rect 22592 21352 22644 21361
rect 23236 21395 23288 21404
rect 23236 21361 23245 21395
rect 23245 21361 23279 21395
rect 23279 21361 23288 21395
rect 23236 21352 23288 21361
rect 24156 21352 24208 21404
rect 27008 21395 27060 21404
rect 27008 21361 27017 21395
rect 27017 21361 27051 21395
rect 27051 21361 27060 21395
rect 27008 21352 27060 21361
rect 27468 21352 27520 21404
rect 27744 21395 27796 21404
rect 27744 21361 27753 21395
rect 27753 21361 27787 21395
rect 27787 21361 27796 21395
rect 27744 21352 27796 21361
rect 16244 21216 16296 21268
rect 18728 21284 18780 21336
rect 22868 21327 22920 21336
rect 22868 21293 22877 21327
rect 22877 21293 22911 21327
rect 22911 21293 22920 21327
rect 22868 21284 22920 21293
rect 24524 21327 24576 21336
rect 24524 21293 24533 21327
rect 24533 21293 24567 21327
rect 24567 21293 24576 21327
rect 25812 21327 25864 21336
rect 24524 21284 24576 21293
rect 25812 21293 25821 21327
rect 25821 21293 25855 21327
rect 25855 21293 25864 21327
rect 25812 21284 25864 21293
rect 26732 21284 26784 21336
rect 27652 21284 27704 21336
rect 28572 21352 28624 21404
rect 29584 21284 29636 21336
rect 2720 21148 2772 21200
rect 4008 21148 4060 21200
rect 4560 21148 4612 21200
rect 6952 21191 7004 21200
rect 6952 21157 6961 21191
rect 6961 21157 6995 21191
rect 6995 21157 7004 21191
rect 6952 21148 7004 21157
rect 9068 21148 9120 21200
rect 22776 21148 22828 21200
rect 23788 21148 23840 21200
rect 25168 21148 25220 21200
rect 28296 21148 28348 21200
rect 28572 21148 28624 21200
rect 3510 21046 3562 21098
rect 3574 21046 3626 21098
rect 3638 21046 3690 21098
rect 3702 21046 3754 21098
rect 3766 21046 3818 21098
rect 3364 20987 3416 20996
rect 3364 20953 3373 20987
rect 3373 20953 3407 20987
rect 3407 20953 3416 20987
rect 3364 20944 3416 20953
rect 3916 20944 3968 20996
rect 4376 20944 4428 20996
rect 4928 20944 4980 20996
rect 5848 20987 5900 20996
rect 5848 20953 5857 20987
rect 5857 20953 5891 20987
rect 5891 20953 5900 20987
rect 5848 20944 5900 20953
rect 7872 20944 7924 20996
rect 10724 20987 10776 20996
rect 10724 20953 10733 20987
rect 10733 20953 10767 20987
rect 10767 20953 10776 20987
rect 10724 20944 10776 20953
rect 11092 20987 11144 20996
rect 11092 20953 11101 20987
rect 11101 20953 11135 20987
rect 11135 20953 11144 20987
rect 11092 20944 11144 20953
rect 11368 20944 11420 20996
rect 12840 20987 12892 20996
rect 12840 20953 12849 20987
rect 12849 20953 12883 20987
rect 12883 20953 12892 20987
rect 12840 20944 12892 20953
rect 13024 20987 13076 20996
rect 13024 20953 13033 20987
rect 13033 20953 13067 20987
rect 13067 20953 13076 20987
rect 13024 20944 13076 20953
rect 16244 20987 16296 20996
rect 16244 20953 16253 20987
rect 16253 20953 16287 20987
rect 16287 20953 16296 20987
rect 16244 20944 16296 20953
rect 16428 20987 16480 20996
rect 16428 20953 16437 20987
rect 16437 20953 16471 20987
rect 16471 20953 16480 20987
rect 16428 20944 16480 20953
rect 17072 20944 17124 20996
rect 17164 20987 17216 20996
rect 17164 20953 17173 20987
rect 17173 20953 17207 20987
rect 17207 20953 17216 20987
rect 17164 20944 17216 20953
rect 18360 20944 18412 20996
rect 21948 20987 22000 20996
rect 21948 20953 21957 20987
rect 21957 20953 21991 20987
rect 21991 20953 22000 20987
rect 21948 20944 22000 20953
rect 22132 20987 22184 20996
rect 22132 20953 22141 20987
rect 22141 20953 22175 20987
rect 22175 20953 22184 20987
rect 22132 20944 22184 20953
rect 2720 20851 2772 20860
rect 2720 20817 2729 20851
rect 2729 20817 2763 20851
rect 2763 20817 2772 20851
rect 2720 20808 2772 20817
rect 4008 20808 4060 20860
rect 4192 20851 4244 20860
rect 4192 20817 4201 20851
rect 4201 20817 4235 20851
rect 4235 20817 4244 20851
rect 4192 20808 4244 20817
rect 696 20783 748 20792
rect 696 20749 705 20783
rect 705 20749 739 20783
rect 739 20749 748 20783
rect 696 20740 748 20749
rect 4100 20740 4152 20792
rect 4468 20808 4520 20860
rect 4744 20808 4796 20860
rect 4928 20740 4980 20792
rect 788 20604 840 20656
rect 1432 20672 1484 20724
rect 6308 20876 6360 20928
rect 8700 20876 8752 20928
rect 7228 20851 7280 20860
rect 7228 20817 7237 20851
rect 7237 20817 7271 20851
rect 7271 20817 7280 20851
rect 7228 20808 7280 20817
rect 6216 20783 6268 20792
rect 6216 20749 6225 20783
rect 6225 20749 6259 20783
rect 6259 20749 6268 20783
rect 6216 20740 6268 20749
rect 7688 20783 7740 20792
rect 7688 20749 7697 20783
rect 7697 20749 7731 20783
rect 7731 20749 7740 20783
rect 7688 20740 7740 20749
rect 7872 20783 7924 20792
rect 7872 20749 7881 20783
rect 7881 20749 7915 20783
rect 7915 20749 7924 20783
rect 7872 20740 7924 20749
rect 7044 20672 7096 20724
rect 12656 20808 12708 20860
rect 22592 20876 22644 20928
rect 22776 20919 22828 20928
rect 22776 20885 22785 20919
rect 22785 20885 22819 20919
rect 22819 20885 22828 20919
rect 22776 20876 22828 20885
rect 23420 20944 23472 20996
rect 24156 20944 24208 20996
rect 24524 20987 24576 20996
rect 24524 20953 24533 20987
rect 24533 20953 24567 20987
rect 24567 20953 24576 20987
rect 24524 20944 24576 20953
rect 26732 20944 26784 20996
rect 27468 20944 27520 20996
rect 27652 20987 27704 20996
rect 27652 20953 27661 20987
rect 27661 20953 27695 20987
rect 27695 20953 27704 20987
rect 27652 20944 27704 20953
rect 29308 20944 29360 20996
rect 17716 20808 17768 20860
rect 23236 20808 23288 20860
rect 9068 20783 9120 20792
rect 9068 20749 9077 20783
rect 9077 20749 9111 20783
rect 9111 20749 9120 20783
rect 9068 20740 9120 20749
rect 9528 20783 9580 20792
rect 9528 20749 9537 20783
rect 9537 20749 9571 20783
rect 9571 20749 9580 20783
rect 9528 20740 9580 20749
rect 10540 20740 10592 20792
rect 11460 20740 11512 20792
rect 6952 20647 7004 20656
rect 6952 20613 6961 20647
rect 6961 20613 6995 20647
rect 6995 20613 7004 20647
rect 6952 20604 7004 20613
rect 7136 20604 7188 20656
rect 10908 20672 10960 20724
rect 17164 20740 17216 20792
rect 17348 20783 17400 20792
rect 17348 20749 17357 20783
rect 17357 20749 17391 20783
rect 17391 20749 17400 20783
rect 17348 20740 17400 20749
rect 18084 20672 18136 20724
rect 19372 20715 19424 20724
rect 19372 20681 19381 20715
rect 19381 20681 19415 20715
rect 19415 20681 19424 20715
rect 19372 20672 19424 20681
rect 9804 20604 9856 20656
rect 10264 20604 10316 20656
rect 10816 20604 10868 20656
rect 11184 20604 11236 20656
rect 11644 20604 11696 20656
rect 16520 20647 16572 20656
rect 16520 20613 16529 20647
rect 16529 20613 16563 20647
rect 16563 20613 16572 20647
rect 16520 20604 16572 20613
rect 22868 20740 22920 20792
rect 23420 20783 23472 20792
rect 23420 20749 23429 20783
rect 23429 20749 23463 20783
rect 23463 20749 23472 20783
rect 23420 20740 23472 20749
rect 23604 20783 23656 20792
rect 23604 20749 23613 20783
rect 23613 20749 23647 20783
rect 23647 20749 23656 20783
rect 23604 20740 23656 20749
rect 22316 20715 22368 20724
rect 22316 20681 22325 20715
rect 22325 20681 22359 20715
rect 22359 20681 22368 20715
rect 22316 20672 22368 20681
rect 22132 20604 22184 20656
rect 27560 20876 27612 20928
rect 28480 20876 28532 20928
rect 23788 20808 23840 20860
rect 27008 20808 27060 20860
rect 28572 20851 28624 20860
rect 28572 20817 28581 20851
rect 28581 20817 28615 20851
rect 28615 20817 28624 20851
rect 28572 20808 28624 20817
rect 24616 20740 24668 20792
rect 27744 20740 27796 20792
rect 25996 20672 26048 20724
rect 27652 20672 27704 20724
rect 29308 20672 29360 20724
rect 28112 20647 28164 20656
rect 28112 20613 28121 20647
rect 28121 20613 28155 20647
rect 28155 20613 28164 20647
rect 28112 20604 28164 20613
rect 28296 20647 28348 20656
rect 28296 20613 28305 20647
rect 28305 20613 28339 20647
rect 28339 20613 28348 20647
rect 28296 20604 28348 20613
rect 18870 20502 18922 20554
rect 18934 20502 18986 20554
rect 18998 20502 19050 20554
rect 19062 20502 19114 20554
rect 19126 20502 19178 20554
rect 1432 20400 1484 20452
rect 2628 20400 2680 20452
rect 5756 20400 5808 20452
rect 8700 20443 8752 20452
rect 8700 20409 8709 20443
rect 8709 20409 8743 20443
rect 8743 20409 8752 20443
rect 8700 20400 8752 20409
rect 9068 20400 9120 20452
rect 16520 20400 16572 20452
rect 1340 20375 1392 20384
rect 1340 20341 1349 20375
rect 1349 20341 1383 20375
rect 1383 20341 1392 20375
rect 1340 20332 1392 20341
rect 7780 20375 7832 20384
rect 7780 20341 7789 20375
rect 7789 20341 7823 20375
rect 7823 20341 7832 20375
rect 7780 20332 7832 20341
rect 2720 20264 2772 20316
rect 3180 20264 3232 20316
rect 6400 20264 6452 20316
rect 7044 20307 7096 20316
rect 7044 20273 7053 20307
rect 7053 20273 7087 20307
rect 7087 20273 7096 20307
rect 7044 20264 7096 20273
rect 7320 20264 7372 20316
rect 9252 20307 9304 20316
rect 9252 20273 9261 20307
rect 9261 20273 9295 20307
rect 9295 20273 9304 20307
rect 9252 20264 9304 20273
rect 14956 20332 15008 20384
rect 17072 20400 17124 20452
rect 23420 20400 23472 20452
rect 27192 20400 27244 20452
rect 28388 20400 28440 20452
rect 18084 20375 18136 20384
rect 18084 20341 18093 20375
rect 18093 20341 18127 20375
rect 18127 20341 18136 20375
rect 18084 20332 18136 20341
rect 21396 20332 21448 20384
rect 21764 20332 21816 20384
rect 21856 20332 21908 20384
rect 23604 20332 23656 20384
rect 6676 20196 6728 20248
rect 8976 20196 9028 20248
rect 11184 20264 11236 20316
rect 11644 20307 11696 20316
rect 11644 20273 11653 20307
rect 11653 20273 11687 20307
rect 11687 20273 11696 20307
rect 11644 20264 11696 20273
rect 16428 20264 16480 20316
rect 11092 20239 11144 20248
rect 11092 20205 11101 20239
rect 11101 20205 11135 20239
rect 11135 20205 11144 20239
rect 11092 20196 11144 20205
rect 11736 20239 11788 20248
rect 11736 20205 11745 20239
rect 11745 20205 11779 20239
rect 11779 20205 11788 20239
rect 11736 20196 11788 20205
rect 11828 20196 11880 20248
rect 17440 20264 17492 20316
rect 17808 20307 17860 20316
rect 17808 20273 17817 20307
rect 17817 20273 17851 20307
rect 17851 20273 17860 20307
rect 17808 20264 17860 20273
rect 21028 20264 21080 20316
rect 21672 20264 21724 20316
rect 23236 20264 23288 20316
rect 26548 20264 26600 20316
rect 27376 20307 27428 20316
rect 27376 20273 27385 20307
rect 27385 20273 27419 20307
rect 27419 20273 27428 20307
rect 27376 20264 27428 20273
rect 28020 20332 28072 20384
rect 28848 20332 28900 20384
rect 27836 20307 27888 20316
rect 27836 20273 27845 20307
rect 27845 20273 27879 20307
rect 27879 20273 27888 20307
rect 27836 20264 27888 20273
rect 28388 20307 28440 20316
rect 28388 20273 28408 20307
rect 28408 20273 28440 20307
rect 696 20128 748 20180
rect 6860 20128 6912 20180
rect 7320 20171 7372 20180
rect 7320 20137 7329 20171
rect 7329 20137 7363 20171
rect 7363 20137 7372 20171
rect 7320 20128 7372 20137
rect 11368 20128 11420 20180
rect 12012 20171 12064 20180
rect 12012 20137 12021 20171
rect 12021 20137 12055 20171
rect 12055 20137 12064 20171
rect 12012 20128 12064 20137
rect 12196 20128 12248 20180
rect 14680 20128 14732 20180
rect 17348 20128 17400 20180
rect 22040 20239 22092 20248
rect 22040 20205 22049 20239
rect 22049 20205 22083 20239
rect 22083 20205 22092 20239
rect 22040 20196 22092 20205
rect 27468 20196 27520 20248
rect 28388 20264 28440 20273
rect 28204 20196 28256 20248
rect 29492 20196 29544 20248
rect 30136 20196 30188 20248
rect 28296 20128 28348 20180
rect 788 20103 840 20112
rect 788 20069 797 20103
rect 797 20069 831 20103
rect 831 20069 840 20103
rect 788 20060 840 20069
rect 3272 20060 3324 20112
rect 4836 20060 4888 20112
rect 7688 20060 7740 20112
rect 8148 20060 8200 20112
rect 9804 20060 9856 20112
rect 12104 20103 12156 20112
rect 12104 20069 12113 20103
rect 12113 20069 12147 20103
rect 12147 20069 12156 20103
rect 12104 20060 12156 20069
rect 20752 20060 20804 20112
rect 3510 19958 3562 20010
rect 3574 19958 3626 20010
rect 3638 19958 3690 20010
rect 3702 19958 3754 20010
rect 3766 19958 3818 20010
rect 1156 19899 1208 19908
rect 1156 19865 1165 19899
rect 1165 19865 1199 19899
rect 1199 19865 1208 19899
rect 1156 19856 1208 19865
rect 3180 19856 3232 19908
rect 6308 19856 6360 19908
rect 7228 19899 7280 19908
rect 7228 19865 7237 19899
rect 7237 19865 7271 19899
rect 7271 19865 7280 19899
rect 7228 19856 7280 19865
rect 9252 19899 9304 19908
rect 9252 19865 9261 19899
rect 9261 19865 9295 19899
rect 9295 19865 9304 19899
rect 9252 19856 9304 19865
rect 9804 19899 9856 19908
rect 9804 19865 9813 19899
rect 9813 19865 9847 19899
rect 9847 19865 9856 19899
rect 9804 19856 9856 19865
rect 10356 19856 10408 19908
rect 788 19788 840 19840
rect 7320 19788 7372 19840
rect 7872 19788 7924 19840
rect 9528 19788 9580 19840
rect 2628 19695 2680 19704
rect 2628 19661 2637 19695
rect 2637 19661 2671 19695
rect 2671 19661 2680 19695
rect 2628 19652 2680 19661
rect 2720 19652 2772 19704
rect 3364 19652 3416 19704
rect 6676 19652 6728 19704
rect 7412 19652 7464 19704
rect 8148 19695 8200 19746
rect 8148 19694 8157 19695
rect 8157 19694 8191 19695
rect 8191 19694 8200 19695
rect 3272 19584 3324 19636
rect 7136 19584 7188 19636
rect 10356 19720 10408 19772
rect 8516 19695 8568 19704
rect 8516 19661 8525 19695
rect 8525 19661 8559 19695
rect 8559 19661 8568 19695
rect 8516 19652 8568 19661
rect 9528 19652 9580 19704
rect 9988 19695 10040 19704
rect 9988 19661 9997 19695
rect 9997 19661 10031 19695
rect 10031 19661 10040 19695
rect 9988 19652 10040 19661
rect 10172 19695 10224 19704
rect 10172 19661 10181 19695
rect 10181 19661 10215 19695
rect 10215 19661 10224 19695
rect 10172 19652 10224 19661
rect 12012 19856 12064 19908
rect 12288 19856 12340 19908
rect 14680 19899 14732 19908
rect 14680 19865 14689 19899
rect 14689 19865 14723 19899
rect 14723 19865 14732 19899
rect 14680 19856 14732 19865
rect 14956 19856 15008 19908
rect 16520 19856 16572 19908
rect 18084 19856 18136 19908
rect 21856 19856 21908 19908
rect 11184 19831 11236 19840
rect 11184 19797 11193 19831
rect 11193 19797 11227 19831
rect 11227 19797 11236 19831
rect 11184 19788 11236 19797
rect 17808 19788 17860 19840
rect 18544 19788 18596 19840
rect 19924 19788 19976 19840
rect 21212 19788 21264 19840
rect 21672 19788 21724 19840
rect 11092 19695 11144 19704
rect 11092 19661 11101 19695
rect 11101 19661 11135 19695
rect 11135 19661 11144 19695
rect 11092 19652 11144 19661
rect 11736 19695 11788 19704
rect 11736 19661 11745 19695
rect 11745 19661 11779 19695
rect 11779 19661 11788 19695
rect 11736 19652 11788 19661
rect 20752 19763 20804 19772
rect 20752 19729 20761 19763
rect 20761 19729 20795 19763
rect 20795 19729 20804 19763
rect 20752 19720 20804 19729
rect 12104 19652 12156 19704
rect 12380 19652 12432 19704
rect 12840 19652 12892 19704
rect 20292 19652 20344 19704
rect 21212 19695 21264 19704
rect 21212 19661 21221 19695
rect 21221 19661 21255 19695
rect 21255 19661 21264 19695
rect 21212 19652 21264 19661
rect 24156 19856 24208 19908
rect 27192 19899 27244 19908
rect 27192 19865 27201 19899
rect 27201 19865 27235 19899
rect 27235 19865 27244 19899
rect 27192 19856 27244 19865
rect 28112 19856 28164 19908
rect 27376 19788 27428 19840
rect 28020 19831 28072 19840
rect 28020 19797 28029 19831
rect 28029 19797 28063 19831
rect 28063 19797 28072 19831
rect 28020 19788 28072 19797
rect 28572 19720 28624 19772
rect 12932 19584 12984 19636
rect 27928 19652 27980 19704
rect 22040 19584 22092 19636
rect 7872 19516 7924 19568
rect 8976 19559 9028 19568
rect 8976 19525 8985 19559
rect 8985 19525 9019 19559
rect 9019 19525 9028 19559
rect 8976 19516 9028 19525
rect 9528 19516 9580 19568
rect 10356 19516 10408 19568
rect 16428 19516 16480 19568
rect 18084 19516 18136 19568
rect 19832 19559 19884 19568
rect 19832 19525 19841 19559
rect 19841 19525 19875 19559
rect 19875 19525 19884 19559
rect 19832 19516 19884 19525
rect 20200 19516 20252 19568
rect 26732 19584 26784 19636
rect 27836 19584 27888 19636
rect 26456 19516 26508 19568
rect 27376 19559 27428 19568
rect 27376 19525 27385 19559
rect 27385 19525 27419 19559
rect 27419 19525 27428 19559
rect 27376 19516 27428 19525
rect 18870 19414 18922 19466
rect 18934 19414 18986 19466
rect 18998 19414 19050 19466
rect 19062 19414 19114 19466
rect 19126 19414 19178 19466
rect 1892 19312 1944 19364
rect 2628 19312 2680 19364
rect 7044 19355 7096 19364
rect 7044 19321 7053 19355
rect 7053 19321 7087 19355
rect 7087 19321 7096 19355
rect 7044 19312 7096 19321
rect 7596 19355 7648 19364
rect 7596 19321 7605 19355
rect 7605 19321 7639 19355
rect 7639 19321 7648 19355
rect 7596 19312 7648 19321
rect 8516 19312 8568 19364
rect 9068 19312 9120 19364
rect 10172 19312 10224 19364
rect 11644 19312 11696 19364
rect 11736 19312 11788 19364
rect 12288 19312 12340 19364
rect 2720 19244 2772 19296
rect 3272 19244 3324 19296
rect 5388 19244 5440 19296
rect 6492 19244 6544 19296
rect 7412 19244 7464 19296
rect 9988 19244 10040 19296
rect 12104 19244 12156 19296
rect 12748 19244 12800 19296
rect 3364 19219 3416 19228
rect 3364 19185 3373 19219
rect 3373 19185 3407 19219
rect 3407 19185 3416 19219
rect 3364 19176 3416 19185
rect 4836 19176 4888 19228
rect 6308 19219 6360 19228
rect 6308 19185 6317 19219
rect 6317 19185 6351 19219
rect 6351 19185 6360 19219
rect 7872 19219 7924 19228
rect 6308 19176 6360 19185
rect 7872 19185 7881 19219
rect 7881 19185 7915 19219
rect 7915 19185 7924 19219
rect 7872 19176 7924 19185
rect 10540 19219 10592 19228
rect 10540 19185 10549 19219
rect 10549 19185 10583 19219
rect 10583 19185 10592 19219
rect 10540 19176 10592 19185
rect 11552 19219 11604 19228
rect 11552 19185 11561 19219
rect 11561 19185 11595 19219
rect 11595 19185 11604 19219
rect 11552 19176 11604 19185
rect 12840 19176 12892 19228
rect 15232 19244 15284 19296
rect 17808 19312 17860 19364
rect 20292 19355 20344 19364
rect 20292 19321 20301 19355
rect 20301 19321 20335 19355
rect 20335 19321 20344 19355
rect 20292 19312 20344 19321
rect 20752 19312 20804 19364
rect 21396 19355 21448 19364
rect 21396 19321 21405 19355
rect 21405 19321 21439 19355
rect 21439 19321 21448 19355
rect 21396 19312 21448 19321
rect 23420 19312 23472 19364
rect 16888 19287 16940 19296
rect 16888 19253 16897 19287
rect 16897 19253 16931 19287
rect 16931 19253 16940 19287
rect 16888 19244 16940 19253
rect 28204 19244 28256 19296
rect 28664 19244 28716 19296
rect 29400 19244 29452 19296
rect 16152 19219 16204 19228
rect 16152 19185 16161 19219
rect 16161 19185 16195 19219
rect 16195 19185 16204 19219
rect 16152 19176 16204 19185
rect 16612 19219 16664 19228
rect 16612 19185 16621 19219
rect 16621 19185 16655 19219
rect 16655 19185 16664 19219
rect 16612 19176 16664 19185
rect 20660 19176 20712 19228
rect 22040 19176 22092 19228
rect 23236 19219 23288 19228
rect 23236 19185 23245 19219
rect 23245 19185 23279 19219
rect 23279 19185 23288 19219
rect 23236 19176 23288 19185
rect 26916 19176 26968 19228
rect 27928 19219 27980 19228
rect 27928 19185 27937 19219
rect 27937 19185 27971 19219
rect 27971 19185 27980 19219
rect 27928 19176 27980 19185
rect 29124 19219 29176 19228
rect 29124 19185 29133 19219
rect 29133 19185 29167 19219
rect 29167 19185 29176 19219
rect 29124 19176 29176 19185
rect 30504 19219 30556 19228
rect 30504 19185 30513 19219
rect 30513 19185 30547 19219
rect 30547 19185 30556 19219
rect 30504 19176 30556 19185
rect 5296 19151 5348 19160
rect 5296 19117 5305 19151
rect 5305 19117 5339 19151
rect 5339 19117 5348 19151
rect 5296 19108 5348 19117
rect 11736 19108 11788 19160
rect 13484 19151 13536 19160
rect 13484 19117 13493 19151
rect 13493 19117 13527 19151
rect 13527 19117 13536 19151
rect 13484 19108 13536 19117
rect 15048 19151 15100 19160
rect 15048 19117 15057 19151
rect 15057 19117 15091 19151
rect 15091 19117 15100 19151
rect 15048 19108 15100 19117
rect 22132 19151 22184 19160
rect 22132 19117 22141 19151
rect 22141 19117 22175 19151
rect 22175 19117 22184 19151
rect 22132 19108 22184 19117
rect 26732 19108 26784 19160
rect 27652 19151 27704 19160
rect 27652 19117 27661 19151
rect 27661 19117 27695 19151
rect 27695 19117 27704 19151
rect 27652 19108 27704 19117
rect 28112 19151 28164 19160
rect 28112 19117 28121 19151
rect 28121 19117 28155 19151
rect 28155 19117 28164 19151
rect 28112 19108 28164 19117
rect 29584 19108 29636 19160
rect 10264 19040 10316 19092
rect 10356 19015 10408 19024
rect 10356 18981 10365 19015
rect 10365 18981 10399 19015
rect 10399 18981 10408 19015
rect 10356 18972 10408 18981
rect 21028 18972 21080 19024
rect 24156 18972 24208 19024
rect 24708 18972 24760 19024
rect 25168 18972 25220 19024
rect 3510 18870 3562 18922
rect 3574 18870 3626 18922
rect 3638 18870 3690 18922
rect 3702 18870 3754 18922
rect 3766 18870 3818 18922
rect 3364 18811 3416 18820
rect 3364 18777 3373 18811
rect 3373 18777 3407 18811
rect 3407 18777 3416 18811
rect 3364 18768 3416 18777
rect 5296 18811 5348 18820
rect 5296 18777 5305 18811
rect 5305 18777 5339 18811
rect 5339 18777 5348 18811
rect 5296 18768 5348 18777
rect 6308 18811 6360 18820
rect 6308 18777 6317 18811
rect 6317 18777 6351 18811
rect 6351 18777 6360 18811
rect 6308 18768 6360 18777
rect 6492 18811 6544 18820
rect 6492 18777 6501 18811
rect 6501 18777 6535 18811
rect 6535 18777 6544 18811
rect 6492 18768 6544 18777
rect 10540 18768 10592 18820
rect 11276 18811 11328 18820
rect 11276 18777 11285 18811
rect 11285 18777 11319 18811
rect 11319 18777 11328 18811
rect 11276 18768 11328 18777
rect 11552 18811 11604 18820
rect 11552 18777 11561 18811
rect 11561 18777 11595 18811
rect 11595 18777 11604 18811
rect 11552 18768 11604 18777
rect 12104 18768 12156 18820
rect 12748 18768 12800 18820
rect 13484 18768 13536 18820
rect 3272 18700 3324 18752
rect 9804 18700 9856 18752
rect 5480 18632 5532 18684
rect 8976 18632 9028 18684
rect 11276 18632 11328 18684
rect 12840 18632 12892 18684
rect 6676 18564 6728 18616
rect 10356 18564 10408 18616
rect 12104 18564 12156 18616
rect 13116 18564 13168 18616
rect 1616 18428 1668 18480
rect 5940 18496 5992 18548
rect 13668 18539 13720 18548
rect 13668 18505 13677 18539
rect 13677 18505 13711 18539
rect 13711 18505 13720 18539
rect 13668 18496 13720 18505
rect 4836 18428 4888 18480
rect 13944 18632 13996 18684
rect 15048 18768 15100 18820
rect 15232 18768 15284 18820
rect 16152 18811 16204 18820
rect 16152 18777 16161 18811
rect 16161 18777 16195 18811
rect 16195 18777 16204 18811
rect 16152 18768 16204 18777
rect 16888 18768 16940 18820
rect 23236 18811 23288 18820
rect 23236 18777 23245 18811
rect 23245 18777 23279 18811
rect 23279 18777 23288 18811
rect 23236 18768 23288 18777
rect 23512 18811 23564 18820
rect 23512 18777 23521 18811
rect 23521 18777 23555 18811
rect 23555 18777 23564 18811
rect 25904 18811 25956 18820
rect 23512 18768 23564 18777
rect 25904 18777 25913 18811
rect 25913 18777 25947 18811
rect 25947 18777 25956 18811
rect 25904 18768 25956 18777
rect 26732 18811 26784 18820
rect 26732 18777 26741 18811
rect 26741 18777 26775 18811
rect 26775 18777 26784 18811
rect 26732 18768 26784 18777
rect 26916 18811 26968 18820
rect 26916 18777 26925 18811
rect 26925 18777 26959 18811
rect 26959 18777 26968 18811
rect 26916 18768 26968 18777
rect 28112 18768 28164 18820
rect 29124 18768 29176 18820
rect 29492 18768 29544 18820
rect 29584 18768 29636 18820
rect 30504 18768 30556 18820
rect 14680 18700 14732 18752
rect 15232 18564 15284 18616
rect 16704 18564 16756 18616
rect 23420 18700 23472 18752
rect 27652 18743 27704 18752
rect 27652 18709 27661 18743
rect 27661 18709 27695 18743
rect 27695 18709 27704 18743
rect 27652 18700 27704 18709
rect 28204 18700 28256 18752
rect 24156 18675 24208 18684
rect 22040 18607 22092 18616
rect 22040 18573 22049 18607
rect 22049 18573 22083 18607
rect 22083 18573 22092 18607
rect 22040 18564 22092 18573
rect 23788 18607 23840 18616
rect 23788 18573 23797 18607
rect 23797 18573 23831 18607
rect 23831 18573 23840 18607
rect 23788 18564 23840 18573
rect 24156 18641 24165 18675
rect 24165 18641 24199 18675
rect 24199 18641 24208 18675
rect 24156 18632 24208 18641
rect 29032 18700 29084 18752
rect 29400 18632 29452 18684
rect 14588 18428 14640 18480
rect 16612 18428 16664 18480
rect 17072 18428 17124 18480
rect 22132 18471 22184 18480
rect 22132 18437 22141 18471
rect 22141 18437 22175 18471
rect 22175 18437 22184 18471
rect 22132 18428 22184 18437
rect 23696 18471 23748 18480
rect 23696 18437 23705 18471
rect 23705 18437 23739 18471
rect 23739 18437 23748 18471
rect 23696 18428 23748 18437
rect 24708 18496 24760 18548
rect 27744 18564 27796 18616
rect 28204 18564 28256 18616
rect 26640 18496 26692 18548
rect 28112 18471 28164 18480
rect 28112 18437 28121 18471
rect 28121 18437 28155 18471
rect 28155 18437 28164 18471
rect 28112 18428 28164 18437
rect 29400 18471 29452 18480
rect 29400 18437 29409 18471
rect 29409 18437 29443 18471
rect 29443 18437 29452 18471
rect 29400 18428 29452 18437
rect 18870 18326 18922 18378
rect 18934 18326 18986 18378
rect 18998 18326 19050 18378
rect 19062 18326 19114 18378
rect 19126 18326 19178 18378
rect 4008 18224 4060 18276
rect 6124 18224 6176 18276
rect 4376 18156 4428 18208
rect 6952 18156 7004 18208
rect 14588 18199 14640 18208
rect 14588 18165 14597 18199
rect 14597 18165 14631 18199
rect 14631 18165 14640 18199
rect 14588 18156 14640 18165
rect 16152 18156 16204 18208
rect 21120 18156 21172 18208
rect 26640 18199 26692 18208
rect 26640 18165 26649 18199
rect 26649 18165 26683 18199
rect 26683 18165 26692 18199
rect 26640 18156 26692 18165
rect 28388 18156 28440 18208
rect 28756 18156 28808 18208
rect 4744 18088 4796 18140
rect 6492 18088 6544 18140
rect 7320 18088 7372 18140
rect 12748 18088 12800 18140
rect 12932 18131 12984 18140
rect 12932 18097 12941 18131
rect 12941 18097 12975 18131
rect 12975 18097 12984 18131
rect 13116 18131 13168 18140
rect 12932 18088 12984 18097
rect 13116 18097 13125 18131
rect 13125 18097 13159 18131
rect 13159 18097 13168 18131
rect 13116 18088 13168 18097
rect 14772 18131 14824 18140
rect 14772 18097 14781 18131
rect 14781 18097 14815 18131
rect 14815 18097 14824 18131
rect 14772 18088 14824 18097
rect 15232 18088 15284 18140
rect 16612 18131 16664 18140
rect 16612 18097 16621 18131
rect 16621 18097 16655 18131
rect 16655 18097 16664 18131
rect 16612 18088 16664 18097
rect 17072 18131 17124 18140
rect 17072 18097 17081 18131
rect 17081 18097 17115 18131
rect 17115 18097 17124 18131
rect 17072 18088 17124 18097
rect 17440 18088 17492 18140
rect 26456 18088 26508 18140
rect 28020 18131 28072 18140
rect 28020 18097 28029 18131
rect 28029 18097 28063 18131
rect 28063 18097 28072 18131
rect 28020 18088 28072 18097
rect 5480 18020 5532 18072
rect 6676 18020 6728 18072
rect 13576 18063 13628 18072
rect 13576 18029 13585 18063
rect 13585 18029 13619 18063
rect 13619 18029 13628 18063
rect 17164 18063 17216 18072
rect 13576 18020 13628 18029
rect 17164 18029 17173 18063
rect 17173 18029 17207 18063
rect 17207 18029 17216 18063
rect 17164 18020 17216 18029
rect 17808 18020 17860 18072
rect 20752 18063 20804 18072
rect 20752 18029 20761 18063
rect 20761 18029 20795 18063
rect 20795 18029 20804 18063
rect 20752 18020 20804 18029
rect 21672 18020 21724 18072
rect 30044 18063 30096 18072
rect 30044 18029 30053 18063
rect 30053 18029 30087 18063
rect 30087 18029 30096 18063
rect 30044 18020 30096 18029
rect 5388 17952 5440 18004
rect 6308 17952 6360 18004
rect 5296 17927 5348 17936
rect 5296 17893 5305 17927
rect 5305 17893 5339 17927
rect 5339 17893 5348 17927
rect 5296 17884 5348 17893
rect 6768 17884 6820 17936
rect 7228 17884 7280 17936
rect 18176 17884 18228 17936
rect 19832 17884 19884 17936
rect 20936 17884 20988 17936
rect 23420 17884 23472 17936
rect 23788 17927 23840 17936
rect 23788 17893 23797 17927
rect 23797 17893 23831 17927
rect 23831 17893 23840 17927
rect 23788 17884 23840 17893
rect 23972 17884 24024 17936
rect 24248 17884 24300 17936
rect 26916 17927 26968 17936
rect 26916 17893 26925 17927
rect 26925 17893 26959 17927
rect 26959 17893 26968 17927
rect 26916 17884 26968 17893
rect 3510 17782 3562 17834
rect 3574 17782 3626 17834
rect 3638 17782 3690 17834
rect 3702 17782 3754 17834
rect 3766 17782 3818 17834
rect 2352 17476 2404 17528
rect 5296 17680 5348 17732
rect 6492 17723 6544 17732
rect 6492 17689 6501 17723
rect 6501 17689 6535 17723
rect 6535 17689 6544 17723
rect 6492 17680 6544 17689
rect 6676 17723 6728 17732
rect 6676 17689 6685 17723
rect 6685 17689 6719 17723
rect 6719 17689 6728 17723
rect 6676 17680 6728 17689
rect 6768 17723 6820 17732
rect 6768 17689 6777 17723
rect 6777 17689 6811 17723
rect 6811 17689 6820 17723
rect 6952 17723 7004 17732
rect 6768 17680 6820 17689
rect 6952 17689 6961 17723
rect 6961 17689 6995 17723
rect 6995 17689 7004 17723
rect 6952 17680 7004 17689
rect 4744 17612 4796 17664
rect 1616 17451 1668 17460
rect 1616 17417 1625 17451
rect 1625 17417 1659 17451
rect 1659 17417 1668 17451
rect 1616 17408 1668 17417
rect 1248 17340 1300 17392
rect 1800 17340 1852 17392
rect 2352 17383 2404 17392
rect 2352 17349 2361 17383
rect 2361 17349 2395 17383
rect 2395 17349 2404 17383
rect 2352 17340 2404 17349
rect 3916 17340 3968 17392
rect 4468 17408 4520 17460
rect 4560 17408 4612 17460
rect 11552 17680 11604 17732
rect 12748 17723 12800 17732
rect 12748 17689 12757 17723
rect 12757 17689 12791 17723
rect 12791 17689 12800 17723
rect 12748 17680 12800 17689
rect 13024 17680 13076 17732
rect 4836 17408 4888 17460
rect 5204 17340 5256 17392
rect 5480 17476 5532 17528
rect 8424 17519 8476 17528
rect 8424 17485 8433 17519
rect 8433 17485 8467 17519
rect 8467 17485 8476 17519
rect 11920 17612 11972 17664
rect 12932 17612 12984 17664
rect 13668 17680 13720 17732
rect 14772 17680 14824 17732
rect 17164 17680 17216 17732
rect 20200 17680 20252 17732
rect 20752 17680 20804 17732
rect 20844 17680 20896 17732
rect 22132 17680 22184 17732
rect 23880 17680 23932 17732
rect 26916 17680 26968 17732
rect 30044 17680 30096 17732
rect 14588 17612 14640 17664
rect 19924 17655 19976 17664
rect 19924 17621 19933 17655
rect 19933 17621 19967 17655
rect 19967 17621 19976 17655
rect 19924 17612 19976 17621
rect 21672 17612 21724 17664
rect 26456 17612 26508 17664
rect 28020 17612 28072 17664
rect 18176 17587 18228 17596
rect 8424 17476 8476 17485
rect 12748 17476 12800 17528
rect 13668 17476 13720 17528
rect 18176 17553 18185 17587
rect 18185 17553 18219 17587
rect 18219 17553 18228 17587
rect 18176 17544 18228 17553
rect 23972 17587 24024 17596
rect 23972 17553 23981 17587
rect 23981 17553 24015 17587
rect 24015 17553 24024 17587
rect 23972 17544 24024 17553
rect 24248 17544 24300 17596
rect 25536 17544 25588 17596
rect 26640 17544 26692 17596
rect 28388 17544 28440 17596
rect 17808 17519 17860 17528
rect 17808 17485 17817 17519
rect 17817 17485 17851 17519
rect 17851 17485 17860 17519
rect 17808 17476 17860 17485
rect 20844 17519 20896 17528
rect 20844 17485 20853 17519
rect 20853 17485 20887 17519
rect 20887 17485 20896 17519
rect 20844 17476 20896 17485
rect 20936 17519 20988 17528
rect 20936 17485 20945 17519
rect 20945 17485 20979 17519
rect 20979 17485 20988 17519
rect 20936 17476 20988 17485
rect 22500 17476 22552 17528
rect 25904 17476 25956 17528
rect 9068 17408 9120 17460
rect 13760 17451 13812 17460
rect 13760 17417 13769 17451
rect 13769 17417 13803 17451
rect 13803 17417 13812 17451
rect 13760 17408 13812 17417
rect 14588 17451 14640 17460
rect 14588 17417 14597 17451
rect 14597 17417 14631 17451
rect 14631 17417 14640 17451
rect 14588 17408 14640 17417
rect 16428 17408 16480 17460
rect 17072 17408 17124 17460
rect 20108 17451 20160 17460
rect 7228 17383 7280 17392
rect 7228 17349 7237 17383
rect 7237 17349 7271 17383
rect 7271 17349 7280 17383
rect 7228 17340 7280 17349
rect 14128 17383 14180 17392
rect 14128 17349 14137 17383
rect 14137 17349 14171 17383
rect 14171 17349 14180 17383
rect 14128 17340 14180 17349
rect 14312 17340 14364 17392
rect 15968 17340 16020 17392
rect 16060 17340 16112 17392
rect 16612 17383 16664 17392
rect 16612 17349 16621 17383
rect 16621 17349 16655 17383
rect 16655 17349 16664 17383
rect 16612 17340 16664 17349
rect 17532 17383 17584 17392
rect 17532 17349 17541 17383
rect 17541 17349 17575 17383
rect 17575 17349 17584 17383
rect 17532 17340 17584 17349
rect 20108 17417 20117 17451
rect 20117 17417 20151 17451
rect 20151 17417 20160 17451
rect 21396 17451 21448 17460
rect 20108 17408 20160 17417
rect 21396 17417 21405 17451
rect 21405 17417 21439 17451
rect 21439 17417 21448 17451
rect 21396 17408 21448 17417
rect 22592 17408 22644 17460
rect 23696 17408 23748 17460
rect 20200 17340 20252 17392
rect 21120 17340 21172 17392
rect 21856 17383 21908 17392
rect 21856 17349 21865 17383
rect 21865 17349 21899 17383
rect 21899 17349 21908 17383
rect 23420 17383 23472 17392
rect 21856 17340 21908 17349
rect 23420 17349 23429 17383
rect 23429 17349 23463 17383
rect 23463 17349 23472 17383
rect 23420 17340 23472 17349
rect 23604 17383 23656 17392
rect 23604 17349 23613 17383
rect 23613 17349 23647 17383
rect 23647 17349 23656 17383
rect 23604 17340 23656 17349
rect 24708 17408 24760 17460
rect 28480 17408 28532 17460
rect 27192 17383 27244 17392
rect 27192 17349 27201 17383
rect 27201 17349 27235 17383
rect 27235 17349 27244 17383
rect 27192 17340 27244 17349
rect 28572 17383 28624 17392
rect 28572 17349 28581 17383
rect 28581 17349 28615 17383
rect 28615 17349 28624 17383
rect 28572 17340 28624 17349
rect 18870 17238 18922 17290
rect 18934 17238 18986 17290
rect 18998 17238 19050 17290
rect 19062 17238 19114 17290
rect 19126 17238 19178 17290
rect 1248 17179 1300 17188
rect 1248 17145 1257 17179
rect 1257 17145 1291 17179
rect 1291 17145 1300 17179
rect 1248 17136 1300 17145
rect 4744 17136 4796 17188
rect 1616 17043 1668 17052
rect 1616 17009 1625 17043
rect 1625 17009 1659 17043
rect 1659 17009 1668 17043
rect 1616 17000 1668 17009
rect 2352 17000 2404 17052
rect 4284 17000 4336 17052
rect 4468 17000 4520 17052
rect 5204 17043 5256 17052
rect 5204 17009 5213 17043
rect 5213 17009 5247 17043
rect 5247 17009 5256 17043
rect 5204 17000 5256 17009
rect 5388 17000 5440 17052
rect 5480 17043 5532 17052
rect 5480 17009 5489 17043
rect 5489 17009 5523 17043
rect 5523 17009 5532 17043
rect 13576 17136 13628 17188
rect 14128 17136 14180 17188
rect 15232 17136 15284 17188
rect 18176 17179 18228 17188
rect 18176 17145 18185 17179
rect 18185 17145 18219 17179
rect 18219 17145 18228 17179
rect 18176 17136 18228 17145
rect 20752 17136 20804 17188
rect 27192 17136 27244 17188
rect 12748 17068 12800 17120
rect 14956 17068 15008 17120
rect 5480 17000 5532 17009
rect 7412 17000 7464 17052
rect 9068 17043 9120 17052
rect 9068 17009 9077 17043
rect 9077 17009 9111 17043
rect 9111 17009 9120 17043
rect 9068 17000 9120 17009
rect 9160 17000 9212 17052
rect 11276 17000 11328 17052
rect 12932 17000 12984 17052
rect 15968 17043 16020 17052
rect 15968 17009 15977 17043
rect 15977 17009 16011 17043
rect 16011 17009 16020 17043
rect 15968 17000 16020 17009
rect 16428 17043 16480 17052
rect 16428 17009 16437 17043
rect 16437 17009 16471 17043
rect 16471 17009 16480 17043
rect 16428 17000 16480 17009
rect 17716 17000 17768 17052
rect 19556 17068 19608 17120
rect 27836 17111 27888 17120
rect 18820 17000 18872 17052
rect 20108 17000 20160 17052
rect 27836 17077 27845 17111
rect 27845 17077 27879 17111
rect 27879 17077 27888 17111
rect 27836 17068 27888 17077
rect 20936 17000 20988 17052
rect 21396 17000 21448 17052
rect 22960 17043 23012 17052
rect 22960 17009 22969 17043
rect 22969 17009 23003 17043
rect 23003 17009 23012 17043
rect 22960 17000 23012 17009
rect 23328 17043 23380 17052
rect 23328 17009 23337 17043
rect 23337 17009 23371 17043
rect 23371 17009 23380 17043
rect 23328 17000 23380 17009
rect 27744 17043 27796 17052
rect 27744 17009 27753 17043
rect 27753 17009 27787 17043
rect 27787 17009 27796 17043
rect 27744 17000 27796 17009
rect 28020 17000 28072 17052
rect 1708 16975 1760 16984
rect 1708 16941 1717 16975
rect 1717 16941 1751 16975
rect 1751 16941 1760 16975
rect 1708 16932 1760 16941
rect 3916 16975 3968 16984
rect 3916 16941 3925 16975
rect 3925 16941 3959 16975
rect 3959 16941 3968 16975
rect 3916 16932 3968 16941
rect 4100 16932 4152 16984
rect 4376 16975 4428 16984
rect 4376 16941 4385 16975
rect 4385 16941 4419 16975
rect 4419 16941 4428 16975
rect 4376 16932 4428 16941
rect 5756 16975 5808 16984
rect 5756 16941 5765 16975
rect 5765 16941 5799 16975
rect 5799 16941 5808 16975
rect 5756 16932 5808 16941
rect 6768 16975 6820 16984
rect 6768 16941 6777 16975
rect 6777 16941 6811 16975
rect 6811 16941 6820 16975
rect 6768 16932 6820 16941
rect 7136 16932 7188 16984
rect 7596 16932 7648 16984
rect 9804 16975 9856 16984
rect 9804 16941 9813 16975
rect 9813 16941 9847 16975
rect 9847 16941 9856 16975
rect 9804 16932 9856 16941
rect 16520 16975 16572 16984
rect 16520 16941 16529 16975
rect 16529 16941 16563 16975
rect 16563 16941 16572 16975
rect 16520 16932 16572 16941
rect 18544 16975 18596 16984
rect 18544 16941 18553 16975
rect 18553 16941 18587 16975
rect 18587 16941 18596 16975
rect 18544 16932 18596 16941
rect 19004 16975 19056 16984
rect 19004 16941 19013 16975
rect 19013 16941 19047 16975
rect 19047 16941 19056 16975
rect 19004 16932 19056 16941
rect 19924 16932 19976 16984
rect 20476 16932 20528 16984
rect 4468 16864 4520 16916
rect 9528 16864 9580 16916
rect 17808 16907 17860 16916
rect 17808 16873 17817 16907
rect 17817 16873 17851 16907
rect 17851 16873 17860 16907
rect 17808 16864 17860 16873
rect 20292 16864 20344 16916
rect 21672 16932 21724 16984
rect 22500 16932 22552 16984
rect 23144 16932 23196 16984
rect 23236 16864 23288 16916
rect 2536 16796 2588 16848
rect 9712 16796 9764 16848
rect 14772 16839 14824 16848
rect 14772 16805 14781 16839
rect 14781 16805 14815 16839
rect 14815 16805 14824 16839
rect 14772 16796 14824 16805
rect 17716 16796 17768 16848
rect 19372 16839 19424 16848
rect 19372 16805 19381 16839
rect 19381 16805 19415 16839
rect 19415 16805 19424 16839
rect 19372 16796 19424 16805
rect 24064 16839 24116 16848
rect 24064 16805 24073 16839
rect 24073 16805 24107 16839
rect 24107 16805 24116 16839
rect 24064 16796 24116 16805
rect 27928 16796 27980 16848
rect 3510 16694 3562 16746
rect 3574 16694 3626 16746
rect 3638 16694 3690 16746
rect 3702 16694 3754 16746
rect 3766 16694 3818 16746
rect 3916 16635 3968 16644
rect 3916 16601 3925 16635
rect 3925 16601 3959 16635
rect 3959 16601 3968 16635
rect 3916 16592 3968 16601
rect 4100 16635 4152 16644
rect 4100 16601 4109 16635
rect 4109 16601 4143 16635
rect 4143 16601 4152 16635
rect 4100 16592 4152 16601
rect 4284 16635 4336 16644
rect 4284 16601 4293 16635
rect 4293 16601 4327 16635
rect 4327 16601 4336 16635
rect 4284 16592 4336 16601
rect 4468 16635 4520 16644
rect 4468 16601 4477 16635
rect 4477 16601 4511 16635
rect 4511 16601 4520 16635
rect 4468 16592 4520 16601
rect 5204 16635 5256 16644
rect 5204 16601 5213 16635
rect 5213 16601 5247 16635
rect 5247 16601 5256 16635
rect 5204 16592 5256 16601
rect 5388 16592 5440 16644
rect 5756 16635 5808 16644
rect 5756 16601 5765 16635
rect 5765 16601 5799 16635
rect 5799 16601 5808 16635
rect 5756 16592 5808 16601
rect 7412 16635 7464 16644
rect 7412 16601 7421 16635
rect 7421 16601 7455 16635
rect 7455 16601 7464 16635
rect 7412 16592 7464 16601
rect 7596 16635 7648 16644
rect 7596 16601 7605 16635
rect 7605 16601 7639 16635
rect 7639 16601 7648 16635
rect 7596 16592 7648 16601
rect 14956 16592 15008 16644
rect 15968 16635 16020 16644
rect 15968 16601 15977 16635
rect 15977 16601 16011 16635
rect 16011 16601 16020 16635
rect 15968 16592 16020 16601
rect 16520 16592 16572 16644
rect 18176 16592 18228 16644
rect 20292 16635 20344 16644
rect 20292 16601 20301 16635
rect 20301 16601 20335 16635
rect 20335 16601 20344 16635
rect 20292 16592 20344 16601
rect 20752 16592 20804 16644
rect 21396 16592 21448 16644
rect 22500 16635 22552 16644
rect 22500 16601 22509 16635
rect 22509 16601 22543 16635
rect 22543 16601 22552 16635
rect 22500 16592 22552 16601
rect 23236 16635 23288 16644
rect 23236 16601 23245 16635
rect 23245 16601 23279 16635
rect 23279 16601 23288 16635
rect 23236 16592 23288 16601
rect 24156 16592 24208 16644
rect 26916 16635 26968 16644
rect 26916 16601 26925 16635
rect 26925 16601 26959 16635
rect 26959 16601 26968 16635
rect 26916 16592 26968 16601
rect 27836 16635 27888 16644
rect 27836 16601 27845 16635
rect 27845 16601 27879 16635
rect 27879 16601 27888 16635
rect 27836 16592 27888 16601
rect 27928 16592 27980 16644
rect 1800 16431 1852 16440
rect 1800 16397 1809 16431
rect 1809 16397 1843 16431
rect 1843 16397 1852 16431
rect 1800 16388 1852 16397
rect 1892 16388 1944 16440
rect 2536 16431 2588 16440
rect 2536 16397 2545 16431
rect 2545 16397 2579 16431
rect 2579 16397 2588 16431
rect 2536 16388 2588 16397
rect 972 16295 1024 16304
rect 972 16261 981 16295
rect 981 16261 1015 16295
rect 1015 16261 1024 16295
rect 1708 16320 1760 16372
rect 5480 16567 5532 16576
rect 5480 16533 5489 16567
rect 5489 16533 5523 16567
rect 5523 16533 5532 16567
rect 5480 16524 5532 16533
rect 3272 16388 3324 16440
rect 4376 16456 4428 16508
rect 11736 16524 11788 16576
rect 6860 16456 6912 16508
rect 4284 16388 4336 16440
rect 7228 16431 7280 16440
rect 7228 16397 7237 16431
rect 7237 16397 7271 16431
rect 7271 16397 7280 16431
rect 7228 16388 7280 16397
rect 8240 16456 8292 16508
rect 8424 16431 8476 16440
rect 8424 16397 8433 16431
rect 8433 16397 8467 16431
rect 8467 16397 8476 16431
rect 8424 16388 8476 16397
rect 9712 16388 9764 16440
rect 13944 16456 13996 16508
rect 16428 16456 16480 16508
rect 17532 16524 17584 16576
rect 19004 16524 19056 16576
rect 20936 16567 20988 16576
rect 20936 16533 20945 16567
rect 20945 16533 20979 16567
rect 20979 16533 20988 16567
rect 20936 16524 20988 16533
rect 23512 16524 23564 16576
rect 19280 16499 19332 16508
rect 19280 16465 19289 16499
rect 19289 16465 19323 16499
rect 19323 16465 19332 16499
rect 19280 16456 19332 16465
rect 23328 16456 23380 16508
rect 24064 16524 24116 16576
rect 11736 16431 11788 16440
rect 11736 16397 11745 16431
rect 11745 16397 11779 16431
rect 11779 16397 11788 16431
rect 11736 16388 11788 16397
rect 12564 16388 12616 16440
rect 17440 16431 17492 16440
rect 17440 16397 17449 16431
rect 17449 16397 17483 16431
rect 17483 16397 17492 16431
rect 17440 16388 17492 16397
rect 17716 16431 17768 16440
rect 17716 16397 17725 16431
rect 17725 16397 17759 16431
rect 17759 16397 17768 16431
rect 17716 16388 17768 16397
rect 19372 16431 19424 16440
rect 19372 16397 19381 16431
rect 19381 16397 19415 16431
rect 19415 16397 19424 16431
rect 19372 16388 19424 16397
rect 3364 16320 3416 16372
rect 7320 16363 7372 16372
rect 7320 16329 7329 16363
rect 7329 16329 7363 16363
rect 7363 16329 7372 16363
rect 7320 16320 7372 16329
rect 7964 16320 8016 16372
rect 12104 16363 12156 16372
rect 12104 16329 12113 16363
rect 12113 16329 12147 16363
rect 12147 16329 12156 16363
rect 12104 16320 12156 16329
rect 19464 16320 19516 16372
rect 6768 16295 6820 16304
rect 972 16252 1024 16261
rect 6768 16261 6777 16295
rect 6777 16261 6811 16295
rect 6811 16261 6820 16295
rect 6768 16252 6820 16261
rect 10540 16252 10592 16304
rect 14772 16252 14824 16304
rect 18452 16252 18504 16304
rect 19832 16431 19884 16440
rect 19832 16397 19841 16431
rect 19841 16397 19875 16431
rect 19875 16397 19884 16431
rect 19832 16388 19884 16397
rect 21580 16320 21632 16372
rect 23144 16388 23196 16440
rect 24156 16388 24208 16440
rect 24616 16431 24668 16440
rect 24616 16397 24625 16431
rect 24625 16397 24659 16431
rect 24659 16397 24668 16431
rect 24616 16388 24668 16397
rect 26180 16456 26232 16508
rect 27744 16567 27796 16576
rect 27744 16533 27753 16567
rect 27753 16533 27787 16567
rect 27787 16533 27796 16567
rect 27744 16524 27796 16533
rect 25260 16388 25312 16440
rect 25444 16388 25496 16440
rect 22960 16320 23012 16372
rect 20476 16252 20528 16304
rect 26180 16320 26232 16372
rect 30044 16388 30096 16440
rect 28020 16295 28072 16304
rect 28020 16261 28029 16295
rect 28029 16261 28063 16295
rect 28063 16261 28072 16295
rect 28020 16252 28072 16261
rect 29952 16295 30004 16304
rect 29952 16261 29961 16295
rect 29961 16261 29995 16295
rect 29995 16261 30004 16295
rect 29952 16252 30004 16261
rect 18870 16150 18922 16202
rect 18934 16150 18986 16202
rect 18998 16150 19050 16202
rect 19062 16150 19114 16202
rect 19126 16150 19178 16202
rect 1708 16091 1760 16100
rect 1708 16057 1717 16091
rect 1717 16057 1751 16091
rect 1751 16057 1760 16091
rect 1708 16048 1760 16057
rect 7320 16048 7372 16100
rect 9804 16048 9856 16100
rect 18728 16048 18780 16100
rect 19280 16091 19332 16100
rect 19280 16057 19289 16091
rect 19289 16057 19323 16091
rect 19323 16057 19332 16091
rect 19280 16048 19332 16057
rect 22132 16048 22184 16100
rect 1616 16023 1668 16032
rect 1616 15989 1625 16023
rect 1625 15989 1659 16023
rect 1659 15989 1668 16023
rect 1616 15980 1668 15989
rect 6768 15980 6820 16032
rect 1156 15955 1208 15964
rect 1156 15921 1165 15955
rect 1165 15921 1199 15955
rect 1199 15921 1208 15955
rect 1156 15912 1208 15921
rect 1984 15955 2036 15964
rect 1984 15921 1993 15955
rect 1993 15921 2027 15955
rect 2027 15921 2036 15955
rect 1984 15912 2036 15921
rect 3272 15912 3324 15964
rect 4008 15912 4060 15964
rect 5756 15912 5808 15964
rect 6308 15955 6360 15964
rect 2260 15887 2312 15896
rect 2260 15853 2269 15887
rect 2269 15853 2303 15887
rect 2303 15853 2312 15887
rect 2260 15844 2312 15853
rect 5848 15887 5900 15896
rect 5848 15853 5857 15887
rect 5857 15853 5891 15887
rect 5891 15853 5900 15887
rect 5848 15844 5900 15853
rect 6308 15921 6317 15955
rect 6317 15921 6351 15955
rect 6351 15921 6360 15955
rect 6308 15912 6360 15921
rect 6492 15955 6544 15964
rect 6492 15921 6501 15955
rect 6501 15921 6535 15955
rect 6535 15921 6544 15955
rect 8240 15980 8292 16032
rect 8424 16023 8476 16032
rect 8424 15989 8433 16023
rect 8433 15989 8467 16023
rect 8467 15989 8476 16023
rect 8424 15980 8476 15989
rect 8792 15980 8844 16032
rect 9160 15980 9212 16032
rect 12564 15980 12616 16032
rect 13760 15980 13812 16032
rect 6492 15912 6544 15921
rect 7688 15912 7740 15964
rect 10724 15955 10776 15964
rect 6952 15844 7004 15896
rect 7412 15844 7464 15896
rect 7044 15776 7096 15828
rect 10724 15921 10733 15955
rect 10733 15921 10767 15955
rect 10767 15921 10776 15955
rect 10724 15912 10776 15921
rect 11000 15912 11052 15964
rect 12104 15955 12156 15964
rect 12104 15921 12113 15955
rect 12113 15921 12147 15955
rect 12147 15921 12156 15955
rect 12104 15912 12156 15921
rect 15232 15980 15284 16032
rect 15600 15912 15652 15964
rect 15968 15980 16020 16032
rect 17440 15980 17492 16032
rect 17716 15980 17768 16032
rect 22592 15980 22644 16032
rect 24064 16048 24116 16100
rect 26732 16091 26784 16100
rect 26732 16057 26741 16091
rect 26741 16057 26775 16091
rect 26775 16057 26784 16091
rect 26732 16048 26784 16057
rect 27284 16048 27336 16100
rect 25444 15980 25496 16032
rect 27560 16023 27612 16032
rect 27560 15989 27569 16023
rect 27569 15989 27603 16023
rect 27603 15989 27612 16023
rect 27560 15980 27612 15989
rect 19464 15955 19516 15964
rect 19464 15921 19473 15955
rect 19473 15921 19507 15955
rect 19507 15921 19516 15955
rect 19464 15912 19516 15921
rect 22316 15912 22368 15964
rect 23880 15912 23932 15964
rect 25812 15912 25864 15964
rect 28204 15955 28256 15964
rect 28204 15921 28213 15955
rect 28213 15921 28247 15955
rect 28247 15921 28256 15955
rect 28204 15912 28256 15921
rect 28480 15912 28532 15964
rect 12288 15844 12340 15896
rect 18544 15844 18596 15896
rect 19832 15844 19884 15896
rect 21856 15887 21908 15896
rect 21856 15853 21865 15887
rect 21865 15853 21899 15887
rect 21899 15853 21908 15887
rect 21856 15844 21908 15853
rect 22224 15887 22276 15896
rect 22224 15853 22233 15887
rect 22233 15853 22267 15887
rect 22267 15853 22276 15887
rect 22224 15844 22276 15853
rect 28112 15887 28164 15896
rect 28112 15853 28121 15887
rect 28121 15853 28155 15887
rect 28155 15853 28164 15887
rect 28112 15844 28164 15853
rect 28388 15844 28440 15896
rect 8332 15776 8384 15828
rect 9068 15776 9120 15828
rect 24616 15776 24668 15828
rect 3364 15708 3416 15760
rect 4744 15751 4796 15760
rect 4744 15717 4753 15751
rect 4753 15717 4787 15751
rect 4787 15717 4796 15751
rect 4744 15708 4796 15717
rect 5388 15751 5440 15760
rect 5388 15717 5397 15751
rect 5397 15717 5431 15751
rect 5431 15717 5440 15751
rect 5388 15708 5440 15717
rect 9528 15751 9580 15760
rect 9528 15717 9537 15751
rect 9537 15717 9571 15751
rect 9571 15717 9580 15751
rect 9528 15708 9580 15717
rect 11000 15751 11052 15760
rect 11000 15717 11009 15751
rect 11009 15717 11043 15751
rect 11043 15717 11052 15751
rect 11000 15708 11052 15717
rect 18912 15751 18964 15760
rect 18912 15717 18921 15751
rect 18921 15717 18955 15751
rect 18955 15717 18964 15751
rect 18912 15708 18964 15717
rect 19004 15708 19056 15760
rect 21856 15708 21908 15760
rect 22408 15708 22460 15760
rect 24064 15751 24116 15760
rect 24064 15717 24073 15751
rect 24073 15717 24107 15751
rect 24107 15717 24116 15751
rect 26548 15751 26600 15760
rect 24064 15708 24116 15717
rect 26548 15717 26557 15751
rect 26557 15717 26591 15751
rect 26591 15717 26600 15751
rect 26548 15708 26600 15717
rect 3510 15606 3562 15658
rect 3574 15606 3626 15658
rect 3638 15606 3690 15658
rect 3702 15606 3754 15658
rect 3766 15606 3818 15658
rect 1156 15504 1208 15556
rect 1984 15547 2036 15556
rect 1984 15513 1993 15547
rect 1993 15513 2027 15547
rect 2027 15513 2036 15547
rect 1984 15504 2036 15513
rect 4468 15504 4520 15556
rect 4744 15504 4796 15556
rect 5756 15547 5808 15556
rect 5756 15513 5765 15547
rect 5765 15513 5799 15547
rect 5799 15513 5808 15547
rect 5756 15504 5808 15513
rect 6492 15504 6544 15556
rect 6952 15547 7004 15556
rect 6952 15513 6961 15547
rect 6961 15513 6995 15547
rect 6995 15513 7004 15547
rect 6952 15504 7004 15513
rect 7964 15547 8016 15556
rect 7964 15513 7973 15547
rect 7973 15513 8007 15547
rect 8007 15513 8016 15547
rect 7964 15504 8016 15513
rect 10724 15547 10776 15556
rect 10724 15513 10733 15547
rect 10733 15513 10767 15547
rect 10767 15513 10776 15547
rect 10724 15504 10776 15513
rect 11000 15547 11052 15556
rect 11000 15513 11009 15547
rect 11009 15513 11043 15547
rect 11043 15513 11052 15547
rect 11000 15504 11052 15513
rect 4008 15436 4060 15488
rect 4100 15479 4152 15488
rect 4100 15445 4109 15479
rect 4109 15445 4143 15479
rect 4143 15445 4152 15479
rect 4100 15436 4152 15445
rect 4836 15436 4888 15488
rect 5848 15479 5900 15488
rect 5848 15445 5857 15479
rect 5857 15445 5891 15479
rect 5891 15445 5900 15479
rect 5848 15436 5900 15445
rect 2260 15343 2312 15352
rect 2260 15309 2269 15343
rect 2269 15309 2303 15343
rect 2303 15309 2312 15343
rect 2260 15300 2312 15309
rect 4284 15368 4336 15420
rect 7780 15368 7832 15420
rect 8240 15411 8292 15420
rect 8240 15377 8249 15411
rect 8249 15377 8283 15411
rect 8283 15377 8292 15411
rect 8240 15368 8292 15377
rect 8332 15343 8384 15352
rect 3272 15232 3324 15284
rect 8332 15309 8341 15343
rect 8341 15309 8375 15343
rect 8375 15309 8384 15343
rect 8332 15300 8384 15309
rect 9528 15436 9580 15488
rect 12104 15504 12156 15556
rect 14956 15504 15008 15556
rect 15968 15547 16020 15556
rect 15968 15513 15977 15547
rect 15977 15513 16011 15547
rect 16011 15513 16020 15547
rect 15968 15504 16020 15513
rect 22132 15547 22184 15556
rect 22132 15513 22141 15547
rect 22141 15513 22175 15547
rect 22175 15513 22184 15547
rect 22132 15504 22184 15513
rect 22316 15504 22368 15556
rect 22408 15547 22460 15556
rect 22408 15513 22417 15547
rect 22417 15513 22451 15547
rect 22451 15513 22460 15547
rect 22408 15504 22460 15513
rect 24248 15504 24300 15556
rect 26732 15504 26784 15556
rect 11736 15436 11788 15488
rect 11920 15436 11972 15488
rect 23604 15436 23656 15488
rect 17808 15368 17860 15420
rect 18544 15368 18596 15420
rect 19004 15368 19056 15420
rect 20568 15411 20620 15420
rect 20568 15377 20577 15411
rect 20577 15377 20611 15411
rect 20611 15377 20620 15411
rect 20568 15368 20620 15377
rect 26088 15436 26140 15488
rect 27192 15504 27244 15556
rect 28112 15504 28164 15556
rect 28848 15547 28900 15556
rect 28848 15513 28857 15547
rect 28857 15513 28891 15547
rect 28891 15513 28900 15547
rect 28848 15504 28900 15513
rect 26916 15436 26968 15488
rect 28204 15436 28256 15488
rect 11920 15343 11972 15352
rect 6400 15232 6452 15284
rect 7688 15232 7740 15284
rect 11920 15309 11929 15343
rect 11929 15309 11963 15343
rect 11963 15309 11972 15343
rect 11920 15300 11972 15309
rect 18912 15300 18964 15352
rect 24156 15300 24208 15352
rect 24892 15343 24944 15352
rect 24892 15309 24901 15343
rect 24901 15309 24935 15343
rect 24935 15309 24944 15343
rect 24892 15300 24944 15309
rect 25260 15343 25312 15352
rect 25260 15309 25269 15343
rect 25269 15309 25303 15343
rect 25303 15309 25312 15343
rect 25260 15300 25312 15309
rect 25536 15368 25588 15420
rect 26548 15368 26600 15420
rect 27560 15411 27612 15420
rect 27560 15377 27569 15411
rect 27569 15377 27603 15411
rect 27603 15377 27612 15411
rect 27560 15368 27612 15377
rect 27836 15368 27888 15420
rect 27100 15343 27152 15352
rect 27100 15309 27109 15343
rect 27109 15309 27143 15343
rect 27143 15309 27152 15343
rect 27100 15300 27152 15309
rect 27192 15343 27244 15352
rect 27192 15309 27201 15343
rect 27201 15309 27235 15343
rect 27235 15309 27244 15343
rect 27192 15300 27244 15309
rect 13116 15232 13168 15284
rect 5296 15207 5348 15216
rect 5296 15173 5305 15207
rect 5305 15173 5339 15207
rect 5339 15173 5348 15207
rect 5296 15164 5348 15173
rect 14864 15232 14916 15284
rect 18452 15275 18504 15284
rect 18452 15241 18461 15275
rect 18461 15241 18495 15275
rect 18495 15241 18504 15275
rect 18452 15232 18504 15241
rect 22592 15232 22644 15284
rect 14956 15164 15008 15216
rect 15232 15164 15284 15216
rect 15692 15207 15744 15216
rect 15692 15173 15701 15207
rect 15701 15173 15735 15207
rect 15735 15173 15744 15207
rect 15692 15164 15744 15173
rect 18268 15164 18320 15216
rect 20292 15164 20344 15216
rect 22224 15207 22276 15216
rect 22224 15173 22233 15207
rect 22233 15173 22267 15207
rect 22267 15173 22276 15207
rect 22224 15164 22276 15173
rect 24708 15164 24760 15216
rect 26180 15164 26232 15216
rect 28480 15300 28532 15352
rect 28664 15343 28716 15352
rect 28664 15309 28673 15343
rect 28673 15309 28707 15343
rect 28707 15309 28716 15343
rect 28664 15300 28716 15309
rect 27652 15232 27704 15284
rect 28388 15232 28440 15284
rect 18870 15062 18922 15114
rect 18934 15062 18986 15114
rect 18998 15062 19050 15114
rect 19062 15062 19114 15114
rect 19126 15062 19178 15114
rect 1984 14960 2036 15012
rect 3364 15003 3416 15012
rect 3364 14969 3373 15003
rect 3373 14969 3407 15003
rect 3407 14969 3416 15003
rect 3364 14960 3416 14969
rect 5388 14960 5440 15012
rect 6492 14960 6544 15012
rect 7780 15003 7832 15012
rect 7780 14969 7789 15003
rect 7789 14969 7823 15003
rect 7823 14969 7832 15003
rect 7780 14960 7832 14969
rect 7964 15003 8016 15012
rect 7964 14969 7973 15003
rect 7973 14969 8007 15003
rect 8007 14969 8016 15003
rect 7964 14960 8016 14969
rect 8332 14960 8384 15012
rect 12564 14960 12616 15012
rect 18636 14960 18688 15012
rect 20108 14960 20160 15012
rect 27100 14960 27152 15012
rect 28848 14960 28900 15012
rect 10724 14892 10776 14944
rect 11184 14892 11236 14944
rect 14680 14935 14732 14944
rect 14680 14901 14689 14935
rect 14689 14901 14723 14935
rect 14723 14901 14732 14935
rect 14680 14892 14732 14901
rect 14956 14892 15008 14944
rect 18360 14892 18412 14944
rect 18544 14892 18596 14944
rect 25996 14892 26048 14944
rect 27744 14935 27796 14944
rect 4468 14867 4520 14876
rect 4468 14833 4477 14867
rect 4477 14833 4511 14867
rect 4511 14833 4520 14867
rect 4468 14824 4520 14833
rect 4560 14824 4612 14876
rect 4744 14867 4796 14876
rect 4744 14833 4753 14867
rect 4753 14833 4787 14867
rect 4787 14833 4796 14867
rect 4744 14824 4796 14833
rect 4836 14867 4888 14876
rect 4836 14833 4845 14867
rect 4845 14833 4879 14867
rect 4879 14833 4888 14867
rect 4836 14824 4888 14833
rect 6400 14824 6452 14876
rect 11736 14824 11788 14876
rect 23420 14867 23472 14876
rect 23420 14833 23429 14867
rect 23429 14833 23463 14867
rect 23463 14833 23472 14867
rect 23420 14824 23472 14833
rect 26272 14824 26324 14876
rect 26456 14824 26508 14876
rect 27008 14867 27060 14876
rect 27008 14833 27017 14867
rect 27017 14833 27051 14867
rect 27051 14833 27060 14867
rect 27008 14824 27060 14833
rect 27192 14824 27244 14876
rect 27744 14901 27753 14935
rect 27753 14901 27787 14935
rect 27787 14901 27796 14935
rect 27744 14892 27796 14901
rect 4008 14799 4060 14808
rect 4008 14765 4017 14799
rect 4017 14765 4051 14799
rect 4051 14765 4060 14799
rect 4008 14756 4060 14765
rect 4100 14756 4152 14808
rect 5388 14799 5440 14808
rect 1432 14620 1484 14672
rect 5388 14765 5397 14799
rect 5397 14765 5431 14799
rect 5431 14765 5440 14799
rect 5388 14756 5440 14765
rect 11092 14756 11144 14808
rect 14496 14756 14548 14808
rect 24248 14756 24300 14808
rect 26180 14756 26232 14808
rect 10724 14688 10776 14740
rect 6676 14620 6728 14672
rect 26272 14688 26324 14740
rect 14956 14663 15008 14672
rect 14956 14629 14965 14663
rect 14965 14629 14999 14663
rect 14999 14629 15008 14663
rect 14956 14620 15008 14629
rect 19188 14663 19240 14672
rect 19188 14629 19197 14663
rect 19197 14629 19231 14663
rect 19231 14629 19240 14663
rect 19188 14620 19240 14629
rect 24156 14620 24208 14672
rect 3510 14518 3562 14570
rect 3574 14518 3626 14570
rect 3638 14518 3690 14570
rect 3702 14518 3754 14570
rect 3766 14518 3818 14570
rect 4008 14459 4060 14468
rect 4008 14425 4017 14459
rect 4017 14425 4051 14459
rect 4051 14425 4060 14459
rect 4008 14416 4060 14425
rect 4744 14416 4796 14468
rect 6492 14459 6544 14468
rect 6492 14425 6501 14459
rect 6501 14425 6535 14459
rect 6535 14425 6544 14459
rect 6492 14416 6544 14425
rect 6676 14459 6728 14468
rect 6676 14425 6685 14459
rect 6685 14425 6719 14459
rect 6719 14425 6728 14459
rect 6676 14416 6728 14425
rect 11092 14459 11144 14468
rect 11092 14425 11101 14459
rect 11101 14425 11135 14459
rect 11135 14425 11144 14459
rect 11092 14416 11144 14425
rect 11184 14459 11236 14468
rect 11184 14425 11193 14459
rect 11193 14425 11227 14459
rect 11227 14425 11236 14459
rect 11184 14416 11236 14425
rect 11736 14416 11788 14468
rect 12104 14416 12156 14468
rect 14956 14416 15008 14468
rect 15600 14416 15652 14468
rect 16704 14459 16756 14468
rect 16704 14425 16713 14459
rect 16713 14425 16747 14459
rect 16747 14425 16756 14459
rect 16704 14416 16756 14425
rect 17532 14416 17584 14468
rect 18728 14459 18780 14468
rect 18728 14425 18737 14459
rect 18737 14425 18771 14459
rect 18771 14425 18780 14459
rect 18728 14416 18780 14425
rect 26088 14459 26140 14468
rect 26088 14425 26097 14459
rect 26097 14425 26131 14459
rect 26131 14425 26140 14459
rect 26088 14416 26140 14425
rect 26916 14459 26968 14468
rect 26916 14425 26925 14459
rect 26925 14425 26959 14459
rect 26959 14425 26968 14459
rect 26916 14416 26968 14425
rect 5388 14348 5440 14400
rect 1984 14280 2036 14332
rect 4100 14280 4152 14332
rect 4836 14280 4888 14332
rect 5848 14280 5900 14332
rect 696 14255 748 14264
rect 696 14221 705 14255
rect 705 14221 739 14255
rect 739 14221 748 14255
rect 696 14212 748 14221
rect 4560 14255 4612 14264
rect 4560 14221 4569 14255
rect 4569 14221 4603 14255
rect 4603 14221 4612 14255
rect 4560 14212 4612 14221
rect 5480 14212 5532 14264
rect 11184 14212 11236 14264
rect 12104 14212 12156 14264
rect 972 14187 1024 14196
rect 972 14153 981 14187
rect 981 14153 1015 14187
rect 1015 14153 1024 14187
rect 972 14144 1024 14153
rect 1708 14144 1760 14196
rect 8240 14187 8292 14196
rect 8240 14153 8249 14187
rect 8249 14153 8283 14187
rect 8283 14153 8292 14187
rect 8240 14144 8292 14153
rect 15416 14348 15468 14400
rect 16060 14348 16112 14400
rect 3916 14076 3968 14128
rect 4284 14076 4336 14128
rect 5296 14076 5348 14128
rect 6400 14076 6452 14128
rect 11828 14076 11880 14128
rect 14220 14119 14272 14128
rect 14220 14085 14229 14119
rect 14229 14085 14263 14119
rect 14263 14085 14272 14119
rect 14220 14076 14272 14085
rect 15048 14119 15100 14128
rect 15048 14085 15057 14119
rect 15057 14085 15091 14119
rect 15091 14085 15100 14119
rect 15048 14076 15100 14085
rect 16060 14255 16112 14264
rect 16060 14221 16069 14255
rect 16069 14221 16103 14255
rect 16103 14221 16112 14255
rect 18544 14323 18596 14332
rect 18544 14289 18553 14323
rect 18553 14289 18587 14323
rect 18587 14289 18596 14323
rect 18544 14280 18596 14289
rect 16060 14212 16112 14221
rect 15600 14144 15652 14196
rect 15876 14187 15928 14196
rect 15876 14153 15885 14187
rect 15885 14153 15919 14187
rect 15919 14153 15928 14187
rect 15876 14144 15928 14153
rect 15968 14076 16020 14128
rect 17900 14076 17952 14128
rect 18452 14076 18504 14128
rect 19188 14280 19240 14332
rect 20016 14280 20068 14332
rect 19464 14212 19516 14264
rect 20108 14255 20160 14264
rect 20108 14221 20117 14255
rect 20117 14221 20151 14255
rect 20151 14221 20160 14255
rect 20108 14212 20160 14221
rect 26824 14348 26876 14400
rect 28664 14416 28716 14468
rect 25260 14280 25312 14332
rect 20568 14212 20620 14264
rect 22408 14144 22460 14196
rect 26824 14212 26876 14264
rect 24708 14144 24760 14196
rect 27008 14144 27060 14196
rect 23420 14076 23472 14128
rect 24248 14119 24300 14128
rect 24248 14085 24257 14119
rect 24257 14085 24291 14119
rect 24291 14085 24300 14119
rect 24248 14076 24300 14085
rect 25996 14076 26048 14128
rect 26272 14076 26324 14128
rect 28848 14076 28900 14128
rect 29400 14076 29452 14128
rect 18870 13974 18922 14026
rect 18934 13974 18986 14026
rect 18998 13974 19050 14026
rect 19062 13974 19114 14026
rect 19126 13974 19178 14026
rect 972 13872 1024 13924
rect 2628 13872 2680 13924
rect 14680 13915 14732 13924
rect 4100 13804 4152 13856
rect 11828 13847 11880 13856
rect 11828 13813 11837 13847
rect 11837 13813 11871 13847
rect 11871 13813 11880 13847
rect 11828 13804 11880 13813
rect 14680 13881 14689 13915
rect 14689 13881 14723 13915
rect 14723 13881 14732 13915
rect 14680 13872 14732 13881
rect 18268 13872 18320 13924
rect 20108 13872 20160 13924
rect 21028 13872 21080 13924
rect 21672 13915 21724 13924
rect 21672 13881 21681 13915
rect 21681 13881 21715 13915
rect 21715 13881 21724 13915
rect 21672 13872 21724 13881
rect 22224 13872 22276 13924
rect 24800 13915 24852 13924
rect 24800 13881 24809 13915
rect 24809 13881 24843 13915
rect 24843 13881 24852 13915
rect 24800 13872 24852 13881
rect 26364 13872 26416 13924
rect 26916 13872 26968 13924
rect 15140 13804 15192 13856
rect 15324 13804 15376 13856
rect 16060 13804 16112 13856
rect 19372 13804 19424 13856
rect 29124 13804 29176 13856
rect 12840 13779 12892 13788
rect 12840 13745 12849 13779
rect 12849 13745 12883 13779
rect 12883 13745 12892 13779
rect 12840 13736 12892 13745
rect 13116 13736 13168 13788
rect 15048 13736 15100 13788
rect 18636 13779 18688 13788
rect 18636 13745 18645 13779
rect 18645 13745 18679 13779
rect 18679 13745 18688 13779
rect 18636 13736 18688 13745
rect 18728 13779 18780 13788
rect 18728 13745 18737 13779
rect 18737 13745 18771 13779
rect 18771 13745 18780 13779
rect 18728 13736 18780 13745
rect 20016 13736 20068 13788
rect 22132 13736 22184 13788
rect 22408 13779 22460 13788
rect 22408 13745 22417 13779
rect 22417 13745 22451 13779
rect 22451 13745 22460 13779
rect 22408 13736 22460 13745
rect 23420 13779 23472 13788
rect 23420 13745 23429 13779
rect 23429 13745 23463 13779
rect 23463 13745 23472 13779
rect 23420 13736 23472 13745
rect 25812 13779 25864 13788
rect 25812 13745 25821 13779
rect 25821 13745 25855 13779
rect 25855 13745 25864 13779
rect 25812 13736 25864 13745
rect 25904 13779 25956 13788
rect 25904 13745 25913 13779
rect 25913 13745 25947 13779
rect 25947 13745 25956 13779
rect 25904 13736 25956 13745
rect 3364 13711 3416 13720
rect 3364 13677 3373 13711
rect 3373 13677 3407 13711
rect 3407 13677 3416 13711
rect 3364 13668 3416 13677
rect 4008 13668 4060 13720
rect 5388 13711 5440 13720
rect 5388 13677 5397 13711
rect 5397 13677 5431 13711
rect 5431 13677 5440 13711
rect 5388 13668 5440 13677
rect 14404 13668 14456 13720
rect 14864 13668 14916 13720
rect 16336 13668 16388 13720
rect 17348 13711 17400 13720
rect 17348 13677 17357 13711
rect 17357 13677 17391 13711
rect 17391 13677 17400 13711
rect 17348 13668 17400 13677
rect 21856 13711 21908 13720
rect 21856 13677 21865 13711
rect 21865 13677 21899 13711
rect 21899 13677 21908 13711
rect 21856 13668 21908 13677
rect 22316 13711 22368 13720
rect 22316 13677 22325 13711
rect 22325 13677 22359 13711
rect 22359 13677 22368 13711
rect 22316 13668 22368 13677
rect 24156 13668 24208 13720
rect 28388 13711 28440 13720
rect 28388 13677 28397 13711
rect 28397 13677 28431 13711
rect 28431 13677 28440 13711
rect 28388 13668 28440 13677
rect 28756 13711 28808 13720
rect 28756 13677 28765 13711
rect 28765 13677 28799 13711
rect 28799 13677 28808 13711
rect 28756 13668 28808 13677
rect 29032 13668 29084 13720
rect 12380 13600 12432 13652
rect 696 13532 748 13584
rect 972 13575 1024 13584
rect 972 13541 981 13575
rect 981 13541 1015 13575
rect 1015 13541 1024 13575
rect 972 13532 1024 13541
rect 12748 13532 12800 13584
rect 24708 13600 24760 13652
rect 13392 13532 13444 13584
rect 18452 13575 18504 13584
rect 18452 13541 18461 13575
rect 18461 13541 18495 13575
rect 18495 13541 18504 13575
rect 18452 13532 18504 13541
rect 19556 13532 19608 13584
rect 19740 13532 19792 13584
rect 25536 13532 25588 13584
rect 26180 13532 26232 13584
rect 3510 13430 3562 13482
rect 3574 13430 3626 13482
rect 3638 13430 3690 13482
rect 3702 13430 3754 13482
rect 3766 13430 3818 13482
rect 4008 13328 4060 13380
rect 13116 13371 13168 13380
rect 13116 13337 13125 13371
rect 13125 13337 13159 13371
rect 13159 13337 13168 13371
rect 13116 13328 13168 13337
rect 13392 13371 13444 13380
rect 13392 13337 13401 13371
rect 13401 13337 13435 13371
rect 13435 13337 13444 13371
rect 13392 13328 13444 13337
rect 15324 13328 15376 13380
rect 16336 13328 16388 13380
rect 18452 13371 18504 13380
rect 18452 13337 18461 13371
rect 18461 13337 18495 13371
rect 18495 13337 18504 13371
rect 18452 13328 18504 13337
rect 18636 13371 18688 13380
rect 18636 13337 18645 13371
rect 18645 13337 18679 13371
rect 18679 13337 18688 13371
rect 18636 13328 18688 13337
rect 19372 13328 19424 13380
rect 20108 13371 20160 13380
rect 20108 13337 20117 13371
rect 20117 13337 20151 13371
rect 20151 13337 20160 13371
rect 20108 13328 20160 13337
rect 21672 13371 21724 13380
rect 21672 13337 21681 13371
rect 21681 13337 21715 13371
rect 21715 13337 21724 13371
rect 21672 13328 21724 13337
rect 22132 13371 22184 13380
rect 22132 13337 22141 13371
rect 22141 13337 22175 13371
rect 22175 13337 22184 13371
rect 22132 13328 22184 13337
rect 23420 13328 23472 13380
rect 24248 13371 24300 13380
rect 24248 13337 24257 13371
rect 24257 13337 24291 13371
rect 24291 13337 24300 13371
rect 24248 13328 24300 13337
rect 24800 13371 24852 13380
rect 24800 13337 24809 13371
rect 24809 13337 24843 13371
rect 24843 13337 24852 13371
rect 24800 13328 24852 13337
rect 25812 13371 25864 13380
rect 25812 13337 25821 13371
rect 25821 13337 25855 13371
rect 25855 13337 25864 13371
rect 25812 13328 25864 13337
rect 26180 13371 26232 13380
rect 26180 13337 26189 13371
rect 26189 13337 26223 13371
rect 26223 13337 26232 13371
rect 26180 13328 26232 13337
rect 28756 13328 28808 13380
rect 29308 13328 29360 13380
rect 3364 13260 3416 13312
rect 3916 13303 3968 13312
rect 3916 13269 3925 13303
rect 3925 13269 3959 13303
rect 3959 13269 3968 13303
rect 3916 13260 3968 13269
rect 12288 13260 12340 13312
rect 5388 13192 5440 13244
rect 12840 13260 12892 13312
rect 3916 13124 3968 13176
rect 8792 13124 8844 13176
rect 12380 13167 12432 13176
rect 12380 13133 12389 13167
rect 12389 13133 12423 13167
rect 12423 13133 12432 13167
rect 12380 13124 12432 13133
rect 12748 13167 12800 13176
rect 12748 13133 12757 13167
rect 12757 13133 12791 13167
rect 12791 13133 12800 13167
rect 12748 13124 12800 13133
rect 12840 13167 12892 13176
rect 12840 13133 12849 13167
rect 12849 13133 12883 13167
rect 12883 13133 12892 13167
rect 12840 13124 12892 13133
rect 4100 13056 4152 13108
rect 10816 13056 10868 13108
rect 16060 13260 16112 13312
rect 16428 13260 16480 13312
rect 18728 13260 18780 13312
rect 14220 13167 14272 13176
rect 14220 13133 14229 13167
rect 14229 13133 14263 13167
rect 14263 13133 14272 13167
rect 14220 13124 14272 13133
rect 14312 13056 14364 13108
rect 14680 13056 14732 13108
rect 15784 13167 15836 13176
rect 15784 13133 15793 13167
rect 15793 13133 15827 13167
rect 15827 13133 15836 13167
rect 15784 13124 15836 13133
rect 16152 13167 16204 13176
rect 16152 13133 16161 13167
rect 16161 13133 16195 13167
rect 16195 13133 16204 13167
rect 16152 13124 16204 13133
rect 16612 13192 16664 13244
rect 17256 13192 17308 13244
rect 19372 13192 19424 13244
rect 17532 13167 17584 13176
rect 17532 13133 17541 13167
rect 17541 13133 17575 13167
rect 17575 13133 17584 13167
rect 17532 13124 17584 13133
rect 19740 13167 19792 13176
rect 19740 13133 19749 13167
rect 19749 13133 19783 13167
rect 19783 13133 19792 13167
rect 19740 13124 19792 13133
rect 22316 13260 22368 13312
rect 20752 13124 20804 13176
rect 21856 13124 21908 13176
rect 26548 13260 26600 13312
rect 24156 13124 24208 13176
rect 25536 13167 25588 13176
rect 15048 13056 15100 13108
rect 9252 12988 9304 13040
rect 9896 12988 9948 13040
rect 11460 13031 11512 13040
rect 11460 12997 11469 13031
rect 11469 12997 11503 13031
rect 11503 12997 11512 13031
rect 11460 12988 11512 12997
rect 14036 13031 14088 13040
rect 14036 12997 14045 13031
rect 14045 12997 14079 13031
rect 14079 12997 14088 13031
rect 14036 12988 14088 12997
rect 14864 12988 14916 13040
rect 17624 13031 17676 13040
rect 17624 12997 17633 13031
rect 17633 12997 17667 13031
rect 17667 12997 17676 13031
rect 17624 12988 17676 12997
rect 19464 13031 19516 13040
rect 19464 12997 19473 13031
rect 19473 12997 19507 13031
rect 19507 12997 19516 13031
rect 19464 12988 19516 12997
rect 19740 12988 19792 13040
rect 21672 12988 21724 13040
rect 22408 13056 22460 13108
rect 25536 13133 25545 13167
rect 25545 13133 25579 13167
rect 25579 13133 25588 13167
rect 25536 13124 25588 13133
rect 25812 13124 25864 13176
rect 27376 13124 27428 13176
rect 23972 13031 24024 13040
rect 23972 12997 23981 13031
rect 23981 12997 24015 13031
rect 24015 12997 24024 13031
rect 23972 12988 24024 12997
rect 25904 13056 25956 13108
rect 28388 13056 28440 13108
rect 26732 12988 26784 13040
rect 28572 13031 28624 13040
rect 28572 12997 28581 13031
rect 28581 12997 28615 13031
rect 28615 12997 28624 13031
rect 28572 12988 28624 12997
rect 29032 12988 29084 13040
rect 18870 12886 18922 12938
rect 18934 12886 18986 12938
rect 18998 12886 19050 12938
rect 19062 12886 19114 12938
rect 19126 12886 19178 12938
rect 1156 12691 1208 12700
rect 1156 12657 1165 12691
rect 1165 12657 1199 12691
rect 1199 12657 1208 12691
rect 1156 12648 1208 12657
rect 14956 12784 15008 12836
rect 16152 12784 16204 12836
rect 27008 12784 27060 12836
rect 28664 12784 28716 12836
rect 8056 12759 8108 12768
rect 4652 12691 4704 12700
rect 4652 12657 4661 12691
rect 4661 12657 4695 12691
rect 4695 12657 4704 12691
rect 4652 12648 4704 12657
rect 8056 12725 8065 12759
rect 8065 12725 8099 12759
rect 8099 12725 8108 12759
rect 8056 12716 8108 12725
rect 11460 12716 11512 12768
rect 7412 12648 7464 12700
rect 7964 12648 8016 12700
rect 11276 12648 11328 12700
rect 12288 12716 12340 12768
rect 12380 12716 12432 12768
rect 12472 12648 12524 12700
rect 12840 12648 12892 12700
rect 14220 12648 14272 12700
rect 15784 12716 15836 12768
rect 14772 12691 14824 12700
rect 14772 12657 14781 12691
rect 14781 12657 14815 12691
rect 14815 12657 14824 12691
rect 14772 12648 14824 12657
rect 14956 12648 15008 12700
rect 15232 12648 15284 12700
rect 16336 12648 16388 12700
rect 17348 12716 17400 12768
rect 18544 12716 18596 12768
rect 18820 12648 18872 12700
rect 29124 12716 29176 12768
rect 21948 12648 22000 12700
rect 23420 12648 23472 12700
rect 24340 12691 24392 12700
rect 24340 12657 24349 12691
rect 24349 12657 24383 12691
rect 24383 12657 24392 12691
rect 24340 12648 24392 12657
rect 24708 12691 24760 12700
rect 24708 12657 24717 12691
rect 24717 12657 24751 12691
rect 24751 12657 24760 12691
rect 24708 12648 24760 12657
rect 1708 12580 1760 12632
rect 3272 12580 3324 12632
rect 4836 12623 4888 12632
rect 4836 12589 4845 12623
rect 4845 12589 4879 12623
rect 4879 12589 4888 12623
rect 4836 12580 4888 12589
rect 5848 12580 5900 12632
rect 6124 12580 6176 12632
rect 6308 12623 6360 12632
rect 6308 12589 6317 12623
rect 6317 12589 6351 12623
rect 6351 12589 6360 12623
rect 6308 12580 6360 12589
rect 9896 12623 9948 12632
rect 9896 12589 9905 12623
rect 9905 12589 9939 12623
rect 9939 12589 9948 12623
rect 9896 12580 9948 12589
rect 10816 12580 10868 12632
rect 13300 12623 13352 12632
rect 13300 12589 13309 12623
rect 13309 12589 13343 12623
rect 13343 12589 13352 12623
rect 13300 12580 13352 12589
rect 16612 12580 16664 12632
rect 16980 12623 17032 12632
rect 16980 12589 16989 12623
rect 16989 12589 17023 12623
rect 17023 12589 17032 12623
rect 16980 12580 17032 12589
rect 17348 12623 17400 12632
rect 17348 12589 17357 12623
rect 17357 12589 17391 12623
rect 17391 12589 17400 12623
rect 17348 12580 17400 12589
rect 18176 12580 18228 12632
rect 19556 12580 19608 12632
rect 24156 12623 24208 12632
rect 24156 12589 24165 12623
rect 24165 12589 24199 12623
rect 24199 12589 24208 12623
rect 24156 12580 24208 12589
rect 23144 12512 23196 12564
rect 25260 12648 25312 12700
rect 27376 12648 27428 12700
rect 26364 12580 26416 12632
rect 28388 12623 28440 12632
rect 28388 12589 28397 12623
rect 28397 12589 28431 12623
rect 28431 12589 28440 12623
rect 28388 12580 28440 12589
rect 28756 12623 28808 12632
rect 28756 12589 28765 12623
rect 28765 12589 28799 12623
rect 28799 12589 28808 12623
rect 28756 12580 28808 12589
rect 30136 12623 30188 12632
rect 30136 12589 30145 12623
rect 30145 12589 30179 12623
rect 30179 12589 30188 12623
rect 30136 12580 30188 12589
rect 8516 12444 8568 12496
rect 16428 12444 16480 12496
rect 18452 12444 18504 12496
rect 19464 12444 19516 12496
rect 20568 12444 20620 12496
rect 21764 12487 21816 12496
rect 21764 12453 21773 12487
rect 21773 12453 21807 12487
rect 21807 12453 21816 12487
rect 21764 12444 21816 12453
rect 23880 12444 23932 12496
rect 3510 12342 3562 12394
rect 3574 12342 3626 12394
rect 3638 12342 3690 12394
rect 3702 12342 3754 12394
rect 3766 12342 3818 12394
rect 1708 12283 1760 12292
rect 1708 12249 1717 12283
rect 1717 12249 1751 12283
rect 1751 12249 1760 12283
rect 1708 12240 1760 12249
rect 1248 12147 1300 12156
rect 1248 12113 1257 12147
rect 1257 12113 1291 12147
rect 1291 12113 1300 12147
rect 4100 12240 4152 12292
rect 4652 12283 4704 12292
rect 4652 12249 4661 12283
rect 4661 12249 4695 12283
rect 4695 12249 4704 12283
rect 4652 12240 4704 12249
rect 6308 12240 6360 12292
rect 10540 12240 10592 12292
rect 10816 12283 10868 12292
rect 10816 12249 10825 12283
rect 10825 12249 10859 12283
rect 10859 12249 10868 12283
rect 10816 12240 10868 12249
rect 12380 12240 12432 12292
rect 13300 12283 13352 12292
rect 13300 12249 13309 12283
rect 13309 12249 13343 12283
rect 13343 12249 13352 12283
rect 14772 12283 14824 12292
rect 13300 12240 13352 12249
rect 14772 12249 14781 12283
rect 14781 12249 14815 12283
rect 14815 12249 14824 12283
rect 14772 12240 14824 12249
rect 15232 12283 15284 12292
rect 15232 12249 15241 12283
rect 15241 12249 15275 12283
rect 15275 12249 15284 12283
rect 15232 12240 15284 12249
rect 16152 12283 16204 12292
rect 16152 12249 16161 12283
rect 16161 12249 16195 12283
rect 16195 12249 16204 12283
rect 16152 12240 16204 12249
rect 16612 12283 16664 12292
rect 16612 12249 16621 12283
rect 16621 12249 16655 12283
rect 16655 12249 16664 12283
rect 16612 12240 16664 12249
rect 16980 12240 17032 12292
rect 18452 12283 18504 12292
rect 18452 12249 18461 12283
rect 18461 12249 18495 12283
rect 18495 12249 18504 12283
rect 18452 12240 18504 12249
rect 18728 12240 18780 12292
rect 21948 12283 22000 12292
rect 21948 12249 21957 12283
rect 21957 12249 21991 12283
rect 21991 12249 22000 12283
rect 21948 12240 22000 12249
rect 24708 12240 24760 12292
rect 27008 12240 27060 12292
rect 28756 12240 28808 12292
rect 11460 12172 11512 12224
rect 14220 12172 14272 12224
rect 18544 12215 18596 12224
rect 18544 12181 18553 12215
rect 18553 12181 18587 12215
rect 18587 12181 18596 12215
rect 18544 12172 18596 12181
rect 21028 12172 21080 12224
rect 23144 12215 23196 12224
rect 23144 12181 23153 12215
rect 23153 12181 23187 12215
rect 23187 12181 23196 12215
rect 23144 12172 23196 12181
rect 28388 12172 28440 12224
rect 1248 12104 1300 12113
rect 5112 12104 5164 12156
rect 8148 12147 8200 12156
rect 1156 11900 1208 11952
rect 2444 11900 2496 11952
rect 3272 12036 3324 12088
rect 6124 12036 6176 12088
rect 6584 12079 6636 12088
rect 6584 12045 6593 12079
rect 6593 12045 6627 12079
rect 6627 12045 6636 12079
rect 6584 12036 6636 12045
rect 6768 12079 6820 12088
rect 6768 12045 6777 12079
rect 6777 12045 6811 12079
rect 6811 12045 6820 12079
rect 6768 12036 6820 12045
rect 8148 12113 8157 12147
rect 8157 12113 8191 12147
rect 8191 12113 8200 12147
rect 8148 12104 8200 12113
rect 8516 12147 8568 12156
rect 8516 12113 8525 12147
rect 8525 12113 8559 12147
rect 8559 12113 8568 12147
rect 8516 12104 8568 12113
rect 9804 12104 9856 12156
rect 8056 12036 8108 12088
rect 11276 12104 11328 12156
rect 14036 12104 14088 12156
rect 12380 12079 12432 12088
rect 7872 11968 7924 12020
rect 4836 11943 4888 11952
rect 4836 11909 4845 11943
rect 4845 11909 4879 11943
rect 4879 11909 4888 11943
rect 4836 11900 4888 11909
rect 5940 11943 5992 11952
rect 5940 11909 5949 11943
rect 5949 11909 5983 11943
rect 5983 11909 5992 11943
rect 5940 11900 5992 11909
rect 7688 11900 7740 11952
rect 7964 11900 8016 11952
rect 8792 11900 8844 11952
rect 12380 12045 12389 12079
rect 12389 12045 12423 12079
rect 12423 12045 12432 12079
rect 12380 12036 12432 12045
rect 17348 12104 17400 12156
rect 17624 12104 17676 12156
rect 14036 11968 14088 12020
rect 17440 12036 17492 12088
rect 18820 12036 18872 12088
rect 23236 12104 23288 12156
rect 24248 12104 24300 12156
rect 25260 12147 25312 12156
rect 25260 12113 25269 12147
rect 25269 12113 25303 12147
rect 25303 12113 25312 12147
rect 25260 12104 25312 12113
rect 26824 12104 26876 12156
rect 28940 12104 28992 12156
rect 17808 11968 17860 12020
rect 20752 12036 20804 12088
rect 21304 12079 21356 12088
rect 21304 12045 21313 12079
rect 21313 12045 21347 12079
rect 21347 12045 21356 12079
rect 21304 12036 21356 12045
rect 21672 12079 21724 12088
rect 21672 12045 21681 12079
rect 21681 12045 21715 12079
rect 21715 12045 21724 12079
rect 21672 12036 21724 12045
rect 21856 12079 21908 12088
rect 21856 12045 21865 12079
rect 21865 12045 21899 12079
rect 21899 12045 21908 12079
rect 21856 12036 21908 12045
rect 23052 12036 23104 12088
rect 23512 12079 23564 12088
rect 23512 12045 23521 12079
rect 23521 12045 23555 12079
rect 23555 12045 23564 12079
rect 23512 12036 23564 12045
rect 23880 12079 23932 12088
rect 23880 12045 23889 12079
rect 23889 12045 23923 12079
rect 23923 12045 23932 12079
rect 23880 12036 23932 12045
rect 27284 12079 27336 12088
rect 20660 12011 20712 12020
rect 20660 11977 20669 12011
rect 20669 11977 20703 12011
rect 20703 11977 20712 12011
rect 20660 11968 20712 11977
rect 12564 11900 12616 11952
rect 14956 11943 15008 11952
rect 14956 11909 14965 11943
rect 14965 11909 14999 11943
rect 14999 11909 15008 11943
rect 14956 11900 15008 11909
rect 19464 11900 19516 11952
rect 20108 11943 20160 11952
rect 20108 11909 20117 11943
rect 20117 11909 20151 11943
rect 20151 11909 20160 11943
rect 20108 11900 20160 11909
rect 20568 11900 20620 11952
rect 21764 11968 21816 12020
rect 23236 11900 23288 11952
rect 24248 11968 24300 12020
rect 26732 12011 26784 12020
rect 26732 11977 26741 12011
rect 26741 11977 26775 12011
rect 26775 11977 26784 12011
rect 27284 12045 27293 12079
rect 27293 12045 27327 12079
rect 27327 12045 27336 12079
rect 27284 12036 27336 12045
rect 29216 12079 29268 12088
rect 26732 11968 26784 11977
rect 27192 11968 27244 12020
rect 28572 11968 28624 12020
rect 29216 12045 29225 12079
rect 29225 12045 29259 12079
rect 29259 12045 29268 12079
rect 29216 12036 29268 12045
rect 29584 12079 29636 12088
rect 29584 12045 29593 12079
rect 29593 12045 29627 12079
rect 29627 12045 29636 12079
rect 29584 12036 29636 12045
rect 30136 12036 30188 12088
rect 29124 11968 29176 12020
rect 27376 11943 27428 11952
rect 27376 11909 27385 11943
rect 27385 11909 27419 11943
rect 27419 11909 27428 11943
rect 27376 11900 27428 11909
rect 18870 11798 18922 11850
rect 18934 11798 18986 11850
rect 18998 11798 19050 11850
rect 19062 11798 19114 11850
rect 19126 11798 19178 11850
rect 6308 11739 6360 11748
rect 6308 11705 6317 11739
rect 6317 11705 6351 11739
rect 6351 11705 6360 11739
rect 6308 11696 6360 11705
rect 8148 11739 8200 11748
rect 8148 11705 8157 11739
rect 8157 11705 8191 11739
rect 8191 11705 8200 11739
rect 8148 11696 8200 11705
rect 9896 11696 9948 11748
rect 16336 11739 16388 11748
rect 8516 11628 8568 11680
rect 9160 11628 9212 11680
rect 16336 11705 16345 11739
rect 16345 11705 16379 11739
rect 16379 11705 16388 11739
rect 16336 11696 16388 11705
rect 16428 11739 16480 11748
rect 16428 11705 16437 11739
rect 16437 11705 16471 11739
rect 16471 11705 16480 11739
rect 16428 11696 16480 11705
rect 16980 11696 17032 11748
rect 17532 11696 17584 11748
rect 18728 11696 18780 11748
rect 20108 11696 20160 11748
rect 21304 11696 21356 11748
rect 23052 11739 23104 11748
rect 23052 11705 23061 11739
rect 23061 11705 23095 11739
rect 23095 11705 23104 11739
rect 23052 11696 23104 11705
rect 23144 11696 23196 11748
rect 23880 11739 23932 11748
rect 23880 11705 23889 11739
rect 23889 11705 23923 11739
rect 23923 11705 23932 11739
rect 24156 11739 24208 11748
rect 23880 11696 23932 11705
rect 24156 11705 24165 11739
rect 24165 11705 24199 11739
rect 24199 11705 24208 11739
rect 24156 11696 24208 11705
rect 14404 11628 14456 11680
rect 19280 11628 19332 11680
rect 21672 11628 21724 11680
rect 24064 11628 24116 11680
rect 27192 11628 27244 11680
rect 28756 11696 28808 11748
rect 29124 11628 29176 11680
rect 29308 11671 29360 11680
rect 29308 11637 29317 11671
rect 29317 11637 29351 11671
rect 29351 11637 29360 11671
rect 29308 11628 29360 11637
rect 1340 11560 1392 11612
rect 9068 11560 9120 11612
rect 9988 11603 10040 11612
rect 9988 11569 9997 11603
rect 9997 11569 10031 11603
rect 10031 11569 10040 11603
rect 9988 11560 10040 11569
rect 12564 11603 12616 11612
rect 12564 11569 12573 11603
rect 12573 11569 12607 11603
rect 12607 11569 12616 11603
rect 12564 11560 12616 11569
rect 17624 11603 17676 11612
rect 17624 11569 17633 11603
rect 17633 11569 17667 11603
rect 17667 11569 17676 11603
rect 17624 11560 17676 11569
rect 20660 11560 20712 11612
rect 21304 11603 21356 11612
rect 21304 11569 21313 11603
rect 21313 11569 21347 11603
rect 21347 11569 21356 11603
rect 21304 11560 21356 11569
rect 6768 11535 6820 11544
rect 6768 11501 6777 11535
rect 6777 11501 6811 11535
rect 6811 11501 6820 11535
rect 6768 11492 6820 11501
rect 9528 11492 9580 11544
rect 9712 11535 9764 11544
rect 9712 11501 9721 11535
rect 9721 11501 9755 11535
rect 9755 11501 9764 11535
rect 9712 11492 9764 11501
rect 6584 11467 6636 11476
rect 6584 11433 6593 11467
rect 6593 11433 6627 11467
rect 6627 11433 6636 11467
rect 6584 11424 6636 11433
rect 7596 11424 7648 11476
rect 8884 11424 8936 11476
rect 9804 11424 9856 11476
rect 12380 11492 12432 11544
rect 14036 11492 14088 11544
rect 18360 11492 18412 11544
rect 21488 11492 21540 11544
rect 22500 11492 22552 11544
rect 23512 11535 23564 11544
rect 23512 11501 23521 11535
rect 23521 11501 23555 11535
rect 23555 11501 23564 11535
rect 23512 11492 23564 11501
rect 26364 11535 26416 11544
rect 26364 11501 26373 11535
rect 26373 11501 26407 11535
rect 26407 11501 26416 11535
rect 26364 11492 26416 11501
rect 26732 11535 26784 11544
rect 26732 11501 26741 11535
rect 26741 11501 26775 11535
rect 26775 11501 26784 11535
rect 26732 11492 26784 11501
rect 28112 11535 28164 11544
rect 28112 11501 28121 11535
rect 28121 11501 28155 11535
rect 28155 11501 28164 11535
rect 28112 11492 28164 11501
rect 28204 11492 28256 11544
rect 29216 11492 29268 11544
rect 29860 11560 29912 11612
rect 29676 11492 29728 11544
rect 30228 11535 30280 11544
rect 30228 11501 30237 11535
rect 30237 11501 30271 11535
rect 30271 11501 30280 11535
rect 30228 11492 30280 11501
rect 12656 11424 12708 11476
rect 20660 11467 20712 11476
rect 20660 11433 20669 11467
rect 20669 11433 20703 11467
rect 20703 11433 20712 11467
rect 20660 11424 20712 11433
rect 27468 11424 27520 11476
rect 29584 11424 29636 11476
rect 30044 11424 30096 11476
rect 1432 11399 1484 11408
rect 1432 11365 1441 11399
rect 1441 11365 1475 11399
rect 1475 11365 1484 11399
rect 1432 11356 1484 11365
rect 6400 11356 6452 11408
rect 12748 11399 12800 11408
rect 12748 11365 12757 11399
rect 12757 11365 12791 11399
rect 12791 11365 12800 11399
rect 12748 11356 12800 11365
rect 24340 11399 24392 11408
rect 24340 11365 24349 11399
rect 24349 11365 24383 11399
rect 24383 11365 24392 11399
rect 24340 11356 24392 11365
rect 28664 11356 28716 11408
rect 3510 11254 3562 11306
rect 3574 11254 3626 11306
rect 3638 11254 3690 11306
rect 3702 11254 3754 11306
rect 3766 11254 3818 11306
rect 1340 11195 1392 11204
rect 1340 11161 1349 11195
rect 1349 11161 1383 11195
rect 1383 11161 1392 11195
rect 1340 11152 1392 11161
rect 7688 11152 7740 11204
rect 8884 11152 8936 11204
rect 9160 11195 9212 11204
rect 9160 11161 9169 11195
rect 9169 11161 9203 11195
rect 9203 11161 9212 11195
rect 9160 11152 9212 11161
rect 12564 11152 12616 11204
rect 13116 11152 13168 11204
rect 14956 11152 15008 11204
rect 15416 11195 15468 11204
rect 15416 11161 15425 11195
rect 15425 11161 15459 11195
rect 15459 11161 15468 11195
rect 15416 11152 15468 11161
rect 15692 11152 15744 11204
rect 17532 11195 17584 11204
rect 17532 11161 17541 11195
rect 17541 11161 17575 11195
rect 17575 11161 17584 11195
rect 17532 11152 17584 11161
rect 17624 11152 17676 11204
rect 21304 11195 21356 11204
rect 21304 11161 21313 11195
rect 21313 11161 21347 11195
rect 21347 11161 21356 11195
rect 21304 11152 21356 11161
rect 21488 11195 21540 11204
rect 21488 11161 21497 11195
rect 21497 11161 21531 11195
rect 21531 11161 21540 11195
rect 21488 11152 21540 11161
rect 26732 11195 26784 11204
rect 26732 11161 26741 11195
rect 26741 11161 26775 11195
rect 26775 11161 26784 11195
rect 26732 11152 26784 11161
rect 29308 11152 29360 11204
rect 29860 11195 29912 11204
rect 29860 11161 29869 11195
rect 29869 11161 29903 11195
rect 29903 11161 29912 11195
rect 29860 11152 29912 11161
rect 30044 11195 30096 11204
rect 30044 11161 30053 11195
rect 30053 11161 30087 11195
rect 30087 11161 30096 11195
rect 30044 11152 30096 11161
rect 7596 11084 7648 11136
rect 9712 11084 9764 11136
rect 12380 11127 12432 11136
rect 12380 11093 12389 11127
rect 12389 11093 12423 11127
rect 12423 11093 12432 11127
rect 12380 11084 12432 11093
rect 12656 11084 12708 11136
rect 17440 11084 17492 11136
rect 6400 11016 6452 11068
rect 7872 11016 7924 11068
rect 9988 11016 10040 11068
rect 12564 11016 12616 11068
rect 2444 10991 2496 11000
rect 2444 10957 2453 10991
rect 2453 10957 2487 10991
rect 2487 10957 2496 10991
rect 2444 10948 2496 10957
rect 6124 10991 6176 11000
rect 6124 10957 6133 10991
rect 6133 10957 6167 10991
rect 6167 10957 6176 10991
rect 6124 10948 6176 10957
rect 1432 10855 1484 10864
rect 1432 10821 1441 10855
rect 1441 10821 1475 10855
rect 1475 10821 1484 10855
rect 1432 10812 1484 10821
rect 7412 10880 7464 10932
rect 2996 10855 3048 10864
rect 2996 10821 3005 10855
rect 3005 10821 3039 10855
rect 3039 10821 3048 10855
rect 2996 10812 3048 10821
rect 5664 10855 5716 10864
rect 5664 10821 5673 10855
rect 5673 10821 5707 10855
rect 5707 10821 5716 10855
rect 5664 10812 5716 10821
rect 5940 10855 5992 10864
rect 5940 10821 5949 10855
rect 5949 10821 5983 10855
rect 5983 10821 5992 10855
rect 5940 10812 5992 10821
rect 7780 10812 7832 10864
rect 13300 10991 13352 11000
rect 13300 10957 13309 10991
rect 13309 10957 13343 10991
rect 13343 10957 13352 10991
rect 13300 10948 13352 10957
rect 13760 10991 13812 11000
rect 13760 10957 13769 10991
rect 13769 10957 13803 10991
rect 13803 10957 13812 10991
rect 15692 11016 15744 11068
rect 17716 11127 17768 11136
rect 17716 11093 17725 11127
rect 17725 11093 17759 11127
rect 17759 11093 17768 11127
rect 17716 11084 17768 11093
rect 17808 11084 17860 11136
rect 13760 10948 13812 10957
rect 14772 10948 14824 11000
rect 15416 10948 15468 11000
rect 17808 10991 17860 11000
rect 17808 10957 17817 10991
rect 17817 10957 17851 10991
rect 17851 10957 17860 10991
rect 17808 10948 17860 10957
rect 21856 11084 21908 11136
rect 25352 11084 25404 11136
rect 27008 11016 27060 11068
rect 28112 11016 28164 11068
rect 29124 11016 29176 11068
rect 29308 11016 29360 11068
rect 24892 10948 24944 11000
rect 26640 10948 26692 11000
rect 27100 10991 27152 11000
rect 27100 10957 27109 10991
rect 27109 10957 27143 10991
rect 27143 10957 27152 10991
rect 27100 10948 27152 10957
rect 27468 10991 27520 11000
rect 27468 10957 27477 10991
rect 27477 10957 27511 10991
rect 27511 10957 27520 10991
rect 27468 10948 27520 10957
rect 28756 10948 28808 11000
rect 29676 10991 29728 11000
rect 29676 10957 29685 10991
rect 29685 10957 29719 10991
rect 29719 10957 29728 10991
rect 29676 10948 29728 10957
rect 10172 10855 10224 10864
rect 10172 10821 10181 10855
rect 10181 10821 10215 10855
rect 10215 10821 10224 10855
rect 10172 10812 10224 10821
rect 10264 10812 10316 10864
rect 13576 10812 13628 10864
rect 16060 10880 16112 10932
rect 18728 10880 18780 10932
rect 21948 10880 22000 10932
rect 27192 10880 27244 10932
rect 19924 10812 19976 10864
rect 20292 10812 20344 10864
rect 21672 10812 21724 10864
rect 23236 10812 23288 10864
rect 26916 10812 26968 10864
rect 27468 10812 27520 10864
rect 29124 10812 29176 10864
rect 30228 10880 30280 10932
rect 18870 10710 18922 10762
rect 18934 10710 18986 10762
rect 18998 10710 19050 10762
rect 19062 10710 19114 10762
rect 19126 10710 19178 10762
rect 12564 10608 12616 10660
rect 13116 10651 13168 10660
rect 13116 10617 13125 10651
rect 13125 10617 13159 10651
rect 13159 10617 13168 10651
rect 13116 10608 13168 10617
rect 14864 10608 14916 10660
rect 18452 10608 18504 10660
rect 19280 10608 19332 10660
rect 26732 10608 26784 10660
rect 27100 10608 27152 10660
rect 28020 10608 28072 10660
rect 28664 10608 28716 10660
rect 6400 10540 6452 10592
rect 7044 10540 7096 10592
rect 13760 10540 13812 10592
rect 16244 10583 16296 10592
rect 16244 10549 16253 10583
rect 16253 10549 16287 10583
rect 16287 10549 16296 10583
rect 16244 10540 16296 10549
rect 17624 10540 17676 10592
rect 26640 10583 26692 10592
rect 26640 10549 26649 10583
rect 26649 10549 26683 10583
rect 26683 10549 26692 10583
rect 26640 10540 26692 10549
rect 28204 10540 28256 10592
rect 2996 10472 3048 10524
rect 4468 10472 4520 10524
rect 7872 10515 7924 10524
rect 7872 10481 7881 10515
rect 7881 10481 7915 10515
rect 7915 10481 7924 10515
rect 7872 10472 7924 10481
rect 12748 10472 12800 10524
rect 13576 10515 13628 10524
rect 13576 10481 13585 10515
rect 13585 10481 13619 10515
rect 13619 10481 13628 10515
rect 13576 10472 13628 10481
rect 14680 10472 14732 10524
rect 14772 10515 14824 10524
rect 14772 10481 14781 10515
rect 14781 10481 14815 10515
rect 14815 10481 14824 10515
rect 14772 10472 14824 10481
rect 16336 10515 16388 10524
rect 16336 10481 16345 10515
rect 16345 10481 16379 10515
rect 16379 10481 16388 10515
rect 16336 10472 16388 10481
rect 17716 10472 17768 10524
rect 18636 10472 18688 10524
rect 18820 10472 18872 10524
rect 26088 10515 26140 10524
rect 26088 10481 26097 10515
rect 26097 10481 26131 10515
rect 26131 10481 26140 10515
rect 26088 10472 26140 10481
rect 29768 10472 29820 10524
rect 1984 10404 2036 10456
rect 4100 10404 4152 10456
rect 7412 10404 7464 10456
rect 7596 10447 7648 10456
rect 7596 10413 7605 10447
rect 7605 10413 7639 10447
rect 7639 10413 7648 10447
rect 7596 10404 7648 10413
rect 7780 10447 7832 10456
rect 7780 10413 7789 10447
rect 7789 10413 7823 10447
rect 7823 10413 7832 10447
rect 7780 10404 7832 10413
rect 18452 10404 18504 10456
rect 13300 10336 13352 10388
rect 18912 10404 18964 10456
rect 19464 10404 19516 10456
rect 22960 10447 23012 10456
rect 22960 10413 22969 10447
rect 22969 10413 23003 10447
rect 23003 10413 23012 10447
rect 22960 10404 23012 10413
rect 23788 10404 23840 10456
rect 24340 10404 24392 10456
rect 3916 10268 3968 10320
rect 4560 10268 4612 10320
rect 6124 10268 6176 10320
rect 8148 10268 8200 10320
rect 8976 10311 9028 10320
rect 8976 10277 8985 10311
rect 8985 10277 9019 10311
rect 9019 10277 9028 10311
rect 8976 10268 9028 10277
rect 14128 10268 14180 10320
rect 14864 10311 14916 10320
rect 14864 10277 14873 10311
rect 14873 10277 14907 10311
rect 14907 10277 14916 10311
rect 14864 10268 14916 10277
rect 16060 10311 16112 10320
rect 16060 10277 16069 10311
rect 16069 10277 16103 10311
rect 16103 10277 16112 10311
rect 16060 10268 16112 10277
rect 20108 10336 20160 10388
rect 24248 10336 24300 10388
rect 26364 10404 26416 10456
rect 25628 10336 25680 10388
rect 16612 10268 16664 10320
rect 17440 10311 17492 10320
rect 17440 10277 17449 10311
rect 17449 10277 17483 10311
rect 17483 10277 17492 10311
rect 17440 10268 17492 10277
rect 18360 10311 18412 10320
rect 18360 10277 18369 10311
rect 18369 10277 18403 10311
rect 18403 10277 18412 10311
rect 18360 10268 18412 10277
rect 23144 10311 23196 10320
rect 23144 10277 23153 10311
rect 23153 10277 23187 10311
rect 23187 10277 23196 10311
rect 23144 10268 23196 10277
rect 25904 10311 25956 10320
rect 25904 10277 25913 10311
rect 25913 10277 25947 10311
rect 25947 10277 25956 10311
rect 25904 10268 25956 10277
rect 29676 10268 29728 10320
rect 3510 10166 3562 10218
rect 3574 10166 3626 10218
rect 3638 10166 3690 10218
rect 3702 10166 3754 10218
rect 3766 10166 3818 10218
rect 1984 10107 2036 10116
rect 1984 10073 1993 10107
rect 1993 10073 2027 10107
rect 2027 10073 2036 10107
rect 1984 10064 2036 10073
rect 4468 10107 4520 10116
rect 4468 10073 4477 10107
rect 4477 10073 4511 10107
rect 4511 10073 4520 10107
rect 4468 10064 4520 10073
rect 4560 10107 4612 10116
rect 4560 10073 4569 10107
rect 4569 10073 4603 10107
rect 4603 10073 4612 10107
rect 7044 10107 7096 10116
rect 4560 10064 4612 10073
rect 7044 10073 7053 10107
rect 7053 10073 7087 10107
rect 7087 10073 7096 10107
rect 7044 10064 7096 10073
rect 7596 10064 7648 10116
rect 8792 10064 8844 10116
rect 9528 10064 9580 10116
rect 13760 10064 13812 10116
rect 14128 10107 14180 10116
rect 14128 10073 14137 10107
rect 14137 10073 14171 10107
rect 14171 10073 14180 10107
rect 14128 10064 14180 10073
rect 14496 10107 14548 10116
rect 14496 10073 14505 10107
rect 14505 10073 14539 10107
rect 14539 10073 14548 10107
rect 14496 10064 14548 10073
rect 14772 10064 14824 10116
rect 16060 10107 16112 10116
rect 7872 9996 7924 10048
rect 2076 9971 2128 9980
rect 2076 9937 2085 9971
rect 2085 9937 2119 9971
rect 2119 9937 2128 9971
rect 2076 9928 2128 9937
rect 4100 9971 4152 9980
rect 4100 9937 4109 9971
rect 4109 9937 4143 9971
rect 4143 9937 4152 9971
rect 4100 9928 4152 9937
rect 7412 9928 7464 9980
rect 7596 9971 7648 9980
rect 7596 9937 7605 9971
rect 7605 9937 7639 9971
rect 7639 9937 7648 9971
rect 7596 9928 7648 9937
rect 8148 9928 8200 9980
rect 8792 9971 8844 9980
rect 8792 9937 8801 9971
rect 8801 9937 8835 9971
rect 8835 9937 8844 9971
rect 8792 9928 8844 9937
rect 13576 9928 13628 9980
rect 16060 10073 16069 10107
rect 16069 10073 16103 10107
rect 16103 10073 16112 10107
rect 16060 10064 16112 10073
rect 16244 10107 16296 10116
rect 16244 10073 16253 10107
rect 16253 10073 16287 10107
rect 16287 10073 16296 10107
rect 16244 10064 16296 10073
rect 16612 10107 16664 10116
rect 16612 10073 16621 10107
rect 16621 10073 16655 10107
rect 16655 10073 16664 10107
rect 16612 10064 16664 10073
rect 17440 10064 17492 10116
rect 18360 10107 18412 10116
rect 18360 10073 18369 10107
rect 18369 10073 18403 10107
rect 18403 10073 18412 10107
rect 18360 10064 18412 10073
rect 19924 10064 19976 10116
rect 24616 10064 24668 10116
rect 26088 10064 26140 10116
rect 28664 10107 28716 10116
rect 28664 10073 28673 10107
rect 28673 10073 28707 10107
rect 28707 10073 28716 10107
rect 28664 10064 28716 10073
rect 16336 9996 16388 10048
rect 17532 9996 17584 10048
rect 25352 9996 25404 10048
rect 26180 9996 26232 10048
rect 7504 9860 7556 9912
rect 8424 9903 8476 9912
rect 8424 9869 8433 9903
rect 8433 9869 8467 9903
rect 8467 9869 8476 9903
rect 8424 9860 8476 9869
rect 2352 9835 2404 9844
rect 2352 9801 2361 9835
rect 2361 9801 2395 9835
rect 2395 9801 2404 9835
rect 2352 9792 2404 9801
rect 2996 9792 3048 9844
rect 5664 9724 5716 9776
rect 7780 9792 7832 9844
rect 9344 9792 9396 9844
rect 9528 9792 9580 9844
rect 10816 9835 10868 9844
rect 10816 9801 10825 9835
rect 10825 9801 10859 9835
rect 10859 9801 10868 9835
rect 10816 9792 10868 9801
rect 14496 9792 14548 9844
rect 15876 9860 15928 9912
rect 15968 9860 16020 9912
rect 19280 9928 19332 9980
rect 20384 9928 20436 9980
rect 19096 9860 19148 9912
rect 19464 9860 19516 9912
rect 23052 9860 23104 9912
rect 23420 9903 23472 9912
rect 23420 9869 23429 9903
rect 23429 9869 23463 9903
rect 23463 9869 23472 9903
rect 23420 9860 23472 9869
rect 28296 9928 28348 9980
rect 29584 9996 29636 10048
rect 11552 9724 11604 9776
rect 15048 9792 15100 9844
rect 18912 9792 18964 9844
rect 14772 9724 14824 9776
rect 18360 9724 18412 9776
rect 19924 9792 19976 9844
rect 22868 9792 22920 9844
rect 23144 9792 23196 9844
rect 21488 9724 21540 9776
rect 23696 9724 23748 9776
rect 24616 9860 24668 9912
rect 25720 9903 25772 9912
rect 25720 9869 25729 9903
rect 25729 9869 25763 9903
rect 25763 9869 25772 9903
rect 25720 9860 25772 9869
rect 26180 9903 26232 9912
rect 26180 9869 26189 9903
rect 26189 9869 26223 9903
rect 26223 9869 26232 9903
rect 26180 9860 26232 9869
rect 29216 9903 29268 9912
rect 29216 9869 29225 9903
rect 29225 9869 29259 9903
rect 29259 9869 29268 9903
rect 29216 9860 29268 9869
rect 25352 9767 25404 9776
rect 25352 9733 25361 9767
rect 25361 9733 25395 9767
rect 25395 9733 25404 9767
rect 25352 9724 25404 9733
rect 27100 9724 27152 9776
rect 27284 9724 27336 9776
rect 29584 9903 29636 9912
rect 29584 9869 29593 9903
rect 29593 9869 29627 9903
rect 29627 9869 29636 9903
rect 29768 9903 29820 9912
rect 29584 9860 29636 9869
rect 29768 9869 29777 9903
rect 29777 9869 29811 9903
rect 29811 9869 29820 9903
rect 29768 9860 29820 9869
rect 18870 9622 18922 9674
rect 18934 9622 18986 9674
rect 18998 9622 19050 9674
rect 19062 9622 19114 9674
rect 19126 9622 19178 9674
rect 2076 9563 2128 9572
rect 2076 9529 2085 9563
rect 2085 9529 2119 9563
rect 2119 9529 2128 9563
rect 2076 9520 2128 9529
rect 8792 9520 8844 9572
rect 12288 9520 12340 9572
rect 14680 9563 14732 9572
rect 14680 9529 14689 9563
rect 14689 9529 14723 9563
rect 14723 9529 14732 9563
rect 14680 9520 14732 9529
rect 18636 9563 18688 9572
rect 18636 9529 18645 9563
rect 18645 9529 18679 9563
rect 18679 9529 18688 9563
rect 18636 9520 18688 9529
rect 18728 9520 18780 9572
rect 19280 9520 19332 9572
rect 24616 9563 24668 9572
rect 24616 9529 24625 9563
rect 24625 9529 24659 9563
rect 24659 9529 24668 9563
rect 24616 9520 24668 9529
rect 24708 9520 24760 9572
rect 25536 9520 25588 9572
rect 25904 9563 25956 9572
rect 25904 9529 25913 9563
rect 25913 9529 25947 9563
rect 25947 9529 25956 9563
rect 25904 9520 25956 9529
rect 2352 9452 2404 9504
rect 3180 9452 3232 9504
rect 4100 9452 4152 9504
rect 5480 9495 5532 9504
rect 5480 9461 5489 9495
rect 5489 9461 5523 9495
rect 5523 9461 5532 9495
rect 5480 9452 5532 9461
rect 9344 9495 9396 9504
rect 9344 9461 9353 9495
rect 9353 9461 9387 9495
rect 9387 9461 9396 9495
rect 9344 9452 9396 9461
rect 14772 9452 14824 9504
rect 17348 9452 17400 9504
rect 1156 9427 1208 9436
rect 1156 9393 1165 9427
rect 1165 9393 1199 9427
rect 1199 9393 1208 9427
rect 1156 9384 1208 9393
rect 2444 9384 2496 9436
rect 3916 9384 3968 9436
rect 4008 9427 4060 9436
rect 4008 9393 4017 9427
rect 4017 9393 4051 9427
rect 4051 9393 4060 9427
rect 4192 9427 4244 9436
rect 4008 9384 4060 9393
rect 4192 9393 4201 9427
rect 4201 9393 4235 9427
rect 4235 9393 4244 9427
rect 4192 9384 4244 9393
rect 5572 9384 5624 9436
rect 9988 9427 10040 9436
rect 9988 9393 9997 9427
rect 9997 9393 10031 9427
rect 10031 9393 10040 9427
rect 9988 9384 10040 9393
rect 10356 9427 10408 9436
rect 10356 9393 10365 9427
rect 10365 9393 10399 9427
rect 10399 9393 10408 9427
rect 10356 9384 10408 9393
rect 15968 9384 16020 9436
rect 17992 9427 18044 9436
rect 17992 9393 18001 9427
rect 18001 9393 18035 9427
rect 18035 9393 18044 9427
rect 17992 9384 18044 9393
rect 23236 9452 23288 9504
rect 26364 9452 26416 9504
rect 27560 9452 27612 9504
rect 27652 9452 27704 9504
rect 28388 9495 28440 9504
rect 28388 9461 28397 9495
rect 28397 9461 28431 9495
rect 28431 9461 28440 9495
rect 28388 9452 28440 9461
rect 28572 9452 28624 9504
rect 19372 9384 19424 9436
rect 22500 9427 22552 9436
rect 22500 9393 22509 9427
rect 22509 9393 22543 9427
rect 22543 9393 22552 9427
rect 22500 9384 22552 9393
rect 22868 9427 22920 9436
rect 22868 9393 22877 9427
rect 22877 9393 22911 9427
rect 22911 9393 22920 9427
rect 22868 9384 22920 9393
rect 26640 9427 26692 9436
rect 26640 9393 26649 9427
rect 26649 9393 26683 9427
rect 26683 9393 26692 9427
rect 26640 9384 26692 9393
rect 27008 9427 27060 9436
rect 1432 9359 1484 9368
rect 1432 9325 1441 9359
rect 1441 9325 1475 9359
rect 1475 9325 1484 9359
rect 1432 9316 1484 9325
rect 6032 9359 6084 9368
rect 6032 9325 6041 9359
rect 6041 9325 6075 9359
rect 6075 9325 6084 9359
rect 6032 9316 6084 9325
rect 9436 9316 9488 9368
rect 9620 9316 9672 9368
rect 9712 9248 9764 9300
rect 10816 9316 10868 9368
rect 18084 9359 18136 9368
rect 18084 9325 18093 9359
rect 18093 9325 18127 9359
rect 18127 9325 18136 9359
rect 18084 9316 18136 9325
rect 18452 9359 18504 9368
rect 18452 9325 18461 9359
rect 18461 9325 18495 9359
rect 18495 9325 18504 9359
rect 18452 9316 18504 9325
rect 22776 9316 22828 9368
rect 24616 9316 24668 9368
rect 25996 9316 26048 9368
rect 27008 9393 27017 9427
rect 27017 9393 27051 9427
rect 27051 9393 27060 9427
rect 27008 9384 27060 9393
rect 27468 9427 27520 9436
rect 27192 9359 27244 9368
rect 27192 9325 27201 9359
rect 27201 9325 27235 9359
rect 27235 9325 27244 9359
rect 27192 9316 27244 9325
rect 25720 9248 25772 9300
rect 27468 9393 27477 9427
rect 27477 9393 27511 9427
rect 27511 9393 27520 9427
rect 27468 9384 27520 9393
rect 28848 9427 28900 9436
rect 28848 9393 28857 9427
rect 28857 9393 28891 9427
rect 28891 9393 28900 9427
rect 28848 9384 28900 9393
rect 29124 9384 29176 9436
rect 28664 9316 28716 9368
rect 28480 9248 28532 9300
rect 30044 9248 30096 9300
rect 1616 9180 1668 9232
rect 6492 9180 6544 9232
rect 12012 9223 12064 9232
rect 12012 9189 12021 9223
rect 12021 9189 12055 9223
rect 12055 9189 12064 9223
rect 12012 9180 12064 9189
rect 16152 9223 16204 9232
rect 16152 9189 16161 9223
rect 16161 9189 16195 9223
rect 16195 9189 16204 9223
rect 16152 9180 16204 9189
rect 17532 9180 17584 9232
rect 3510 9078 3562 9130
rect 3574 9078 3626 9130
rect 3638 9078 3690 9130
rect 3702 9078 3754 9130
rect 3766 9078 3818 9130
rect 2076 8976 2128 9028
rect 3180 9019 3232 9028
rect 3180 8985 3189 9019
rect 3189 8985 3223 9019
rect 3223 8985 3232 9019
rect 3180 8976 3232 8985
rect 4468 9019 4520 9028
rect 4468 8985 4477 9019
rect 4477 8985 4511 9019
rect 4511 8985 4520 9019
rect 4468 8976 4520 8985
rect 5480 9019 5532 9028
rect 5480 8985 5489 9019
rect 5489 8985 5523 9019
rect 5523 8985 5532 9019
rect 5480 8976 5532 8985
rect 9344 8976 9396 9028
rect 14588 8976 14640 9028
rect 15692 8976 15744 9028
rect 15968 9019 16020 9028
rect 15968 8985 15977 9019
rect 15977 8985 16011 9019
rect 16011 8985 16020 9019
rect 15968 8976 16020 8985
rect 16152 8976 16204 9028
rect 18452 8976 18504 9028
rect 19372 8976 19424 9028
rect 22776 9019 22828 9028
rect 22776 8985 22785 9019
rect 22785 8985 22819 9019
rect 22819 8985 22828 9019
rect 22776 8976 22828 8985
rect 22868 8976 22920 9028
rect 24708 9019 24760 9028
rect 24708 8985 24717 9019
rect 24717 8985 24751 9019
rect 24751 8985 24760 9019
rect 24708 8976 24760 8985
rect 25536 8976 25588 9028
rect 27192 8976 27244 9028
rect 27468 8976 27520 9028
rect 28480 8976 28532 9028
rect 29124 8976 29176 9028
rect 29216 8976 29268 9028
rect 6032 8908 6084 8960
rect 7872 8908 7924 8960
rect 8700 8908 8752 8960
rect 10356 8908 10408 8960
rect 12748 8908 12800 8960
rect 18268 8908 18320 8960
rect 696 8883 748 8892
rect 696 8849 705 8883
rect 705 8849 739 8883
rect 739 8849 748 8883
rect 696 8840 748 8849
rect 1616 8840 1668 8892
rect 4192 8883 4244 8892
rect 4192 8849 4201 8883
rect 4201 8849 4235 8883
rect 4235 8849 4244 8883
rect 4192 8840 4244 8849
rect 4744 8840 4796 8892
rect 6492 8883 6544 8892
rect 3640 8815 3692 8824
rect 3640 8781 3649 8815
rect 3649 8781 3683 8815
rect 3683 8781 3692 8815
rect 3640 8772 3692 8781
rect 4468 8772 4520 8824
rect 6124 8815 6176 8824
rect 6124 8781 6133 8815
rect 6133 8781 6167 8815
rect 6167 8781 6176 8815
rect 6124 8772 6176 8781
rect 6492 8849 6501 8883
rect 6501 8849 6535 8883
rect 6535 8849 6544 8883
rect 6492 8840 6544 8849
rect 7412 8840 7464 8892
rect 8424 8840 8476 8892
rect 9712 8840 9764 8892
rect 9988 8840 10040 8892
rect 12012 8840 12064 8892
rect 12656 8883 12708 8892
rect 12288 8772 12340 8824
rect 12656 8849 12665 8883
rect 12665 8849 12699 8883
rect 12699 8849 12708 8883
rect 12656 8840 12708 8849
rect 17992 8840 18044 8892
rect 22500 8908 22552 8960
rect 12748 8815 12800 8824
rect 12748 8781 12757 8815
rect 12757 8781 12791 8815
rect 12791 8781 12800 8815
rect 12748 8772 12800 8781
rect 972 8747 1024 8756
rect 972 8713 981 8747
rect 981 8713 1015 8747
rect 1015 8713 1024 8747
rect 972 8704 1024 8713
rect 1432 8704 1484 8756
rect 2904 8747 2956 8756
rect 2904 8713 2913 8747
rect 2913 8713 2947 8747
rect 2947 8713 2956 8747
rect 2904 8704 2956 8713
rect 7320 8704 7372 8756
rect 11184 8704 11236 8756
rect 12656 8704 12708 8756
rect 14588 8747 14640 8756
rect 14588 8713 14597 8747
rect 14597 8713 14631 8747
rect 14631 8713 14640 8747
rect 14588 8704 14640 8713
rect 14772 8815 14824 8824
rect 14772 8781 14781 8815
rect 14781 8781 14815 8815
rect 14815 8781 14824 8815
rect 14772 8772 14824 8781
rect 17440 8772 17492 8824
rect 18728 8772 18780 8824
rect 23328 8840 23380 8892
rect 24616 8908 24668 8960
rect 25628 8908 25680 8960
rect 27008 8908 27060 8960
rect 29032 8951 29084 8960
rect 29032 8917 29041 8951
rect 29041 8917 29075 8951
rect 29075 8917 29084 8951
rect 29032 8908 29084 8917
rect 25904 8840 25956 8892
rect 26640 8840 26692 8892
rect 17348 8747 17400 8756
rect 17348 8713 17357 8747
rect 17357 8713 17391 8747
rect 17391 8713 17400 8747
rect 17348 8704 17400 8713
rect 17808 8747 17860 8756
rect 17808 8713 17817 8747
rect 17817 8713 17851 8747
rect 17851 8713 17860 8747
rect 17808 8704 17860 8713
rect 18084 8704 18136 8756
rect 21212 8772 21264 8824
rect 25352 8772 25404 8824
rect 25628 8815 25680 8824
rect 21764 8704 21816 8756
rect 25168 8704 25220 8756
rect 25628 8781 25637 8815
rect 25637 8781 25671 8815
rect 25671 8781 25680 8815
rect 25628 8772 25680 8781
rect 27100 8815 27152 8824
rect 27100 8781 27109 8815
rect 27109 8781 27143 8815
rect 27143 8781 27152 8815
rect 27100 8772 27152 8781
rect 27284 8772 27336 8824
rect 27468 8815 27520 8824
rect 27468 8781 27477 8815
rect 27477 8781 27511 8815
rect 27511 8781 27520 8815
rect 27468 8772 27520 8781
rect 27652 8815 27704 8824
rect 27652 8781 27661 8815
rect 27661 8781 27695 8815
rect 27695 8781 27704 8815
rect 27652 8772 27704 8781
rect 28848 8772 28900 8824
rect 29400 8772 29452 8824
rect 26456 8747 26508 8756
rect 26456 8713 26465 8747
rect 26465 8713 26499 8747
rect 26499 8713 26508 8747
rect 26456 8704 26508 8713
rect 29216 8747 29268 8756
rect 29216 8713 29225 8747
rect 29225 8713 29259 8747
rect 29259 8713 29268 8747
rect 29216 8704 29268 8713
rect 4008 8636 4060 8688
rect 5480 8636 5532 8688
rect 7780 8636 7832 8688
rect 9436 8636 9488 8688
rect 11460 8679 11512 8688
rect 11460 8645 11469 8679
rect 11469 8645 11503 8679
rect 11503 8645 11512 8679
rect 11460 8636 11512 8645
rect 14772 8636 14824 8688
rect 24340 8636 24392 8688
rect 25720 8679 25772 8688
rect 25720 8645 25729 8679
rect 25729 8645 25763 8679
rect 25763 8645 25772 8679
rect 25720 8636 25772 8645
rect 25904 8679 25956 8688
rect 25904 8645 25913 8679
rect 25913 8645 25947 8679
rect 25947 8645 25956 8679
rect 25904 8636 25956 8645
rect 28664 8636 28716 8688
rect 18870 8534 18922 8586
rect 18934 8534 18986 8586
rect 18998 8534 19050 8586
rect 19062 8534 19114 8586
rect 19126 8534 19178 8586
rect 696 8432 748 8484
rect 1432 8432 1484 8484
rect 3916 8475 3968 8484
rect 3916 8441 3925 8475
rect 3925 8441 3959 8475
rect 3959 8441 3968 8475
rect 3916 8432 3968 8441
rect 17992 8432 18044 8484
rect 26364 8475 26416 8484
rect 26364 8441 26373 8475
rect 26373 8441 26407 8475
rect 26407 8441 26416 8475
rect 26364 8432 26416 8441
rect 27100 8475 27152 8484
rect 27100 8441 27109 8475
rect 27109 8441 27143 8475
rect 27143 8441 27152 8475
rect 27100 8432 27152 8441
rect 28388 8475 28440 8484
rect 28388 8441 28397 8475
rect 28397 8441 28431 8475
rect 28431 8441 28440 8475
rect 28388 8432 28440 8441
rect 29400 8475 29452 8484
rect 29400 8441 29409 8475
rect 29409 8441 29443 8475
rect 29443 8441 29452 8475
rect 29400 8432 29452 8441
rect 30044 8475 30096 8484
rect 30044 8441 30053 8475
rect 30053 8441 30087 8475
rect 30087 8441 30096 8475
rect 30044 8432 30096 8441
rect 2904 8364 2956 8416
rect 1800 8228 1852 8280
rect 2352 8339 2404 8348
rect 2352 8305 2361 8339
rect 2361 8305 2395 8339
rect 2395 8305 2404 8339
rect 4008 8364 4060 8416
rect 4192 8364 4244 8416
rect 5296 8407 5348 8416
rect 5296 8373 5305 8407
rect 5305 8373 5339 8407
rect 5339 8373 5348 8407
rect 5296 8364 5348 8373
rect 2352 8296 2404 8305
rect 3364 8296 3416 8348
rect 3640 8339 3692 8348
rect 3640 8305 3649 8339
rect 3649 8305 3683 8339
rect 3683 8305 3692 8339
rect 3640 8296 3692 8305
rect 5480 8339 5532 8348
rect 5480 8305 5489 8339
rect 5489 8305 5523 8339
rect 5523 8305 5532 8339
rect 5480 8296 5532 8305
rect 6216 8296 6268 8348
rect 7136 8296 7188 8348
rect 9988 8364 10040 8416
rect 11552 8364 11604 8416
rect 17532 8407 17584 8416
rect 17532 8373 17541 8407
rect 17541 8373 17575 8407
rect 17575 8373 17584 8407
rect 17532 8364 17584 8373
rect 24616 8364 24668 8416
rect 26456 8364 26508 8416
rect 27376 8364 27428 8416
rect 7872 8339 7924 8348
rect 7872 8305 7881 8339
rect 7881 8305 7915 8339
rect 7915 8305 7924 8339
rect 7872 8296 7924 8305
rect 5848 8271 5900 8280
rect 5848 8237 5857 8271
rect 5857 8237 5891 8271
rect 5891 8237 5900 8271
rect 5848 8228 5900 8237
rect 6860 8271 6912 8280
rect 6860 8237 6869 8271
rect 6869 8237 6903 8271
rect 6903 8237 6912 8271
rect 6860 8228 6912 8237
rect 6952 8228 7004 8280
rect 972 8160 1024 8212
rect 1708 8203 1760 8212
rect 1708 8169 1717 8203
rect 1717 8169 1751 8203
rect 1751 8169 1760 8203
rect 1708 8160 1760 8169
rect 6400 8160 6452 8212
rect 8792 8296 8844 8348
rect 10816 8339 10868 8348
rect 10816 8305 10825 8339
rect 10825 8305 10859 8339
rect 10859 8305 10868 8339
rect 10816 8296 10868 8305
rect 11184 8339 11236 8348
rect 11184 8305 11193 8339
rect 11193 8305 11227 8339
rect 11227 8305 11236 8339
rect 11184 8296 11236 8305
rect 20936 8339 20988 8348
rect 20936 8305 20945 8339
rect 20945 8305 20979 8339
rect 20979 8305 20988 8339
rect 20936 8296 20988 8305
rect 21212 8339 21264 8348
rect 21212 8305 21221 8339
rect 21221 8305 21255 8339
rect 21255 8305 21264 8339
rect 21212 8296 21264 8305
rect 21764 8339 21816 8348
rect 21764 8305 21773 8339
rect 21773 8305 21807 8339
rect 21807 8305 21816 8339
rect 21764 8296 21816 8305
rect 22868 8339 22920 8348
rect 22868 8305 22877 8339
rect 22877 8305 22911 8339
rect 22911 8305 22920 8339
rect 22868 8296 22920 8305
rect 24340 8296 24392 8348
rect 24524 8296 24576 8348
rect 25352 8296 25404 8348
rect 27468 8296 27520 8348
rect 11460 8228 11512 8280
rect 12656 8228 12708 8280
rect 8608 8160 8660 8212
rect 20568 8160 20620 8212
rect 22040 8228 22092 8280
rect 23512 8228 23564 8280
rect 25904 8228 25956 8280
rect 29216 8339 29268 8348
rect 29216 8305 29225 8339
rect 29225 8305 29259 8339
rect 29259 8305 29268 8339
rect 29216 8296 29268 8305
rect 28572 8228 28624 8280
rect 21580 8160 21632 8212
rect 6124 8092 6176 8144
rect 7044 8092 7096 8144
rect 14312 8092 14364 8144
rect 26640 8160 26692 8212
rect 27652 8160 27704 8212
rect 23052 8135 23104 8144
rect 23052 8101 23061 8135
rect 23061 8101 23095 8135
rect 23095 8101 23104 8135
rect 23052 8092 23104 8101
rect 25076 8135 25128 8144
rect 25076 8101 25085 8135
rect 25085 8101 25119 8135
rect 25119 8101 25128 8135
rect 25076 8092 25128 8101
rect 27284 8092 27336 8144
rect 3510 7990 3562 8042
rect 3574 7990 3626 8042
rect 3638 7990 3690 8042
rect 3702 7990 3754 8042
rect 3766 7990 3818 8042
rect 1708 7888 1760 7940
rect 2904 7888 2956 7940
rect 3364 7931 3416 7940
rect 3364 7897 3373 7931
rect 3373 7897 3407 7931
rect 3407 7897 3416 7931
rect 3364 7888 3416 7897
rect 4008 7888 4060 7940
rect 5296 7931 5348 7940
rect 5296 7897 5305 7931
rect 5305 7897 5339 7931
rect 5339 7897 5348 7931
rect 5296 7888 5348 7897
rect 5848 7888 5900 7940
rect 6216 7931 6268 7940
rect 6216 7897 6225 7931
rect 6225 7897 6259 7931
rect 6259 7897 6268 7931
rect 6216 7888 6268 7897
rect 6400 7931 6452 7940
rect 6400 7897 6409 7931
rect 6409 7897 6443 7931
rect 6443 7897 6452 7931
rect 6400 7888 6452 7897
rect 6860 7888 6912 7940
rect 11184 7931 11236 7940
rect 11184 7897 11193 7931
rect 11193 7897 11227 7931
rect 11227 7897 11236 7931
rect 11184 7888 11236 7897
rect 14312 7931 14364 7940
rect 14312 7897 14321 7931
rect 14321 7897 14355 7931
rect 14355 7897 14364 7931
rect 14312 7888 14364 7897
rect 17440 7888 17492 7940
rect 17992 7888 18044 7940
rect 21212 7888 21264 7940
rect 21580 7888 21632 7940
rect 23052 7888 23104 7940
rect 23972 7888 24024 7940
rect 25536 7888 25588 7940
rect 27468 7888 27520 7940
rect 29216 7931 29268 7940
rect 2352 7752 2404 7804
rect 10816 7820 10868 7872
rect 20936 7863 20988 7872
rect 20936 7829 20945 7863
rect 20945 7829 20979 7863
rect 20979 7829 20988 7863
rect 20936 7820 20988 7829
rect 22868 7820 22920 7872
rect 23512 7863 23564 7872
rect 23512 7829 23521 7863
rect 23521 7829 23555 7863
rect 23555 7829 23564 7863
rect 23512 7820 23564 7829
rect 23788 7863 23840 7872
rect 23788 7829 23797 7863
rect 23797 7829 23831 7863
rect 23831 7829 23840 7863
rect 23788 7820 23840 7829
rect 23880 7820 23932 7872
rect 24800 7820 24852 7872
rect 7228 7752 7280 7804
rect 8608 7752 8660 7804
rect 10356 7752 10408 7804
rect 11552 7752 11604 7804
rect 1156 7727 1208 7736
rect 1156 7693 1165 7727
rect 1165 7693 1199 7727
rect 1199 7693 1208 7727
rect 1156 7684 1208 7693
rect 7044 7727 7096 7736
rect 7044 7693 7053 7727
rect 7053 7693 7087 7727
rect 7087 7693 7096 7727
rect 7044 7684 7096 7693
rect 7504 7684 7556 7736
rect 12288 7684 12340 7736
rect 14312 7684 14364 7736
rect 14864 7684 14916 7736
rect 15784 7752 15836 7804
rect 23236 7795 23288 7804
rect 15140 7684 15192 7736
rect 1432 7659 1484 7668
rect 1432 7625 1441 7659
rect 1441 7625 1475 7659
rect 1475 7625 1484 7659
rect 1432 7616 1484 7625
rect 7780 7616 7832 7668
rect 8792 7616 8844 7668
rect 11460 7616 11512 7668
rect 1800 7591 1852 7600
rect 1800 7557 1809 7591
rect 1809 7557 1843 7591
rect 1843 7557 1852 7591
rect 1800 7548 1852 7557
rect 5480 7591 5532 7600
rect 5480 7557 5489 7591
rect 5489 7557 5523 7591
rect 5523 7557 5532 7591
rect 5480 7548 5532 7557
rect 6768 7591 6820 7600
rect 6768 7557 6777 7591
rect 6777 7557 6811 7591
rect 6811 7557 6820 7591
rect 6768 7548 6820 7557
rect 14036 7548 14088 7600
rect 14404 7591 14456 7600
rect 14404 7557 14413 7591
rect 14413 7557 14447 7591
rect 14447 7557 14456 7591
rect 14404 7548 14456 7557
rect 14680 7548 14732 7600
rect 16796 7548 16848 7600
rect 23236 7761 23245 7795
rect 23245 7761 23279 7795
rect 23279 7761 23288 7795
rect 23236 7752 23288 7761
rect 21764 7684 21816 7736
rect 24892 7752 24944 7804
rect 25536 7727 25588 7736
rect 23604 7616 23656 7668
rect 23972 7616 24024 7668
rect 24340 7659 24392 7668
rect 24340 7625 24349 7659
rect 24349 7625 24383 7659
rect 24383 7625 24392 7659
rect 24340 7616 24392 7625
rect 24616 7616 24668 7668
rect 25076 7616 25128 7668
rect 25536 7693 25545 7727
rect 25545 7693 25579 7727
rect 25579 7693 25588 7727
rect 25536 7684 25588 7693
rect 29216 7897 29225 7931
rect 29225 7897 29259 7931
rect 29259 7897 29268 7931
rect 29216 7888 29268 7897
rect 30044 7888 30096 7940
rect 28572 7727 28624 7736
rect 28572 7693 28581 7727
rect 28581 7693 28615 7727
rect 28615 7693 28624 7727
rect 28572 7684 28624 7693
rect 20568 7591 20620 7600
rect 20568 7557 20577 7591
rect 20577 7557 20611 7591
rect 20611 7557 20620 7591
rect 20568 7548 20620 7557
rect 28112 7591 28164 7600
rect 28112 7557 28121 7591
rect 28121 7557 28155 7591
rect 28155 7557 28164 7591
rect 28112 7548 28164 7557
rect 18870 7446 18922 7498
rect 18934 7446 18986 7498
rect 18998 7446 19050 7498
rect 19062 7446 19114 7498
rect 19126 7446 19178 7498
rect 6952 7387 7004 7396
rect 6952 7353 6961 7387
rect 6961 7353 6995 7387
rect 6995 7353 7004 7387
rect 6952 7344 7004 7353
rect 7228 7387 7280 7396
rect 7228 7353 7237 7387
rect 7237 7353 7271 7387
rect 7271 7353 7280 7387
rect 7228 7344 7280 7353
rect 7504 7387 7556 7396
rect 7504 7353 7513 7387
rect 7513 7353 7547 7387
rect 7547 7353 7556 7387
rect 7504 7344 7556 7353
rect 8884 7344 8936 7396
rect 23236 7344 23288 7396
rect 24340 7387 24392 7396
rect 24340 7353 24349 7387
rect 24349 7353 24383 7387
rect 24383 7353 24392 7387
rect 24340 7344 24392 7353
rect 24524 7387 24576 7396
rect 24524 7353 24533 7387
rect 24533 7353 24567 7387
rect 24567 7353 24576 7387
rect 24524 7344 24576 7353
rect 24708 7387 24760 7396
rect 24708 7353 24717 7387
rect 24717 7353 24751 7387
rect 24751 7353 24760 7387
rect 24708 7344 24760 7353
rect 24892 7387 24944 7396
rect 24892 7353 24901 7387
rect 24901 7353 24935 7387
rect 24935 7353 24944 7387
rect 24892 7344 24944 7353
rect 5940 7276 5992 7328
rect 6768 7276 6820 7328
rect 8608 7276 8660 7328
rect 18728 7319 18780 7328
rect 18728 7285 18737 7319
rect 18737 7285 18771 7319
rect 18771 7285 18780 7319
rect 18728 7276 18780 7285
rect 23696 7276 23748 7328
rect 26640 7276 26692 7328
rect 3364 7208 3416 7260
rect 5296 7251 5348 7260
rect 5296 7217 5305 7251
rect 5305 7217 5339 7251
rect 5339 7217 5348 7251
rect 5296 7208 5348 7217
rect 5480 7251 5532 7260
rect 5480 7217 5489 7251
rect 5489 7217 5523 7251
rect 5523 7217 5532 7251
rect 5480 7208 5532 7217
rect 12288 7251 12340 7260
rect 12288 7217 12297 7251
rect 12297 7217 12331 7251
rect 12331 7217 12340 7251
rect 12288 7208 12340 7217
rect 14680 7208 14732 7260
rect 14956 7208 15008 7260
rect 17808 7208 17860 7260
rect 18176 7251 18228 7260
rect 18176 7217 18185 7251
rect 18185 7217 18219 7251
rect 18219 7217 18228 7251
rect 18176 7208 18228 7217
rect 18452 7208 18504 7260
rect 23052 7208 23104 7260
rect 28664 7276 28716 7328
rect 28112 7208 28164 7260
rect 3916 7140 3968 7192
rect 26548 7140 26600 7192
rect 27836 7140 27888 7192
rect 28756 7140 28808 7192
rect 28020 7072 28072 7124
rect 29584 7072 29636 7124
rect 8148 7004 8200 7056
rect 11552 7004 11604 7056
rect 12748 7004 12800 7056
rect 15140 7047 15192 7056
rect 15140 7013 15149 7047
rect 15149 7013 15183 7047
rect 15183 7013 15192 7047
rect 15140 7004 15192 7013
rect 20200 7004 20252 7056
rect 20936 7004 20988 7056
rect 26916 7047 26968 7056
rect 26916 7013 26925 7047
rect 26925 7013 26959 7047
rect 26959 7013 26968 7047
rect 26916 7004 26968 7013
rect 28480 7047 28532 7056
rect 28480 7013 28489 7047
rect 28489 7013 28523 7047
rect 28523 7013 28532 7047
rect 28480 7004 28532 7013
rect 3510 6902 3562 6954
rect 3574 6902 3626 6954
rect 3638 6902 3690 6954
rect 3702 6902 3754 6954
rect 3766 6902 3818 6954
rect 3364 6800 3416 6852
rect 4008 6800 4060 6852
rect 4836 6800 4888 6852
rect 5296 6843 5348 6852
rect 5296 6809 5305 6843
rect 5305 6809 5339 6843
rect 5339 6809 5348 6843
rect 5296 6800 5348 6809
rect 5940 6800 5992 6852
rect 6492 6800 6544 6852
rect 7136 6775 7188 6784
rect 7136 6741 7145 6775
rect 7145 6741 7179 6775
rect 7179 6741 7188 6775
rect 7136 6732 7188 6741
rect 7412 6732 7464 6784
rect 2904 6503 2956 6512
rect 2904 6469 2913 6503
rect 2913 6469 2947 6503
rect 2947 6469 2956 6503
rect 2904 6460 2956 6469
rect 3088 6460 3140 6512
rect 3916 6503 3968 6512
rect 3916 6469 3925 6503
rect 3925 6469 3959 6503
rect 3959 6469 3968 6503
rect 3916 6460 3968 6469
rect 4100 6460 4152 6512
rect 8148 6707 8200 6716
rect 8148 6673 8157 6707
rect 8157 6673 8191 6707
rect 8191 6673 8200 6707
rect 8148 6664 8200 6673
rect 8700 6639 8752 6648
rect 8700 6605 8709 6639
rect 8709 6605 8743 6639
rect 8743 6605 8752 6639
rect 8700 6596 8752 6605
rect 8884 6800 8936 6852
rect 11552 6775 11604 6784
rect 11552 6741 11561 6775
rect 11561 6741 11595 6775
rect 11595 6741 11604 6775
rect 11552 6732 11604 6741
rect 4376 6528 4428 6580
rect 5480 6528 5532 6580
rect 6584 6528 6636 6580
rect 6676 6528 6728 6580
rect 12288 6800 12340 6852
rect 12748 6843 12800 6852
rect 12748 6809 12757 6843
rect 12757 6809 12791 6843
rect 12791 6809 12800 6843
rect 12748 6800 12800 6809
rect 15140 6800 15192 6852
rect 15232 6800 15284 6852
rect 18176 6843 18228 6852
rect 18176 6809 18185 6843
rect 18185 6809 18219 6843
rect 18219 6809 18228 6843
rect 18176 6800 18228 6809
rect 18728 6800 18780 6852
rect 23052 6800 23104 6852
rect 17808 6732 17860 6784
rect 12196 6664 12248 6716
rect 13944 6664 13996 6716
rect 11552 6528 11604 6580
rect 13208 6596 13260 6648
rect 10816 6460 10868 6512
rect 18268 6596 18320 6648
rect 20200 6664 20252 6716
rect 23696 6732 23748 6784
rect 24616 6800 24668 6852
rect 24892 6800 24944 6852
rect 28112 6800 28164 6852
rect 28296 6843 28348 6852
rect 28296 6809 28305 6843
rect 28305 6809 28339 6843
rect 28339 6809 28348 6843
rect 28296 6800 28348 6809
rect 25536 6732 25588 6784
rect 26640 6732 26692 6784
rect 26916 6732 26968 6784
rect 27836 6775 27888 6784
rect 27836 6741 27845 6775
rect 27845 6741 27879 6775
rect 27879 6741 27888 6775
rect 27836 6732 27888 6741
rect 28020 6664 28072 6716
rect 29308 6707 29360 6716
rect 29308 6673 29317 6707
rect 29317 6673 29351 6707
rect 29351 6673 29360 6707
rect 29308 6664 29360 6673
rect 20936 6639 20988 6648
rect 14680 6528 14732 6580
rect 14864 6503 14916 6512
rect 14864 6469 14873 6503
rect 14873 6469 14907 6503
rect 14907 6469 14916 6503
rect 14864 6460 14916 6469
rect 15416 6528 15468 6580
rect 16336 6460 16388 6512
rect 18452 6503 18504 6512
rect 18452 6469 18461 6503
rect 18461 6469 18495 6503
rect 18495 6469 18504 6503
rect 18452 6460 18504 6469
rect 20568 6528 20620 6580
rect 20936 6605 20945 6639
rect 20945 6605 20979 6639
rect 20979 6605 20988 6639
rect 20936 6596 20988 6605
rect 21120 6596 21172 6648
rect 21948 6596 22000 6648
rect 23420 6596 23472 6648
rect 23696 6596 23748 6648
rect 24248 6639 24300 6648
rect 24248 6605 24257 6639
rect 24257 6605 24291 6639
rect 24291 6605 24300 6639
rect 24248 6596 24300 6605
rect 24340 6596 24392 6648
rect 25444 6596 25496 6648
rect 26548 6596 26600 6648
rect 29216 6639 29268 6648
rect 29216 6605 29225 6639
rect 29225 6605 29259 6639
rect 29259 6605 29268 6639
rect 29216 6596 29268 6605
rect 29584 6639 29636 6648
rect 29584 6605 29593 6639
rect 29593 6605 29627 6639
rect 29627 6605 29636 6639
rect 29584 6596 29636 6605
rect 21672 6528 21724 6580
rect 23328 6528 23380 6580
rect 20384 6460 20436 6512
rect 21580 6460 21632 6512
rect 22132 6460 22184 6512
rect 23604 6460 23656 6512
rect 28480 6528 28532 6580
rect 28940 6528 28992 6580
rect 28664 6460 28716 6512
rect 28848 6503 28900 6512
rect 28848 6469 28857 6503
rect 28857 6469 28891 6503
rect 28891 6469 28900 6503
rect 28848 6460 28900 6469
rect 18870 6358 18922 6410
rect 18934 6358 18986 6410
rect 18998 6358 19050 6410
rect 19062 6358 19114 6410
rect 19126 6358 19178 6410
rect 880 6299 932 6308
rect 880 6265 889 6299
rect 889 6265 923 6299
rect 923 6265 932 6299
rect 880 6256 932 6265
rect 8700 6256 8752 6308
rect 9160 6256 9212 6308
rect 11276 6256 11328 6308
rect 12196 6256 12248 6308
rect 15232 6299 15284 6308
rect 15232 6265 15241 6299
rect 15241 6265 15275 6299
rect 15275 6265 15284 6299
rect 15232 6256 15284 6265
rect 24248 6299 24300 6308
rect 24248 6265 24257 6299
rect 24257 6265 24291 6299
rect 24291 6265 24300 6299
rect 24248 6256 24300 6265
rect 28020 6256 28072 6308
rect 29216 6299 29268 6308
rect 29216 6265 29225 6299
rect 29225 6265 29259 6299
rect 29259 6265 29268 6299
rect 29216 6256 29268 6265
rect 696 6188 748 6240
rect 3364 6188 3416 6240
rect 3088 6120 3140 6172
rect 4376 6188 4428 6240
rect 10356 6188 10408 6240
rect 21580 6188 21632 6240
rect 29308 6188 29360 6240
rect 6768 6163 6820 6172
rect 6768 6129 6777 6163
rect 6777 6129 6811 6163
rect 6811 6129 6820 6163
rect 6768 6120 6820 6129
rect 9528 6120 9580 6172
rect 13208 6163 13260 6172
rect 13208 6129 13217 6163
rect 13217 6129 13251 6163
rect 13251 6129 13260 6163
rect 13208 6120 13260 6129
rect 14772 6120 14824 6172
rect 15968 6120 16020 6172
rect 16152 6120 16204 6172
rect 18268 6163 18320 6172
rect 18268 6129 18277 6163
rect 18277 6129 18311 6163
rect 18311 6129 18320 6163
rect 18268 6120 18320 6129
rect 19464 6120 19516 6172
rect 19832 6120 19884 6172
rect 20568 6163 20620 6172
rect 20568 6129 20577 6163
rect 20577 6129 20611 6163
rect 20611 6129 20620 6163
rect 20568 6120 20620 6129
rect 26640 6120 26692 6172
rect 27744 6163 27796 6172
rect 27744 6129 27753 6163
rect 27753 6129 27787 6163
rect 27787 6129 27796 6163
rect 27744 6120 27796 6129
rect 28204 6120 28256 6172
rect 1800 6052 1852 6104
rect 2168 6052 2220 6104
rect 3916 6095 3968 6104
rect 3916 6061 3925 6095
rect 3925 6061 3959 6095
rect 3959 6061 3968 6095
rect 3916 6052 3968 6061
rect 5664 6095 5716 6104
rect 5664 6061 5673 6095
rect 5673 6061 5707 6095
rect 5707 6061 5716 6095
rect 5664 6052 5716 6061
rect 6584 6052 6636 6104
rect 8424 6052 8476 6104
rect 10724 6052 10776 6104
rect 10816 6095 10868 6104
rect 10816 6061 10825 6095
rect 10825 6061 10859 6095
rect 10859 6061 10868 6095
rect 13484 6095 13536 6104
rect 10816 6052 10868 6061
rect 13484 6061 13493 6095
rect 13493 6061 13527 6095
rect 13527 6061 13536 6095
rect 13484 6052 13536 6061
rect 16244 6052 16296 6104
rect 20384 6052 20436 6104
rect 21948 6095 22000 6104
rect 21948 6061 21957 6095
rect 21957 6061 21991 6095
rect 21991 6061 22000 6095
rect 21948 6052 22000 6061
rect 28296 6095 28348 6104
rect 28296 6061 28305 6095
rect 28305 6061 28339 6095
rect 28339 6061 28348 6095
rect 28296 6052 28348 6061
rect 12288 5984 12340 6036
rect 20200 5984 20252 6036
rect 27652 5984 27704 6036
rect 2996 5916 3048 5968
rect 5296 5916 5348 5968
rect 12380 5916 12432 5968
rect 18636 5916 18688 5968
rect 28848 5959 28900 5968
rect 28848 5925 28857 5959
rect 28857 5925 28891 5959
rect 28891 5925 28900 5959
rect 28848 5916 28900 5925
rect 3510 5814 3562 5866
rect 3574 5814 3626 5866
rect 3638 5814 3690 5866
rect 3702 5814 3754 5866
rect 3766 5814 3818 5866
rect 696 5619 748 5628
rect 696 5585 705 5619
rect 705 5585 739 5619
rect 739 5585 748 5619
rect 696 5576 748 5585
rect 2996 5712 3048 5764
rect 3088 5755 3140 5764
rect 3088 5721 3097 5755
rect 3097 5721 3131 5755
rect 3131 5721 3140 5755
rect 3916 5755 3968 5764
rect 3088 5712 3140 5721
rect 3916 5721 3925 5755
rect 3925 5721 3959 5755
rect 3959 5721 3968 5755
rect 3916 5712 3968 5721
rect 6952 5712 7004 5764
rect 11552 5712 11604 5764
rect 13208 5755 13260 5764
rect 13208 5721 13217 5755
rect 13217 5721 13251 5755
rect 13251 5721 13260 5755
rect 13208 5712 13260 5721
rect 14680 5712 14732 5764
rect 15784 5755 15836 5764
rect 15784 5721 15793 5755
rect 15793 5721 15827 5755
rect 15827 5721 15836 5755
rect 15784 5712 15836 5721
rect 15968 5755 16020 5764
rect 15968 5721 15977 5755
rect 15977 5721 16011 5755
rect 16011 5721 16020 5755
rect 15968 5712 16020 5721
rect 18268 5755 18320 5764
rect 18268 5721 18277 5755
rect 18277 5721 18311 5755
rect 18311 5721 18320 5755
rect 18268 5712 18320 5721
rect 19832 5755 19884 5764
rect 19832 5721 19841 5755
rect 19841 5721 19875 5755
rect 19875 5721 19884 5755
rect 19832 5712 19884 5721
rect 20568 5712 20620 5764
rect 21120 5712 21172 5764
rect 21856 5712 21908 5764
rect 24248 5755 24300 5764
rect 24248 5721 24257 5755
rect 24257 5721 24291 5755
rect 24291 5721 24300 5755
rect 24248 5712 24300 5721
rect 8424 5687 8476 5696
rect 8424 5653 8433 5687
rect 8433 5653 8467 5687
rect 8467 5653 8476 5687
rect 8424 5644 8476 5653
rect 9712 5576 9764 5628
rect 10540 5644 10592 5696
rect 11460 5687 11512 5696
rect 11460 5653 11469 5687
rect 11469 5653 11503 5687
rect 11503 5653 11512 5687
rect 11460 5644 11512 5653
rect 4468 5551 4520 5560
rect 4468 5517 4477 5551
rect 4477 5517 4511 5551
rect 4511 5517 4520 5551
rect 4468 5508 4520 5517
rect 4652 5551 4704 5560
rect 4652 5517 4661 5551
rect 4661 5517 4695 5551
rect 4695 5517 4704 5551
rect 4652 5508 4704 5517
rect 4836 5551 4888 5560
rect 4836 5517 4845 5551
rect 4845 5517 4879 5551
rect 4879 5517 4888 5551
rect 4836 5508 4888 5517
rect 6676 5508 6728 5560
rect 6768 5508 6820 5560
rect 7504 5508 7556 5560
rect 9252 5551 9304 5560
rect 9252 5517 9261 5551
rect 9261 5517 9295 5551
rect 9295 5517 9304 5551
rect 10080 5551 10132 5560
rect 9252 5508 9304 5517
rect 972 5483 1024 5492
rect 972 5449 981 5483
rect 981 5449 1015 5483
rect 1015 5449 1024 5483
rect 972 5440 1024 5449
rect 1432 5440 1484 5492
rect 5664 5440 5716 5492
rect 5940 5440 5992 5492
rect 9528 5440 9580 5492
rect 10080 5517 10089 5551
rect 10089 5517 10123 5551
rect 10123 5517 10132 5551
rect 10080 5508 10132 5517
rect 10356 5508 10408 5560
rect 10816 5508 10868 5560
rect 12196 5551 12248 5560
rect 12196 5517 12205 5551
rect 12205 5517 12239 5551
rect 12239 5517 12248 5551
rect 12196 5508 12248 5517
rect 12380 5551 12432 5560
rect 12380 5517 12389 5551
rect 12389 5517 12423 5551
rect 12423 5517 12432 5551
rect 12380 5508 12432 5517
rect 14864 5644 14916 5696
rect 20384 5687 20436 5696
rect 20384 5653 20393 5687
rect 20393 5653 20427 5687
rect 20427 5653 20436 5687
rect 20384 5644 20436 5653
rect 12932 5576 12984 5628
rect 13576 5576 13628 5628
rect 10908 5440 10960 5492
rect 14588 5508 14640 5560
rect 15784 5508 15836 5560
rect 19372 5576 19424 5628
rect 19464 5576 19516 5628
rect 21580 5644 21632 5696
rect 21672 5644 21724 5696
rect 20660 5576 20712 5628
rect 23420 5576 23472 5628
rect 25444 5712 25496 5764
rect 26640 5712 26692 5764
rect 28296 5712 28348 5764
rect 26180 5644 26232 5696
rect 27744 5644 27796 5696
rect 28204 5687 28256 5696
rect 28204 5653 28213 5687
rect 28213 5653 28247 5687
rect 28247 5653 28256 5687
rect 28204 5644 28256 5653
rect 26640 5576 26692 5628
rect 21212 5508 21264 5560
rect 21672 5508 21724 5560
rect 21856 5551 21908 5560
rect 21856 5517 21865 5551
rect 21865 5517 21899 5551
rect 21899 5517 21908 5551
rect 21856 5508 21908 5517
rect 4560 5372 4612 5424
rect 6584 5415 6636 5424
rect 6584 5381 6593 5415
rect 6593 5381 6627 5415
rect 6627 5381 6636 5415
rect 6584 5372 6636 5381
rect 9160 5415 9212 5424
rect 9160 5381 9169 5415
rect 9169 5381 9203 5415
rect 9203 5381 9212 5415
rect 9160 5372 9212 5381
rect 13484 5415 13536 5424
rect 13484 5381 13493 5415
rect 13493 5381 13527 5415
rect 13527 5381 13536 5415
rect 13484 5372 13536 5381
rect 13852 5372 13904 5424
rect 15140 5372 15192 5424
rect 15416 5415 15468 5424
rect 15416 5381 15425 5415
rect 15425 5381 15459 5415
rect 15459 5381 15468 5415
rect 15416 5372 15468 5381
rect 16244 5415 16296 5424
rect 16244 5381 16253 5415
rect 16253 5381 16287 5415
rect 16287 5381 16296 5415
rect 16244 5372 16296 5381
rect 18636 5372 18688 5424
rect 19280 5372 19332 5424
rect 20660 5415 20712 5424
rect 20660 5381 20669 5415
rect 20669 5381 20703 5415
rect 20703 5381 20712 5415
rect 20660 5372 20712 5381
rect 20936 5415 20988 5424
rect 20936 5381 20945 5415
rect 20945 5381 20979 5415
rect 20979 5381 20988 5415
rect 20936 5372 20988 5381
rect 24892 5508 24944 5560
rect 26548 5508 26600 5560
rect 27100 5440 27152 5492
rect 28204 5440 28256 5492
rect 24800 5415 24852 5424
rect 24800 5381 24809 5415
rect 24809 5381 24843 5415
rect 24843 5381 24852 5415
rect 24800 5372 24852 5381
rect 26916 5372 26968 5424
rect 28756 5440 28808 5492
rect 29308 5483 29360 5492
rect 29308 5449 29317 5483
rect 29317 5449 29351 5483
rect 29351 5449 29360 5483
rect 29308 5440 29360 5449
rect 18870 5270 18922 5322
rect 18934 5270 18986 5322
rect 18998 5270 19050 5322
rect 19062 5270 19114 5322
rect 19126 5270 19178 5322
rect 880 5211 932 5220
rect 880 5177 889 5211
rect 889 5177 923 5211
rect 923 5177 932 5211
rect 880 5168 932 5177
rect 1432 5168 1484 5220
rect 4376 5168 4428 5220
rect 9528 5211 9580 5220
rect 9528 5177 9537 5211
rect 9537 5177 9571 5211
rect 9571 5177 9580 5211
rect 9528 5168 9580 5177
rect 9712 5211 9764 5220
rect 9712 5177 9721 5211
rect 9721 5177 9755 5211
rect 9755 5177 9764 5211
rect 9712 5168 9764 5177
rect 972 5100 1024 5152
rect 4836 5100 4888 5152
rect 8148 5100 8200 5152
rect 1616 5032 1668 5084
rect 2168 5032 2220 5084
rect 3272 5032 3324 5084
rect 4008 5032 4060 5084
rect 4744 5032 4796 5084
rect 7320 5075 7372 5084
rect 7320 5041 7329 5075
rect 7329 5041 7363 5075
rect 7363 5041 7372 5075
rect 7320 5032 7372 5041
rect 7504 5075 7556 5084
rect 7504 5041 7513 5075
rect 7513 5041 7547 5075
rect 7547 5041 7556 5075
rect 7504 5032 7556 5041
rect 11276 5100 11328 5152
rect 16888 5100 16940 5152
rect 20752 5168 20804 5220
rect 20936 5211 20988 5220
rect 20936 5177 20945 5211
rect 20945 5177 20979 5211
rect 20979 5177 20988 5211
rect 20936 5168 20988 5177
rect 17624 5100 17676 5152
rect 9804 5032 9856 5084
rect 10908 5075 10960 5084
rect 10908 5041 10917 5075
rect 10917 5041 10951 5075
rect 10951 5041 10960 5075
rect 10908 5032 10960 5041
rect 15416 5075 15468 5084
rect 15416 5041 15425 5075
rect 15425 5041 15459 5075
rect 15459 5041 15468 5075
rect 15416 5032 15468 5041
rect 15876 5075 15928 5084
rect 1984 4964 2036 5016
rect 2352 5007 2404 5016
rect 2352 4973 2361 5007
rect 2361 4973 2395 5007
rect 2395 4973 2404 5007
rect 2352 4964 2404 4973
rect 2904 4964 2956 5016
rect 3364 4896 3416 4948
rect 4008 4896 4060 4948
rect 4560 5007 4612 5016
rect 4560 4973 4569 5007
rect 4569 4973 4603 5007
rect 4603 4973 4612 5007
rect 9160 5007 9212 5016
rect 4560 4964 4612 4973
rect 9160 4973 9169 5007
rect 9169 4973 9203 5007
rect 9203 4973 9212 5007
rect 9160 4964 9212 4973
rect 10724 4964 10776 5016
rect 11460 4964 11512 5016
rect 14680 4964 14732 5016
rect 15876 5041 15885 5075
rect 15885 5041 15919 5075
rect 15919 5041 15928 5075
rect 15876 5032 15928 5041
rect 16336 5075 16388 5084
rect 4652 4896 4704 4948
rect 15324 4896 15376 4948
rect 16336 5041 16354 5075
rect 16354 5041 16388 5075
rect 16336 5032 16388 5041
rect 18360 5075 18412 5084
rect 18360 5041 18369 5075
rect 18369 5041 18403 5075
rect 18403 5041 18412 5075
rect 18360 5032 18412 5041
rect 20660 5100 20712 5152
rect 21120 5100 21172 5152
rect 25260 5168 25312 5220
rect 25812 5168 25864 5220
rect 27652 5211 27704 5220
rect 27652 5177 27661 5211
rect 27661 5177 27695 5211
rect 27695 5177 27704 5211
rect 27652 5168 27704 5177
rect 28756 5168 28808 5220
rect 21764 5100 21816 5152
rect 22132 5100 22184 5152
rect 23420 5143 23472 5152
rect 23420 5109 23429 5143
rect 23429 5109 23463 5143
rect 23463 5109 23472 5143
rect 23420 5100 23472 5109
rect 24432 5100 24484 5152
rect 29124 5100 29176 5152
rect 19832 5032 19884 5084
rect 21396 5075 21448 5084
rect 21396 5041 21405 5075
rect 21405 5041 21439 5075
rect 21439 5041 21448 5075
rect 21396 5032 21448 5041
rect 24248 5075 24300 5084
rect 24248 5041 24257 5075
rect 24257 5041 24291 5075
rect 24291 5041 24300 5075
rect 24248 5032 24300 5041
rect 27100 5075 27152 5084
rect 27100 5041 27109 5075
rect 27109 5041 27143 5075
rect 27143 5041 27152 5075
rect 27100 5032 27152 5041
rect 28020 5032 28072 5084
rect 17072 4964 17124 5016
rect 18544 4964 18596 5016
rect 18636 4964 18688 5016
rect 24432 5007 24484 5016
rect 24432 4973 24441 5007
rect 24441 4973 24475 5007
rect 24475 4973 24484 5007
rect 24432 4964 24484 4973
rect 27284 5007 27336 5016
rect 27284 4973 27293 5007
rect 27293 4973 27327 5007
rect 27327 4973 27336 5007
rect 27284 4964 27336 4973
rect 28940 4964 28992 5016
rect 4468 4828 4520 4880
rect 4928 4828 4980 4880
rect 10080 4828 10132 4880
rect 12380 4828 12432 4880
rect 15140 4828 15192 4880
rect 18268 4828 18320 4880
rect 21212 4828 21264 4880
rect 3510 4726 3562 4778
rect 3574 4726 3626 4778
rect 3638 4726 3690 4778
rect 3702 4726 3754 4778
rect 3766 4726 3818 4778
rect 1616 4667 1668 4676
rect 1616 4633 1625 4667
rect 1625 4633 1659 4667
rect 1659 4633 1668 4667
rect 1616 4624 1668 4633
rect 1984 4624 2036 4676
rect 2168 4624 2220 4676
rect 4744 4667 4796 4676
rect 4744 4633 4753 4667
rect 4753 4633 4787 4667
rect 4787 4633 4796 4667
rect 4744 4624 4796 4633
rect 4928 4667 4980 4676
rect 4928 4633 4937 4667
rect 4937 4633 4971 4667
rect 4971 4633 4980 4667
rect 4928 4624 4980 4633
rect 7504 4667 7556 4676
rect 7504 4633 7513 4667
rect 7513 4633 7547 4667
rect 7547 4633 7556 4667
rect 7504 4624 7556 4633
rect 8148 4624 8200 4676
rect 9160 4624 9212 4676
rect 4560 4556 4612 4608
rect 5940 4556 5992 4608
rect 6584 4420 6636 4472
rect 9712 4624 9764 4676
rect 10448 4624 10500 4676
rect 10908 4667 10960 4676
rect 10908 4633 10917 4667
rect 10917 4633 10951 4667
rect 10951 4633 10960 4667
rect 10908 4624 10960 4633
rect 11276 4624 11328 4676
rect 11920 4624 11972 4676
rect 15324 4667 15376 4676
rect 9804 4599 9856 4608
rect 9804 4565 9813 4599
rect 9813 4565 9847 4599
rect 9847 4565 9856 4599
rect 9804 4556 9856 4565
rect 10540 4556 10592 4608
rect 15324 4633 15333 4667
rect 15333 4633 15367 4667
rect 15367 4633 15376 4667
rect 15324 4624 15376 4633
rect 15876 4667 15928 4676
rect 15876 4633 15885 4667
rect 15885 4633 15919 4667
rect 15919 4633 15928 4667
rect 15876 4624 15928 4633
rect 16888 4667 16940 4676
rect 16888 4633 16897 4667
rect 16897 4633 16931 4667
rect 16931 4633 16940 4667
rect 16888 4624 16940 4633
rect 18636 4624 18688 4676
rect 18728 4624 18780 4676
rect 21212 4624 21264 4676
rect 21764 4667 21816 4676
rect 21764 4633 21773 4667
rect 21773 4633 21807 4667
rect 21807 4633 21816 4667
rect 21764 4624 21816 4633
rect 24248 4667 24300 4676
rect 24248 4633 24257 4667
rect 24257 4633 24291 4667
rect 24291 4633 24300 4667
rect 24248 4624 24300 4633
rect 27100 4667 27152 4676
rect 27100 4633 27109 4667
rect 27109 4633 27143 4667
rect 27143 4633 27152 4667
rect 27100 4624 27152 4633
rect 28940 4667 28992 4676
rect 28940 4633 28949 4667
rect 28949 4633 28983 4667
rect 28983 4633 28992 4667
rect 28940 4624 28992 4633
rect 14588 4599 14640 4608
rect 14588 4565 14597 4599
rect 14597 4565 14631 4599
rect 14631 4565 14640 4599
rect 14588 4556 14640 4565
rect 14680 4599 14732 4608
rect 14680 4565 14689 4599
rect 14689 4565 14723 4599
rect 14723 4565 14732 4599
rect 14680 4556 14732 4565
rect 15232 4556 15284 4608
rect 17624 4599 17676 4608
rect 17624 4565 17633 4599
rect 17633 4565 17667 4599
rect 17667 4565 17676 4599
rect 17624 4556 17676 4565
rect 18176 4599 18228 4608
rect 18176 4565 18185 4599
rect 18185 4565 18219 4599
rect 18219 4565 18228 4599
rect 18176 4556 18228 4565
rect 18544 4556 18596 4608
rect 20660 4556 20712 4608
rect 11092 4488 11144 4540
rect 11920 4488 11972 4540
rect 14404 4488 14456 4540
rect 21120 4488 21172 4540
rect 21396 4488 21448 4540
rect 10172 4420 10224 4472
rect 12288 4420 12340 4472
rect 14496 4420 14548 4472
rect 3272 4284 3324 4336
rect 8976 4352 9028 4404
rect 11736 4352 11788 4404
rect 15692 4463 15744 4472
rect 15692 4429 15701 4463
rect 15701 4429 15735 4463
rect 15735 4429 15744 4463
rect 15692 4420 15744 4429
rect 16060 4420 16112 4472
rect 18360 4463 18412 4472
rect 18360 4429 18369 4463
rect 18369 4429 18403 4463
rect 18403 4429 18412 4463
rect 18360 4420 18412 4429
rect 6400 4327 6452 4336
rect 6400 4293 6409 4327
rect 6409 4293 6443 4327
rect 6443 4293 6452 4327
rect 6400 4284 6452 4293
rect 6584 4284 6636 4336
rect 7136 4284 7188 4336
rect 7320 4284 7372 4336
rect 7504 4284 7556 4336
rect 10724 4284 10776 4336
rect 11184 4327 11236 4336
rect 11184 4293 11193 4327
rect 11193 4293 11227 4327
rect 11227 4293 11236 4327
rect 11184 4284 11236 4293
rect 13392 4284 13444 4336
rect 14404 4327 14456 4336
rect 14404 4293 14413 4327
rect 14413 4293 14447 4327
rect 14447 4293 14456 4327
rect 14404 4284 14456 4293
rect 15048 4284 15100 4336
rect 18636 4420 18688 4472
rect 16336 4284 16388 4336
rect 28020 4420 28072 4472
rect 20568 4352 20620 4404
rect 28756 4395 28808 4404
rect 28756 4361 28765 4395
rect 28765 4361 28799 4395
rect 28799 4361 28808 4395
rect 28756 4352 28808 4361
rect 21028 4284 21080 4336
rect 21580 4284 21632 4336
rect 24064 4284 24116 4336
rect 24432 4327 24484 4336
rect 24432 4293 24441 4327
rect 24441 4293 24475 4327
rect 24475 4293 24484 4327
rect 24432 4284 24484 4293
rect 27284 4327 27336 4336
rect 27284 4293 27293 4327
rect 27293 4293 27327 4327
rect 27327 4293 27336 4327
rect 27284 4284 27336 4293
rect 28664 4327 28716 4336
rect 28664 4293 28673 4327
rect 28673 4293 28707 4327
rect 28707 4293 28716 4327
rect 28664 4284 28716 4293
rect 18870 4182 18922 4234
rect 18934 4182 18986 4234
rect 18998 4182 19050 4234
rect 19062 4182 19114 4234
rect 19126 4182 19178 4234
rect 1248 4123 1300 4132
rect 1248 4089 1257 4123
rect 1257 4089 1291 4123
rect 1291 4089 1300 4123
rect 1248 4080 1300 4089
rect 6400 4080 6452 4132
rect 9436 4080 9488 4132
rect 11000 4080 11052 4132
rect 13852 4123 13904 4132
rect 13852 4089 13861 4123
rect 13861 4089 13895 4123
rect 13895 4089 13904 4123
rect 13852 4080 13904 4089
rect 15416 4080 15468 4132
rect 18176 4080 18228 4132
rect 24800 4080 24852 4132
rect 25168 4123 25220 4132
rect 4652 4012 4704 4064
rect 5480 4012 5532 4064
rect 3916 3944 3968 3996
rect 5664 3944 5716 3996
rect 7596 4012 7648 4064
rect 5940 3987 5992 3996
rect 5940 3953 5949 3987
rect 5949 3953 5983 3987
rect 5983 3953 5992 3987
rect 5940 3944 5992 3953
rect 6952 3987 7004 3996
rect 6952 3953 6961 3987
rect 6961 3953 6995 3987
rect 6995 3953 7004 3987
rect 6952 3944 7004 3953
rect 7136 3987 7188 3996
rect 7136 3953 7145 3987
rect 7145 3953 7179 3987
rect 7179 3953 7188 3987
rect 7136 3944 7188 3953
rect 12380 4012 12432 4064
rect 16796 4012 16848 4064
rect 17348 4012 17400 4064
rect 12012 3987 12064 3996
rect 12012 3953 12021 3987
rect 12021 3953 12055 3987
rect 12055 3953 12064 3987
rect 12012 3944 12064 3953
rect 14956 3944 15008 3996
rect 17900 3987 17952 3996
rect 17900 3953 17909 3987
rect 17909 3953 17943 3987
rect 17943 3953 17952 3987
rect 17900 3944 17952 3953
rect 18360 4012 18412 4064
rect 25168 4089 25177 4123
rect 25177 4089 25211 4123
rect 25211 4089 25220 4123
rect 25168 4080 25220 4089
rect 28020 4080 28072 4132
rect 21672 3987 21724 3996
rect 21672 3953 21681 3987
rect 21681 3953 21715 3987
rect 21715 3953 21724 3987
rect 21672 3944 21724 3953
rect 21856 3944 21908 3996
rect 23880 3944 23932 3996
rect 24064 3987 24116 3996
rect 24064 3953 24073 3987
rect 24073 3953 24107 3987
rect 24107 3953 24116 3987
rect 24064 3944 24116 3953
rect 26180 4012 26232 4064
rect 3272 3876 3324 3928
rect 11736 3919 11788 3928
rect 11736 3885 11745 3919
rect 11745 3885 11779 3919
rect 11779 3885 11788 3919
rect 11736 3876 11788 3885
rect 5388 3851 5440 3860
rect 5388 3817 5397 3851
rect 5397 3817 5431 3851
rect 5431 3817 5440 3851
rect 5388 3808 5440 3817
rect 9160 3808 9212 3860
rect 10172 3808 10224 3860
rect 10632 3808 10684 3860
rect 11644 3808 11696 3860
rect 14404 3876 14456 3928
rect 15692 3876 15744 3928
rect 17808 3919 17860 3928
rect 17808 3885 17817 3919
rect 17817 3885 17851 3919
rect 17851 3885 17860 3919
rect 17808 3876 17860 3885
rect 14496 3808 14548 3860
rect 16060 3808 16112 3860
rect 17532 3808 17584 3860
rect 20476 3876 20528 3928
rect 21488 3919 21540 3928
rect 21488 3885 21497 3919
rect 21497 3885 21531 3919
rect 21531 3885 21540 3919
rect 21488 3876 21540 3885
rect 19188 3808 19240 3860
rect 21028 3808 21080 3860
rect 22224 3876 22276 3928
rect 23788 3919 23840 3928
rect 23788 3885 23797 3919
rect 23797 3885 23831 3919
rect 23831 3885 23840 3919
rect 23788 3876 23840 3885
rect 23144 3808 23196 3860
rect 26088 3944 26140 3996
rect 28664 4080 28716 4132
rect 29124 4012 29176 4064
rect 28756 3919 28808 3928
rect 28756 3885 28765 3919
rect 28765 3885 28799 3919
rect 28799 3885 28808 3919
rect 28756 3876 28808 3885
rect 2352 3783 2404 3792
rect 2352 3749 2361 3783
rect 2361 3749 2395 3783
rect 2395 3749 2404 3783
rect 2352 3740 2404 3749
rect 2904 3740 2956 3792
rect 3364 3740 3416 3792
rect 11276 3783 11328 3792
rect 11276 3749 11285 3783
rect 11285 3749 11319 3783
rect 11319 3749 11328 3783
rect 11276 3740 11328 3749
rect 18912 3783 18964 3792
rect 18912 3749 18921 3783
rect 18921 3749 18955 3783
rect 18955 3749 18964 3783
rect 18912 3740 18964 3749
rect 21304 3783 21356 3792
rect 21304 3749 21313 3783
rect 21313 3749 21347 3783
rect 21347 3749 21356 3783
rect 21304 3740 21356 3749
rect 23328 3783 23380 3792
rect 23328 3749 23337 3783
rect 23337 3749 23371 3783
rect 23371 3749 23380 3783
rect 23328 3740 23380 3749
rect 30504 3783 30556 3792
rect 30504 3749 30513 3783
rect 30513 3749 30547 3783
rect 30547 3749 30556 3783
rect 30504 3740 30556 3749
rect 3510 3638 3562 3690
rect 3574 3638 3626 3690
rect 3638 3638 3690 3690
rect 3702 3638 3754 3690
rect 3766 3638 3818 3690
rect 1248 3579 1300 3588
rect 1248 3545 1257 3579
rect 1257 3545 1291 3579
rect 1291 3545 1300 3579
rect 1248 3536 1300 3545
rect 3916 3536 3968 3588
rect 4376 3536 4428 3588
rect 5388 3579 5440 3588
rect 5388 3545 5397 3579
rect 5397 3545 5431 3579
rect 5431 3545 5440 3579
rect 5388 3536 5440 3545
rect 5480 3579 5532 3588
rect 5480 3545 5489 3579
rect 5489 3545 5523 3579
rect 5523 3545 5532 3579
rect 5480 3536 5532 3545
rect 5664 3536 5716 3588
rect 6952 3579 7004 3588
rect 6952 3545 6961 3579
rect 6961 3545 6995 3579
rect 6995 3545 7004 3579
rect 6952 3536 7004 3545
rect 7136 3579 7188 3588
rect 7136 3545 7145 3579
rect 7145 3545 7179 3579
rect 7179 3545 7188 3579
rect 7136 3536 7188 3545
rect 7596 3536 7648 3588
rect 11276 3579 11328 3588
rect 11276 3545 11285 3579
rect 11285 3545 11319 3579
rect 11319 3545 11328 3579
rect 11276 3536 11328 3545
rect 14956 3536 15008 3588
rect 15508 3536 15560 3588
rect 16060 3579 16112 3588
rect 16060 3545 16069 3579
rect 16069 3545 16103 3579
rect 16103 3545 16112 3579
rect 16060 3536 16112 3545
rect 16796 3579 16848 3588
rect 16796 3545 16805 3579
rect 16805 3545 16839 3579
rect 16839 3545 16848 3579
rect 16796 3536 16848 3545
rect 18452 3536 18504 3588
rect 18912 3536 18964 3588
rect 20200 3536 20252 3588
rect 21028 3579 21080 3588
rect 21028 3545 21037 3579
rect 21037 3545 21071 3579
rect 21071 3545 21080 3579
rect 21028 3536 21080 3545
rect 21304 3579 21356 3588
rect 21304 3545 21313 3579
rect 21313 3545 21347 3579
rect 21347 3545 21356 3579
rect 21304 3536 21356 3545
rect 21856 3536 21908 3588
rect 23328 3579 23380 3588
rect 23328 3545 23337 3579
rect 23337 3545 23371 3579
rect 23371 3545 23380 3579
rect 23328 3536 23380 3545
rect 28756 3536 28808 3588
rect 5940 3468 5992 3520
rect 3364 3400 3416 3452
rect 2904 3375 2956 3384
rect 2904 3341 2913 3375
rect 2913 3341 2947 3375
rect 2947 3341 2956 3375
rect 2904 3332 2956 3341
rect 5848 3400 5900 3452
rect 12012 3468 12064 3520
rect 12380 3468 12432 3520
rect 13116 3468 13168 3520
rect 9896 3400 9948 3452
rect 1064 3264 1116 3316
rect 4376 3332 4428 3384
rect 3272 3196 3324 3248
rect 3916 3239 3968 3248
rect 3916 3205 3925 3239
rect 3925 3205 3959 3239
rect 3959 3205 3968 3239
rect 6032 3332 6084 3384
rect 10172 3400 10224 3452
rect 11736 3400 11788 3452
rect 13852 3468 13904 3520
rect 15416 3468 15468 3520
rect 17808 3468 17860 3520
rect 10356 3375 10408 3384
rect 10356 3341 10365 3375
rect 10365 3341 10399 3375
rect 10399 3341 10408 3375
rect 10356 3332 10408 3341
rect 8148 3264 8200 3316
rect 5664 3239 5716 3248
rect 3916 3196 3968 3205
rect 5664 3205 5673 3239
rect 5673 3205 5707 3239
rect 5707 3205 5716 3239
rect 5664 3196 5716 3205
rect 6032 3196 6084 3248
rect 7504 3196 7556 3248
rect 9252 3239 9304 3248
rect 9252 3205 9261 3239
rect 9261 3205 9295 3239
rect 9295 3205 9304 3239
rect 10540 3332 10592 3384
rect 12104 3332 12156 3384
rect 12288 3332 12340 3384
rect 12380 3375 12432 3384
rect 12380 3341 12389 3375
rect 12389 3341 12423 3375
rect 12423 3341 12432 3375
rect 12380 3332 12432 3341
rect 12932 3375 12984 3384
rect 12932 3341 12941 3375
rect 12941 3341 12975 3375
rect 12975 3341 12984 3375
rect 12932 3332 12984 3341
rect 11736 3264 11788 3316
rect 13484 3307 13536 3316
rect 13484 3273 13493 3307
rect 13493 3273 13527 3307
rect 13527 3273 13536 3307
rect 13484 3264 13536 3273
rect 14404 3375 14456 3384
rect 14404 3341 14413 3375
rect 14413 3341 14447 3375
rect 14447 3341 14456 3375
rect 18636 3443 18688 3452
rect 18636 3409 18645 3443
rect 18645 3409 18679 3443
rect 18679 3409 18688 3443
rect 18636 3400 18688 3409
rect 14772 3375 14824 3384
rect 14404 3332 14456 3341
rect 14772 3341 14781 3375
rect 14781 3341 14815 3375
rect 14815 3341 14824 3375
rect 14772 3332 14824 3341
rect 9252 3196 9304 3205
rect 11644 3196 11696 3248
rect 11828 3239 11880 3248
rect 11828 3205 11837 3239
rect 11837 3205 11871 3239
rect 11871 3205 11880 3239
rect 11828 3196 11880 3205
rect 13576 3239 13628 3248
rect 13576 3205 13585 3239
rect 13585 3205 13619 3239
rect 13619 3205 13628 3239
rect 15692 3332 15744 3384
rect 16980 3375 17032 3384
rect 16980 3341 16989 3375
rect 16989 3341 17023 3375
rect 17023 3341 17032 3375
rect 16980 3332 17032 3341
rect 17900 3332 17952 3384
rect 21212 3468 21264 3520
rect 24892 3511 24944 3520
rect 24892 3477 24901 3511
rect 24901 3477 24935 3511
rect 24935 3477 24944 3511
rect 24892 3468 24944 3477
rect 25168 3468 25220 3520
rect 27284 3468 27336 3520
rect 29216 3468 29268 3520
rect 19188 3443 19240 3452
rect 19188 3409 19197 3443
rect 19197 3409 19231 3443
rect 19231 3409 19240 3443
rect 19188 3400 19240 3409
rect 21488 3443 21540 3452
rect 19280 3332 19332 3384
rect 21488 3409 21497 3443
rect 21497 3409 21531 3443
rect 21531 3409 21540 3443
rect 21488 3400 21540 3409
rect 21856 3400 21908 3452
rect 23788 3400 23840 3452
rect 15048 3264 15100 3316
rect 17348 3239 17400 3248
rect 13576 3196 13628 3205
rect 17348 3205 17357 3239
rect 17357 3205 17391 3239
rect 17391 3205 17400 3239
rect 17348 3196 17400 3205
rect 17532 3239 17584 3248
rect 17532 3205 17541 3239
rect 17541 3205 17575 3239
rect 17575 3205 17584 3239
rect 17532 3196 17584 3205
rect 18636 3264 18688 3316
rect 24064 3332 24116 3384
rect 25536 3375 25588 3384
rect 25536 3341 25545 3375
rect 25545 3341 25579 3375
rect 25579 3341 25588 3375
rect 25536 3332 25588 3341
rect 26088 3375 26140 3384
rect 21672 3264 21724 3316
rect 23144 3239 23196 3248
rect 23144 3205 23153 3239
rect 23153 3205 23187 3239
rect 23187 3205 23196 3239
rect 23144 3196 23196 3205
rect 23420 3239 23472 3248
rect 23420 3205 23429 3239
rect 23429 3205 23463 3239
rect 23463 3205 23472 3239
rect 23420 3196 23472 3205
rect 23880 3239 23932 3248
rect 23880 3205 23889 3239
rect 23889 3205 23923 3239
rect 23923 3205 23932 3239
rect 24800 3239 24852 3248
rect 23880 3196 23932 3205
rect 24800 3205 24809 3239
rect 24809 3205 24843 3239
rect 24843 3205 24852 3239
rect 26088 3341 26097 3375
rect 26097 3341 26131 3375
rect 26131 3341 26140 3375
rect 26088 3332 26140 3341
rect 26548 3375 26600 3384
rect 26548 3341 26557 3375
rect 26557 3341 26591 3375
rect 26591 3341 26600 3375
rect 26548 3332 26600 3341
rect 28296 3332 28348 3384
rect 29216 3375 29268 3384
rect 29216 3341 29225 3375
rect 29225 3341 29259 3375
rect 29259 3341 29268 3375
rect 29216 3332 29268 3341
rect 29308 3332 29360 3384
rect 29584 3375 29636 3384
rect 29584 3341 29593 3375
rect 29593 3341 29627 3375
rect 29627 3341 29636 3375
rect 29584 3332 29636 3341
rect 30504 3332 30556 3384
rect 28296 3239 28348 3248
rect 24800 3196 24852 3205
rect 28296 3205 28305 3239
rect 28305 3205 28339 3239
rect 28339 3205 28348 3239
rect 28296 3196 28348 3205
rect 28756 3196 28808 3248
rect 29584 3196 29636 3248
rect 18870 3094 18922 3146
rect 18934 3094 18986 3146
rect 18998 3094 19050 3146
rect 19062 3094 19114 3146
rect 19126 3094 19178 3146
rect 1064 3035 1116 3044
rect 1064 3001 1073 3035
rect 1073 3001 1107 3035
rect 1107 3001 1116 3035
rect 1064 2992 1116 3001
rect 3364 3035 3416 3044
rect 3364 3001 3373 3035
rect 3373 3001 3407 3035
rect 3407 3001 3416 3035
rect 3364 2992 3416 3001
rect 5664 2992 5716 3044
rect 8148 3035 8200 3044
rect 8148 3001 8157 3035
rect 8157 3001 8191 3035
rect 8191 3001 8200 3035
rect 8148 2992 8200 3001
rect 10356 2992 10408 3044
rect 11828 3035 11880 3044
rect 11828 3001 11837 3035
rect 11837 3001 11871 3035
rect 11871 3001 11880 3035
rect 11828 2992 11880 3001
rect 12012 2992 12064 3044
rect 13392 2992 13444 3044
rect 14772 2992 14824 3044
rect 17808 2992 17860 3044
rect 18176 2992 18228 3044
rect 5388 2924 5440 2976
rect 7504 2967 7556 2976
rect 7504 2933 7513 2967
rect 7513 2933 7547 2967
rect 7547 2933 7556 2967
rect 7504 2924 7556 2933
rect 11736 2967 11788 2976
rect 11736 2933 11745 2967
rect 11745 2933 11779 2967
rect 11779 2933 11788 2967
rect 11736 2924 11788 2933
rect 12104 2967 12156 2976
rect 12104 2933 12113 2967
rect 12113 2933 12147 2967
rect 12147 2933 12156 2967
rect 12104 2924 12156 2933
rect 13116 2967 13168 2976
rect 13116 2933 13125 2967
rect 13125 2933 13159 2967
rect 13159 2933 13168 2967
rect 13116 2924 13168 2933
rect 15508 2967 15560 2976
rect 15508 2933 15517 2967
rect 15517 2933 15551 2967
rect 15551 2933 15560 2967
rect 15508 2924 15560 2933
rect 17072 2967 17124 2976
rect 17072 2933 17081 2967
rect 17081 2933 17115 2967
rect 17115 2933 17124 2967
rect 17072 2924 17124 2933
rect 17900 2924 17952 2976
rect 21212 2992 21264 3044
rect 21580 2992 21632 3044
rect 21304 2924 21356 2976
rect 22224 2992 22276 3044
rect 23328 2992 23380 3044
rect 26180 3035 26232 3044
rect 26180 3001 26189 3035
rect 26189 3001 26223 3035
rect 26223 3001 26232 3035
rect 26180 2992 26232 3001
rect 26088 2967 26140 2976
rect 26088 2933 26097 2967
rect 26097 2933 26131 2967
rect 26131 2933 26140 2967
rect 26088 2924 26140 2933
rect 28756 2924 28808 2976
rect 3364 2856 3416 2908
rect 3916 2856 3968 2908
rect 4468 2899 4520 2908
rect 4468 2865 4477 2899
rect 4477 2865 4511 2899
rect 4511 2865 4520 2899
rect 4468 2856 4520 2865
rect 4652 2856 4704 2908
rect 6860 2856 6912 2908
rect 11092 2856 11144 2908
rect 11644 2856 11696 2908
rect 15692 2899 15744 2908
rect 15692 2865 15701 2899
rect 15701 2865 15735 2899
rect 15735 2865 15744 2899
rect 15692 2856 15744 2865
rect 16244 2856 16296 2908
rect 16888 2899 16940 2908
rect 16888 2865 16897 2899
rect 16897 2865 16931 2899
rect 16931 2865 16940 2899
rect 16888 2856 16940 2865
rect 17164 2899 17216 2908
rect 17164 2865 17173 2899
rect 17173 2865 17207 2899
rect 17207 2865 17216 2899
rect 17164 2856 17216 2865
rect 21120 2899 21172 2908
rect 4008 2788 4060 2840
rect 3916 2763 3968 2772
rect 3916 2729 3925 2763
rect 3925 2729 3959 2763
rect 3959 2729 3968 2763
rect 3916 2720 3968 2729
rect 6124 2788 6176 2840
rect 9712 2831 9764 2840
rect 9712 2797 9721 2831
rect 9721 2797 9755 2831
rect 9755 2797 9764 2831
rect 9712 2788 9764 2797
rect 9988 2831 10040 2840
rect 9988 2797 9997 2831
rect 9997 2797 10031 2831
rect 10031 2797 10040 2831
rect 9988 2788 10040 2797
rect 16060 2831 16112 2840
rect 16060 2797 16069 2831
rect 16069 2797 16103 2831
rect 16103 2797 16112 2831
rect 16060 2788 16112 2797
rect 21120 2865 21129 2899
rect 21129 2865 21163 2899
rect 21163 2865 21172 2899
rect 21120 2856 21172 2865
rect 26548 2856 26600 2908
rect 28020 2899 28072 2908
rect 28020 2865 28029 2899
rect 28029 2865 28063 2899
rect 28063 2865 28072 2899
rect 28020 2856 28072 2865
rect 23696 2788 23748 2840
rect 26824 2788 26876 2840
rect 28848 2788 28900 2840
rect 29308 2788 29360 2840
rect 1708 2652 1760 2704
rect 4560 2652 4612 2704
rect 13392 2695 13444 2704
rect 13392 2661 13401 2695
rect 13401 2661 13435 2695
rect 13435 2661 13444 2695
rect 13392 2652 13444 2661
rect 18452 2695 18504 2704
rect 18452 2661 18461 2695
rect 18461 2661 18495 2695
rect 18495 2661 18504 2695
rect 18452 2652 18504 2661
rect 18636 2652 18688 2704
rect 19096 2652 19148 2704
rect 19740 2652 19792 2704
rect 23604 2652 23656 2704
rect 25812 2695 25864 2704
rect 25812 2661 25821 2695
rect 25821 2661 25855 2695
rect 25855 2661 25864 2695
rect 25812 2652 25864 2661
rect 3510 2550 3562 2602
rect 3574 2550 3626 2602
rect 3638 2550 3690 2602
rect 3702 2550 3754 2602
rect 3766 2550 3818 2602
rect 1064 2448 1116 2500
rect 3364 2491 3416 2500
rect 3364 2457 3373 2491
rect 3373 2457 3407 2491
rect 3407 2457 3416 2491
rect 3364 2448 3416 2457
rect 3916 2448 3968 2500
rect 5388 2448 5440 2500
rect 6124 2491 6176 2500
rect 6124 2457 6133 2491
rect 6133 2457 6167 2491
rect 6167 2457 6176 2491
rect 6124 2448 6176 2457
rect 4468 2380 4520 2432
rect 6032 2380 6084 2432
rect 1708 2312 1760 2364
rect 972 2287 1024 2296
rect 972 2253 981 2287
rect 981 2253 1015 2287
rect 1015 2253 1024 2287
rect 972 2244 1024 2253
rect 1708 2176 1760 2228
rect 4008 2244 4060 2296
rect 4192 2312 4244 2364
rect 6860 2448 6912 2500
rect 9988 2448 10040 2500
rect 11828 2448 11880 2500
rect 13392 2448 13444 2500
rect 15508 2448 15560 2500
rect 16060 2448 16112 2500
rect 17164 2448 17216 2500
rect 11736 2380 11788 2432
rect 17072 2380 17124 2432
rect 19372 2448 19424 2500
rect 21212 2491 21264 2500
rect 21212 2457 21221 2491
rect 21221 2457 21255 2491
rect 21255 2457 21264 2491
rect 21212 2448 21264 2457
rect 21304 2448 21356 2500
rect 23236 2448 23288 2500
rect 24432 2448 24484 2500
rect 25444 2448 25496 2500
rect 21120 2380 21172 2432
rect 4100 2219 4152 2228
rect 4100 2185 4109 2219
rect 4109 2185 4143 2219
rect 4143 2185 4152 2219
rect 4100 2176 4152 2185
rect 4284 2244 4336 2296
rect 6768 2244 6820 2296
rect 4652 2176 4704 2228
rect 3272 2108 3324 2160
rect 7228 2108 7280 2160
rect 9252 2312 9304 2364
rect 13484 2312 13536 2364
rect 16888 2355 16940 2364
rect 16888 2321 16897 2355
rect 16897 2321 16931 2355
rect 16931 2321 16940 2355
rect 16888 2312 16940 2321
rect 8056 2287 8108 2296
rect 8056 2253 8065 2287
rect 8065 2253 8099 2287
rect 8099 2253 8108 2287
rect 8056 2244 8108 2253
rect 8148 2244 8200 2296
rect 10356 2244 10408 2296
rect 11184 2244 11236 2296
rect 18360 2312 18412 2364
rect 21028 2312 21080 2364
rect 9804 2176 9856 2228
rect 11092 2176 11144 2228
rect 11736 2108 11788 2160
rect 13484 2176 13536 2228
rect 18452 2244 18504 2296
rect 18544 2244 18596 2296
rect 19096 2244 19148 2296
rect 23328 2312 23380 2364
rect 23420 2244 23472 2296
rect 15692 2176 15744 2228
rect 18176 2176 18228 2228
rect 17532 2151 17584 2160
rect 17532 2117 17541 2151
rect 17541 2117 17575 2151
rect 17575 2117 17584 2151
rect 17532 2108 17584 2117
rect 19372 2176 19424 2228
rect 22500 2176 22552 2228
rect 23144 2219 23196 2228
rect 23144 2185 23153 2219
rect 23153 2185 23187 2219
rect 23187 2185 23196 2219
rect 23144 2176 23196 2185
rect 19464 2108 19516 2160
rect 20752 2151 20804 2160
rect 20752 2117 20761 2151
rect 20761 2117 20795 2151
rect 20795 2117 20804 2151
rect 20752 2108 20804 2117
rect 23328 2151 23380 2160
rect 23328 2117 23337 2151
rect 23337 2117 23371 2151
rect 23371 2117 23380 2151
rect 23328 2108 23380 2117
rect 24432 2176 24484 2228
rect 25812 2312 25864 2364
rect 26824 2355 26876 2364
rect 26824 2321 26833 2355
rect 26833 2321 26867 2355
rect 26867 2321 26876 2355
rect 26824 2312 26876 2321
rect 27284 2448 27336 2500
rect 28848 2448 28900 2500
rect 27468 2380 27520 2432
rect 28204 2380 28256 2432
rect 29584 2312 29636 2364
rect 27376 2287 27428 2296
rect 27376 2253 27385 2287
rect 27385 2253 27419 2287
rect 27419 2253 27428 2287
rect 27376 2244 27428 2253
rect 27744 2244 27796 2296
rect 28020 2244 28072 2296
rect 25628 2176 25680 2228
rect 27836 2176 27888 2228
rect 28388 2176 28440 2228
rect 29308 2176 29360 2228
rect 27744 2108 27796 2160
rect 18870 2006 18922 2058
rect 18934 2006 18986 2058
rect 18998 2006 19050 2058
rect 19062 2006 19114 2058
rect 19126 2006 19178 2058
rect 972 1904 1024 1956
rect 1156 1811 1208 1820
rect 1156 1777 1165 1811
rect 1165 1777 1199 1811
rect 1199 1777 1208 1811
rect 1156 1768 1208 1777
rect 1708 1904 1760 1956
rect 5572 1904 5624 1956
rect 8056 1904 8108 1956
rect 9712 1904 9764 1956
rect 10356 1904 10408 1956
rect 13576 1904 13628 1956
rect 16980 1947 17032 1956
rect 16980 1913 16989 1947
rect 16989 1913 17023 1947
rect 17023 1913 17032 1947
rect 16980 1904 17032 1913
rect 18360 1947 18412 1956
rect 18360 1913 18369 1947
rect 18369 1913 18403 1947
rect 18403 1913 18412 1947
rect 18360 1904 18412 1913
rect 18452 1904 18504 1956
rect 3916 1836 3968 1888
rect 4652 1836 4704 1888
rect 5848 1836 5900 1888
rect 6768 1811 6820 1820
rect 6768 1777 6777 1811
rect 6777 1777 6811 1811
rect 6811 1777 6820 1811
rect 6768 1768 6820 1777
rect 13116 1836 13168 1888
rect 13484 1879 13536 1888
rect 13484 1845 13493 1879
rect 13493 1845 13527 1879
rect 13527 1845 13536 1879
rect 13484 1836 13536 1845
rect 18636 1836 18688 1888
rect 11092 1768 11144 1820
rect 4560 1700 4612 1752
rect 6952 1743 7004 1752
rect 6952 1709 6961 1743
rect 6961 1709 6995 1743
rect 6995 1709 7004 1743
rect 6952 1700 7004 1709
rect 10080 1700 10132 1752
rect 11276 1700 11328 1752
rect 11736 1743 11788 1752
rect 11736 1709 11745 1743
rect 11745 1709 11779 1743
rect 11779 1709 11788 1743
rect 11736 1700 11788 1709
rect 13944 1700 13996 1752
rect 18452 1768 18504 1820
rect 18728 1811 18780 1820
rect 18728 1777 18737 1811
rect 18737 1777 18771 1811
rect 18771 1777 18780 1811
rect 18728 1768 18780 1777
rect 19096 1811 19148 1820
rect 19096 1777 19105 1811
rect 19105 1777 19139 1811
rect 19139 1777 19148 1811
rect 19096 1768 19148 1777
rect 20200 1768 20252 1820
rect 27376 1904 27428 1956
rect 21212 1836 21264 1888
rect 21764 1836 21816 1888
rect 23052 1768 23104 1820
rect 17348 1700 17400 1752
rect 18176 1700 18228 1752
rect 19464 1700 19516 1752
rect 20660 1743 20712 1752
rect 20660 1709 20669 1743
rect 20669 1709 20703 1743
rect 20703 1709 20712 1743
rect 20660 1700 20712 1709
rect 22040 1743 22092 1752
rect 22040 1709 22049 1743
rect 22049 1709 22083 1743
rect 22083 1709 22092 1743
rect 22040 1700 22092 1709
rect 22592 1700 22644 1752
rect 23696 1743 23748 1752
rect 23696 1709 23705 1743
rect 23705 1709 23739 1743
rect 23739 1709 23748 1743
rect 23696 1700 23748 1709
rect 23880 1811 23932 1820
rect 23880 1777 23889 1811
rect 23889 1777 23923 1811
rect 23923 1777 23932 1811
rect 23880 1768 23932 1777
rect 24064 1768 24116 1820
rect 24800 1768 24852 1820
rect 28204 1836 28256 1888
rect 27836 1811 27888 1820
rect 27836 1777 27845 1811
rect 27845 1777 27879 1811
rect 27879 1777 27888 1811
rect 27836 1768 27888 1777
rect 28020 1700 28072 1752
rect 18544 1632 18596 1684
rect 26548 1632 26600 1684
rect 2168 1607 2220 1616
rect 2168 1573 2177 1607
rect 2177 1573 2211 1607
rect 2211 1573 2220 1607
rect 2168 1564 2220 1573
rect 12748 1607 12800 1616
rect 12748 1573 12757 1607
rect 12757 1573 12791 1607
rect 12791 1573 12800 1607
rect 12748 1564 12800 1573
rect 15140 1607 15192 1616
rect 15140 1573 15149 1607
rect 15149 1573 15183 1607
rect 15183 1573 15192 1607
rect 15140 1564 15192 1573
rect 16612 1564 16664 1616
rect 23696 1564 23748 1616
rect 25996 1607 26048 1616
rect 25996 1573 26005 1607
rect 26005 1573 26039 1607
rect 26039 1573 26048 1607
rect 25996 1564 26048 1573
rect 27744 1564 27796 1616
rect 30780 1564 30832 1616
rect 3510 1462 3562 1514
rect 3574 1462 3626 1514
rect 3638 1462 3690 1514
rect 3702 1462 3754 1514
rect 3766 1462 3818 1514
rect 1156 1360 1208 1412
rect 3916 1360 3968 1412
rect 4652 1360 4704 1412
rect 6952 1360 7004 1412
rect 9804 1403 9856 1412
rect 9804 1369 9813 1403
rect 9813 1369 9847 1403
rect 9847 1369 9856 1403
rect 9804 1360 9856 1369
rect 10080 1403 10132 1412
rect 10080 1369 10089 1403
rect 10089 1369 10123 1403
rect 10123 1369 10132 1403
rect 10080 1360 10132 1369
rect 10356 1403 10408 1412
rect 10356 1369 10365 1403
rect 10365 1369 10399 1403
rect 10399 1369 10408 1403
rect 10356 1360 10408 1369
rect 18176 1403 18228 1412
rect 18176 1369 18185 1403
rect 18185 1369 18219 1403
rect 18219 1369 18228 1403
rect 18176 1360 18228 1369
rect 18452 1403 18504 1412
rect 18452 1369 18461 1403
rect 18461 1369 18495 1403
rect 18495 1369 18504 1403
rect 18452 1360 18504 1369
rect 18728 1403 18780 1412
rect 18728 1369 18737 1403
rect 18737 1369 18771 1403
rect 18771 1369 18780 1403
rect 18728 1360 18780 1369
rect 20660 1360 20712 1412
rect 21764 1360 21816 1412
rect 24064 1360 24116 1412
rect 24432 1360 24484 1412
rect 27468 1403 27520 1412
rect 27468 1369 27477 1403
rect 27477 1369 27511 1403
rect 27511 1369 27520 1403
rect 27468 1360 27520 1369
rect 27836 1403 27888 1412
rect 27836 1369 27845 1403
rect 27845 1369 27879 1403
rect 27879 1369 27888 1403
rect 27836 1360 27888 1369
rect 28020 1403 28072 1412
rect 28020 1369 28029 1403
rect 28029 1369 28063 1403
rect 28063 1369 28072 1403
rect 28020 1360 28072 1369
rect 5848 1292 5900 1344
rect 11736 1292 11788 1344
rect 18360 1335 18412 1344
rect 18360 1301 18369 1335
rect 18369 1301 18403 1335
rect 18403 1301 18412 1335
rect 18360 1292 18412 1301
rect 22592 1335 22644 1344
rect 4560 1267 4612 1276
rect 4560 1233 4569 1267
rect 4569 1233 4603 1267
rect 4603 1233 4612 1267
rect 4560 1224 4612 1233
rect 6768 1224 6820 1276
rect 19096 1224 19148 1276
rect 19648 1267 19700 1276
rect 19648 1233 19657 1267
rect 19657 1233 19691 1267
rect 19691 1233 19700 1267
rect 19648 1224 19700 1233
rect 22592 1301 22601 1335
rect 22601 1301 22635 1335
rect 22635 1301 22644 1335
rect 22592 1292 22644 1301
rect 21212 1224 21264 1276
rect 23328 1292 23380 1344
rect 24800 1292 24852 1344
rect 27744 1335 27796 1344
rect 23696 1267 23748 1276
rect 23696 1233 23705 1267
rect 23705 1233 23739 1267
rect 23739 1233 23748 1267
rect 23696 1224 23748 1233
rect 27744 1301 27753 1335
rect 27753 1301 27787 1335
rect 27787 1301 27796 1335
rect 27744 1292 27796 1301
rect 20200 1199 20252 1208
rect 20200 1165 20209 1199
rect 20209 1165 20243 1199
rect 20243 1165 20252 1199
rect 20200 1156 20252 1165
rect 4468 1088 4520 1140
rect 19280 1088 19332 1140
rect 22040 1156 22092 1208
rect 23420 1199 23472 1208
rect 23420 1165 23429 1199
rect 23429 1165 23463 1199
rect 23463 1165 23472 1199
rect 23420 1156 23472 1165
rect 24432 1088 24484 1140
rect 2168 1020 2220 1072
rect 3180 1020 3232 1072
rect 11460 1020 11512 1072
rect 12748 1020 12800 1072
rect 15140 1020 15192 1072
rect 15508 1020 15560 1072
rect 16612 1063 16664 1072
rect 16612 1029 16621 1063
rect 16621 1029 16655 1063
rect 16655 1029 16664 1063
rect 16612 1020 16664 1029
rect 23052 1063 23104 1072
rect 23052 1029 23061 1063
rect 23061 1029 23095 1063
rect 23095 1029 23104 1063
rect 23052 1020 23104 1029
rect 23788 1020 23840 1072
rect 25996 1020 26048 1072
rect 18870 918 18922 970
rect 18934 918 18986 970
rect 18998 918 19050 970
rect 19062 918 19114 970
rect 19126 918 19178 970
rect 20200 816 20252 868
rect 23696 859 23748 868
rect 23696 825 23705 859
rect 23705 825 23739 859
rect 23739 825 23748 859
rect 23696 816 23748 825
rect 23880 859 23932 868
rect 23880 825 23889 859
rect 23889 825 23923 859
rect 23923 825 23932 859
rect 23880 816 23932 825
rect 19648 748 19700 800
rect 23420 748 23472 800
rect 21028 476 21080 528
rect 23052 476 23104 528
rect 3510 374 3562 426
rect 3574 374 3626 426
rect 3638 374 3690 426
rect 3702 374 3754 426
rect 3766 374 3818 426
<< metal2 >>
rect 1126 31664 1238 32088
rect 2598 31664 2710 32088
rect 3886 31664 3998 32088
rect 5358 31664 5470 32088
rect 6646 31664 6758 32088
rect 8118 31690 8230 32088
rect 7516 31664 8230 31690
rect 9406 31664 9518 32088
rect 10878 31664 10990 32088
rect 12166 31664 12278 32088
rect 13638 31664 13750 32088
rect 14926 31664 15038 32088
rect 16398 31664 16510 32088
rect 17686 31664 17798 32088
rect 19158 31664 19270 32088
rect 20446 31664 20558 32088
rect 21918 31690 22030 32088
rect 21776 31664 22030 31690
rect 23206 31664 23318 32088
rect 418 30960 474 30969
rect 418 30895 474 30904
rect 432 30250 460 30895
rect 1168 30658 1196 31664
rect 2640 30726 2668 31664
rect 3504 30892 3824 30912
rect 3504 30890 3516 30892
rect 3572 30890 3596 30892
rect 3652 30890 3676 30892
rect 3732 30890 3756 30892
rect 3812 30890 3824 30892
rect 3504 30838 3510 30890
rect 3572 30838 3574 30890
rect 3754 30838 3756 30890
rect 3818 30838 3824 30890
rect 3504 30836 3516 30838
rect 3572 30836 3596 30838
rect 3652 30836 3676 30838
rect 3732 30836 3756 30838
rect 3812 30836 3824 30838
rect 3504 30816 3824 30836
rect 2628 30720 2680 30726
rect 2628 30662 2680 30668
rect 1156 30652 1208 30658
rect 1156 30594 1208 30600
rect 3928 30454 3956 31664
rect 5400 30640 5428 31664
rect 5400 30612 5520 30640
rect 4008 30584 4060 30590
rect 4008 30526 4060 30532
rect 3916 30448 3968 30454
rect 3916 30390 3968 30396
rect 420 30244 472 30250
rect 420 30186 472 30192
rect 4020 30182 4048 30526
rect 5020 30516 5072 30522
rect 5020 30458 5072 30464
rect 5388 30516 5440 30522
rect 5388 30458 5440 30464
rect 4008 30176 4060 30182
rect 4008 30118 4060 30124
rect 4468 30176 4520 30182
rect 4468 30118 4520 30124
rect 3180 30040 3232 30046
rect 3180 29982 3232 29988
rect 1156 29972 1208 29978
rect 1156 29914 1208 29920
rect 1168 29434 1196 29914
rect 1248 29904 1300 29910
rect 1248 29846 1300 29852
rect 1260 29570 1288 29846
rect 3192 29706 3220 29982
rect 3504 29804 3824 29824
rect 3504 29802 3516 29804
rect 3572 29802 3596 29804
rect 3652 29802 3676 29804
rect 3732 29802 3756 29804
rect 3812 29802 3824 29804
rect 3504 29750 3510 29802
rect 3572 29750 3574 29802
rect 3754 29750 3756 29802
rect 3818 29750 3824 29802
rect 3504 29748 3516 29750
rect 3572 29748 3596 29750
rect 3652 29748 3676 29750
rect 3732 29748 3756 29750
rect 3812 29748 3824 29750
rect 3504 29728 3824 29748
rect 2352 29700 2404 29706
rect 2352 29642 2404 29648
rect 3180 29700 3232 29706
rect 3180 29642 3232 29648
rect 3364 29700 3416 29706
rect 3364 29642 3416 29648
rect 1248 29564 1300 29570
rect 1248 29506 1300 29512
rect 2364 29502 2392 29642
rect 2352 29496 2404 29502
rect 2352 29438 2404 29444
rect 1156 29428 1208 29434
rect 1156 29370 1208 29376
rect 1168 28618 1196 29370
rect 2364 29162 2392 29438
rect 2996 29406 3048 29412
rect 2996 29348 3048 29354
rect 3272 29360 3324 29366
rect 2352 29156 2404 29162
rect 2352 29098 2404 29104
rect 3008 29026 3036 29348
rect 3272 29302 3324 29308
rect 2996 29020 3048 29026
rect 2996 28962 3048 28968
rect 1892 28816 1944 28822
rect 1614 28784 1670 28793
rect 1892 28758 1944 28764
rect 2076 28816 2128 28822
rect 2076 28758 2128 28764
rect 3180 28816 3232 28822
rect 3180 28758 3232 28764
rect 1614 28719 1670 28728
rect 1156 28612 1208 28618
rect 1156 28554 1208 28560
rect 1340 28272 1392 28278
rect 1340 28214 1392 28220
rect 1352 28006 1380 28214
rect 1340 28000 1392 28006
rect 1340 27942 1392 27948
rect 1432 27388 1484 27394
rect 1432 27330 1484 27336
rect 1156 27184 1208 27190
rect 1156 27126 1208 27132
rect 1444 27172 1472 27330
rect 1524 27184 1576 27190
rect 1444 27144 1524 27172
rect 696 26232 748 26238
rect 696 26174 748 26180
rect 708 25694 736 26174
rect 788 26096 840 26102
rect 788 26038 840 26044
rect 696 25688 748 25694
rect 696 25630 748 25636
rect 708 22974 736 25630
rect 800 25558 828 26038
rect 788 25552 840 25558
rect 788 25494 840 25500
rect 800 25286 828 25494
rect 788 25280 840 25286
rect 788 25222 840 25228
rect 1168 24742 1196 27126
rect 1444 26646 1472 27144
rect 1524 27126 1576 27132
rect 1432 26640 1484 26646
rect 1432 26582 1484 26588
rect 1444 26170 1472 26582
rect 1432 26164 1484 26170
rect 1432 26106 1484 26112
rect 1156 24736 1208 24742
rect 1156 24678 1208 24684
rect 972 24192 1024 24198
rect 972 24134 1024 24140
rect 984 23042 1012 24134
rect 1168 23586 1196 24678
rect 1156 23580 1208 23586
rect 1156 23522 1208 23528
rect 1340 23580 1392 23586
rect 1340 23522 1392 23528
rect 972 23036 1024 23042
rect 972 22978 1024 22984
rect 696 22968 748 22974
rect 696 22910 748 22916
rect 708 22294 736 22910
rect 984 22634 1012 22978
rect 972 22628 1024 22634
rect 972 22570 1024 22576
rect 1352 22294 1380 23522
rect 1432 23512 1484 23518
rect 1432 23454 1484 23460
rect 1444 22906 1472 23454
rect 1432 22900 1484 22906
rect 1432 22842 1484 22848
rect 1444 22634 1472 22842
rect 1432 22628 1484 22634
rect 1432 22570 1484 22576
rect 696 22288 748 22294
rect 696 22230 748 22236
rect 1340 22288 1392 22294
rect 1340 22230 1392 22236
rect 708 20798 736 22230
rect 1352 21410 1380 22230
rect 1340 21404 1392 21410
rect 1340 21346 1392 21352
rect 696 20792 748 20798
rect 696 20734 748 20740
rect 708 20186 736 20734
rect 788 20656 840 20662
rect 788 20598 840 20604
rect 1154 20624 1210 20633
rect 696 20180 748 20186
rect 696 20122 748 20128
rect 800 20118 828 20598
rect 1154 20559 1210 20568
rect 788 20112 840 20118
rect 788 20054 840 20060
rect 800 19846 828 20054
rect 1168 19914 1196 20559
rect 1352 20390 1380 21346
rect 1432 21336 1484 21342
rect 1432 21278 1484 21284
rect 1444 20730 1472 21278
rect 1432 20724 1484 20730
rect 1432 20666 1484 20672
rect 1444 20458 1472 20666
rect 1432 20452 1484 20458
rect 1432 20394 1484 20400
rect 1340 20384 1392 20390
rect 1340 20326 1392 20332
rect 1156 19908 1208 19914
rect 1156 19850 1208 19856
rect 788 19840 840 19846
rect 788 19782 840 19788
rect 1628 18486 1656 28719
rect 1904 28414 1932 28758
rect 2088 28414 2116 28758
rect 3192 28414 3220 28758
rect 1892 28408 1944 28414
rect 1892 28350 1944 28356
rect 2076 28408 2128 28414
rect 2260 28408 2312 28414
rect 2076 28350 2128 28356
rect 2180 28368 2260 28396
rect 1904 25898 1932 28350
rect 1984 27932 2036 27938
rect 1984 27874 2036 27880
rect 1996 27258 2024 27874
rect 2088 27394 2116 28350
rect 2180 27938 2208 28368
rect 2260 28350 2312 28356
rect 3180 28408 3232 28414
rect 3180 28350 3232 28356
rect 3088 28068 3140 28074
rect 3088 28010 3140 28016
rect 2168 27932 2220 27938
rect 2168 27874 2220 27880
rect 2180 27530 2208 27874
rect 2444 27864 2496 27870
rect 2444 27806 2496 27812
rect 2168 27524 2220 27530
rect 2168 27466 2220 27472
rect 2456 27462 2484 27806
rect 2444 27456 2496 27462
rect 2444 27398 2496 27404
rect 2076 27388 2128 27394
rect 2076 27330 2128 27336
rect 2720 27388 2772 27394
rect 2720 27330 2772 27336
rect 1984 27252 2036 27258
rect 1984 27194 2036 27200
rect 2732 26986 2760 27330
rect 3100 27326 3128 28010
rect 3284 27462 3312 29302
rect 3376 28074 3404 29642
rect 4100 29496 4152 29502
rect 4100 29438 4152 29444
rect 4112 29162 4140 29438
rect 4192 29360 4244 29366
rect 4192 29302 4244 29308
rect 4100 29156 4152 29162
rect 4100 29098 4152 29104
rect 4008 29020 4060 29026
rect 4008 28962 4060 28968
rect 3504 28716 3824 28736
rect 3504 28714 3516 28716
rect 3572 28714 3596 28716
rect 3652 28714 3676 28716
rect 3732 28714 3756 28716
rect 3812 28714 3824 28716
rect 3504 28662 3510 28714
rect 3572 28662 3574 28714
rect 3754 28662 3756 28714
rect 3818 28662 3824 28714
rect 3504 28660 3516 28662
rect 3572 28660 3596 28662
rect 3652 28660 3676 28662
rect 3732 28660 3756 28662
rect 3812 28660 3824 28662
rect 3504 28640 3824 28660
rect 3456 28272 3508 28278
rect 3456 28214 3508 28220
rect 3364 28068 3416 28074
rect 3364 28010 3416 28016
rect 3468 27938 3496 28214
rect 4020 27938 4048 28962
rect 4112 28006 4140 29098
rect 4204 28414 4232 29302
rect 4480 29162 4508 30118
rect 4652 30040 4704 30046
rect 4652 29982 4704 29988
rect 4664 29910 4692 29982
rect 4652 29904 4704 29910
rect 4652 29846 4704 29852
rect 4560 29564 4612 29570
rect 4560 29506 4612 29512
rect 4572 29366 4600 29506
rect 4664 29366 4692 29846
rect 5032 29706 5060 30458
rect 5400 30182 5428 30458
rect 5388 30176 5440 30182
rect 5388 30118 5440 30124
rect 5388 30040 5440 30046
rect 5388 29982 5440 29988
rect 5020 29700 5072 29706
rect 5020 29642 5072 29648
rect 5400 29638 5428 29982
rect 5492 29638 5520 30612
rect 6688 30250 6716 31664
rect 7516 31662 8188 31664
rect 6492 30244 6544 30250
rect 6492 30186 6544 30192
rect 6676 30244 6728 30250
rect 6676 30186 6728 30192
rect 6308 30108 6360 30114
rect 6308 30050 6360 30056
rect 5388 29632 5440 29638
rect 5388 29574 5440 29580
rect 5480 29632 5532 29638
rect 5480 29574 5532 29580
rect 6216 29496 6268 29502
rect 6216 29438 6268 29444
rect 5296 29428 5348 29434
rect 5296 29370 5348 29376
rect 4560 29360 4612 29366
rect 4560 29302 4612 29308
rect 4652 29360 4704 29366
rect 4652 29302 4704 29308
rect 5308 29162 5336 29370
rect 4468 29156 4520 29162
rect 4468 29098 4520 29104
rect 5296 29156 5348 29162
rect 5296 29098 5348 29104
rect 4284 29020 4336 29026
rect 4284 28962 4336 28968
rect 4296 28618 4324 28962
rect 4928 28952 4980 28958
rect 4928 28894 4980 28900
rect 4284 28612 4336 28618
rect 4284 28554 4336 28560
rect 4192 28408 4244 28414
rect 4192 28350 4244 28356
rect 4204 28278 4232 28350
rect 4192 28272 4244 28278
rect 4192 28214 4244 28220
rect 4100 28000 4152 28006
rect 4100 27942 4152 27948
rect 3364 27932 3416 27938
rect 3364 27874 3416 27880
rect 3456 27932 3508 27938
rect 3456 27874 3508 27880
rect 4008 27932 4060 27938
rect 4008 27874 4060 27880
rect 3272 27456 3324 27462
rect 3272 27398 3324 27404
rect 2904 27320 2956 27326
rect 2904 27262 2956 27268
rect 3088 27320 3140 27326
rect 3088 27262 3140 27268
rect 2720 26980 2772 26986
rect 2720 26922 2772 26928
rect 2720 26708 2772 26714
rect 2720 26650 2772 26656
rect 2732 26306 2760 26650
rect 2916 26442 2944 27262
rect 3376 27258 3404 27874
rect 3504 27628 3824 27648
rect 3504 27626 3516 27628
rect 3572 27626 3596 27628
rect 3652 27626 3676 27628
rect 3732 27626 3756 27628
rect 3812 27626 3824 27628
rect 3504 27574 3510 27626
rect 3572 27574 3574 27626
rect 3754 27574 3756 27626
rect 3818 27574 3824 27626
rect 3504 27572 3516 27574
rect 3572 27572 3596 27574
rect 3652 27572 3676 27574
rect 3732 27572 3756 27574
rect 3812 27572 3824 27574
rect 3504 27552 3824 27572
rect 3272 27252 3324 27258
rect 3272 27194 3324 27200
rect 3364 27252 3416 27258
rect 3364 27194 3416 27200
rect 3284 26850 3312 27194
rect 3272 26844 3324 26850
rect 3272 26786 3324 26792
rect 2904 26436 2956 26442
rect 2904 26378 2956 26384
rect 2720 26300 2772 26306
rect 2720 26242 2772 26248
rect 3284 26102 3312 26786
rect 3376 26646 3404 27194
rect 4020 27190 4048 27874
rect 4112 27530 4140 27942
rect 4100 27524 4152 27530
rect 4100 27466 4152 27472
rect 4008 27184 4060 27190
rect 4008 27126 4060 27132
rect 3364 26640 3416 26646
rect 3364 26582 3416 26588
rect 3272 26096 3324 26102
rect 3272 26038 3324 26044
rect 3376 26084 3404 26582
rect 3504 26540 3824 26560
rect 3504 26538 3516 26540
rect 3572 26538 3596 26540
rect 3652 26538 3676 26540
rect 3732 26538 3756 26540
rect 3812 26538 3824 26540
rect 3504 26486 3510 26538
rect 3572 26486 3574 26538
rect 3754 26486 3756 26538
rect 3818 26486 3824 26538
rect 3504 26484 3516 26486
rect 3572 26484 3596 26486
rect 3652 26484 3676 26486
rect 3732 26484 3756 26486
rect 3812 26484 3824 26486
rect 3504 26464 3824 26484
rect 3456 26096 3508 26102
rect 3376 26056 3456 26084
rect 1892 25892 1944 25898
rect 1892 25834 1944 25840
rect 2628 25892 2680 25898
rect 2628 25834 2680 25840
rect 2350 25248 2406 25257
rect 2350 25183 2406 25192
rect 2364 25150 2392 25183
rect 2640 25150 2668 25834
rect 3088 25824 3140 25830
rect 3088 25766 3140 25772
rect 2720 25688 2772 25694
rect 2720 25630 2772 25636
rect 2732 25150 2760 25630
rect 2352 25144 2404 25150
rect 2352 25086 2404 25092
rect 2628 25144 2680 25150
rect 2628 25086 2680 25092
rect 2720 25144 2772 25150
rect 2720 25086 2772 25092
rect 2364 24810 2392 25086
rect 1892 24804 1944 24810
rect 1892 24746 1944 24752
rect 2352 24804 2404 24810
rect 2352 24746 2404 24752
rect 1904 19370 1932 24746
rect 2640 24044 2668 25086
rect 3100 25014 3128 25766
rect 3284 25286 3312 26038
rect 3376 25762 3404 26056
rect 3456 26038 3508 26044
rect 3364 25756 3416 25762
rect 3364 25698 3416 25704
rect 3272 25280 3324 25286
rect 3272 25222 3324 25228
rect 3088 25008 3140 25014
rect 3088 24950 3140 24956
rect 3100 24470 3128 24950
rect 3376 24810 3404 25698
rect 3916 25688 3968 25694
rect 4204 25676 4232 28214
rect 4296 28074 4324 28554
rect 4744 28476 4796 28482
rect 4744 28418 4796 28424
rect 4836 28476 4888 28482
rect 4836 28418 4888 28424
rect 4284 28068 4336 28074
rect 4284 28010 4336 28016
rect 4560 26096 4612 26102
rect 4560 26038 4612 26044
rect 4284 25688 4336 25694
rect 4204 25648 4284 25676
rect 3916 25630 3968 25636
rect 4284 25630 4336 25636
rect 3504 25452 3824 25472
rect 3504 25450 3516 25452
rect 3572 25450 3596 25452
rect 3652 25450 3676 25452
rect 3732 25450 3756 25452
rect 3812 25450 3824 25452
rect 3504 25398 3510 25450
rect 3572 25398 3574 25450
rect 3754 25398 3756 25450
rect 3818 25398 3824 25450
rect 3504 25396 3516 25398
rect 3572 25396 3596 25398
rect 3652 25396 3676 25398
rect 3732 25396 3756 25398
rect 3812 25396 3824 25398
rect 3504 25376 3824 25396
rect 3824 25008 3876 25014
rect 3928 24996 3956 25630
rect 4296 25354 4324 25630
rect 4284 25348 4336 25354
rect 4284 25290 4336 25296
rect 4572 25150 4600 26038
rect 4560 25144 4612 25150
rect 4560 25086 4612 25092
rect 4284 25076 4336 25082
rect 4284 25018 4336 25024
rect 3876 24968 3956 24996
rect 3824 24950 3876 24956
rect 3364 24804 3416 24810
rect 3364 24746 3416 24752
rect 3928 24606 3956 24968
rect 4296 24606 4324 25018
rect 4572 25014 4600 25086
rect 4560 25008 4612 25014
rect 4560 24950 4612 24956
rect 4572 24606 4600 24950
rect 4652 24668 4704 24674
rect 4652 24610 4704 24616
rect 3916 24600 3968 24606
rect 3916 24542 3968 24548
rect 4284 24600 4336 24606
rect 4284 24542 4336 24548
rect 4560 24600 4612 24606
rect 4560 24542 4612 24548
rect 3088 24464 3140 24470
rect 3088 24406 3140 24412
rect 3100 24062 3128 24406
rect 3504 24364 3824 24384
rect 3504 24362 3516 24364
rect 3572 24362 3596 24364
rect 3652 24362 3676 24364
rect 3732 24362 3756 24364
rect 3812 24362 3824 24364
rect 3504 24310 3510 24362
rect 3572 24310 3574 24362
rect 3754 24310 3756 24362
rect 3818 24310 3824 24362
rect 3504 24308 3516 24310
rect 3572 24308 3596 24310
rect 3652 24308 3676 24310
rect 3732 24308 3756 24310
rect 3812 24308 3824 24310
rect 3504 24288 3824 24308
rect 3928 24266 3956 24542
rect 3916 24260 3968 24266
rect 3916 24202 3968 24208
rect 2720 24056 2772 24062
rect 2640 24016 2720 24044
rect 2640 23722 2668 24016
rect 2720 23998 2772 24004
rect 3088 24056 3140 24062
rect 3088 23998 3140 24004
rect 2628 23716 2680 23722
rect 2628 23658 2680 23664
rect 1984 23376 2036 23382
rect 1984 23318 2036 23324
rect 1996 23042 2024 23318
rect 1984 23036 2036 23042
rect 1984 22978 2036 22984
rect 2640 22634 2668 23658
rect 3100 23382 3128 23998
rect 3916 23988 3968 23994
rect 3916 23930 3968 23936
rect 3364 23580 3416 23586
rect 3364 23522 3416 23528
rect 3088 23376 3140 23382
rect 3088 23318 3140 23324
rect 3376 23042 3404 23522
rect 3504 23276 3824 23296
rect 3504 23274 3516 23276
rect 3572 23274 3596 23276
rect 3652 23274 3676 23276
rect 3732 23274 3756 23276
rect 3812 23274 3824 23276
rect 3504 23222 3510 23274
rect 3572 23222 3574 23274
rect 3754 23222 3756 23274
rect 3818 23222 3824 23274
rect 3504 23220 3516 23222
rect 3572 23220 3596 23222
rect 3652 23220 3676 23222
rect 3732 23220 3756 23222
rect 3812 23220 3824 23222
rect 3504 23200 3824 23220
rect 3364 23036 3416 23042
rect 3364 22978 3416 22984
rect 2904 22900 2956 22906
rect 2904 22842 2956 22848
rect 2628 22628 2680 22634
rect 2628 22570 2680 22576
rect 2640 20458 2668 22570
rect 2916 22090 2944 22842
rect 3272 22492 3324 22498
rect 3272 22434 3324 22440
rect 3180 22356 3232 22362
rect 3180 22298 3232 22304
rect 2904 22084 2956 22090
rect 2904 22026 2956 22032
rect 3192 21750 3220 22298
rect 3284 22090 3312 22434
rect 3928 22362 3956 23930
rect 4296 23926 4324 24542
rect 4572 24198 4600 24542
rect 4560 24192 4612 24198
rect 4560 24134 4612 24140
rect 4664 24130 4692 24610
rect 4652 24124 4704 24130
rect 4652 24066 4704 24072
rect 4756 24062 4784 28418
rect 4848 27870 4876 28418
rect 4940 28074 4968 28894
rect 5308 28890 5336 29098
rect 5664 29020 5716 29026
rect 5664 28962 5716 28968
rect 5572 28952 5624 28958
rect 5572 28894 5624 28900
rect 5296 28884 5348 28890
rect 5296 28826 5348 28832
rect 5020 28816 5072 28822
rect 5020 28758 5072 28764
rect 5032 28414 5060 28758
rect 5308 28618 5336 28826
rect 5296 28612 5348 28618
rect 5296 28554 5348 28560
rect 5584 28550 5612 28894
rect 5676 28618 5704 28962
rect 6228 28822 6256 29438
rect 6320 29366 6348 30050
rect 6308 29360 6360 29366
rect 6308 29302 6360 29308
rect 6216 28816 6268 28822
rect 6216 28758 6268 28764
rect 6228 28618 6256 28758
rect 5664 28612 5716 28618
rect 5664 28554 5716 28560
rect 6216 28612 6268 28618
rect 6216 28554 6268 28560
rect 5572 28544 5624 28550
rect 5572 28486 5624 28492
rect 5676 28414 5704 28554
rect 5020 28408 5072 28414
rect 5020 28350 5072 28356
rect 5664 28408 5716 28414
rect 5664 28350 5716 28356
rect 4928 28068 4980 28074
rect 4928 28010 4980 28016
rect 5676 27938 5704 28350
rect 5756 28272 5808 28278
rect 5756 28214 5808 28220
rect 5664 27932 5716 27938
rect 5664 27874 5716 27880
rect 4836 27864 4888 27870
rect 4836 27806 4888 27812
rect 5020 27864 5072 27870
rect 5020 27806 5072 27812
rect 4848 27530 4876 27806
rect 4836 27524 4888 27530
rect 4836 27466 4888 27472
rect 5032 27462 5060 27806
rect 5676 27462 5704 27874
rect 5768 27870 5796 28214
rect 5756 27864 5808 27870
rect 5756 27806 5808 27812
rect 5848 27864 5900 27870
rect 5848 27806 5900 27812
rect 5020 27456 5072 27462
rect 5020 27398 5072 27404
rect 5664 27456 5716 27462
rect 5664 27398 5716 27404
rect 5860 27394 5888 27806
rect 6032 27524 6084 27530
rect 6032 27466 6084 27472
rect 5848 27388 5900 27394
rect 5848 27330 5900 27336
rect 5756 25756 5808 25762
rect 5756 25698 5808 25704
rect 4928 25552 4980 25558
rect 4928 25494 4980 25500
rect 4940 25354 4968 25494
rect 4928 25348 4980 25354
rect 4928 25290 4980 25296
rect 5768 25286 5796 25698
rect 5756 25280 5808 25286
rect 5756 25222 5808 25228
rect 5860 25132 5888 27330
rect 6044 25830 6072 27466
rect 6124 26232 6176 26238
rect 6124 26174 6176 26180
rect 6032 25824 6084 25830
rect 6032 25766 6084 25772
rect 6044 25354 6072 25766
rect 6032 25348 6084 25354
rect 6032 25290 6084 25296
rect 5940 25144 5992 25150
rect 5860 25104 5940 25132
rect 5860 24674 5888 25104
rect 5940 25086 5992 25092
rect 5388 24668 5440 24674
rect 5388 24610 5440 24616
rect 5848 24668 5900 24674
rect 5848 24610 5900 24616
rect 4744 24056 4796 24062
rect 4744 23998 4796 24004
rect 4284 23920 4336 23926
rect 4284 23862 4336 23868
rect 4008 23376 4060 23382
rect 4008 23318 4060 23324
rect 4020 22838 4048 23318
rect 4008 22832 4060 22838
rect 4008 22774 4060 22780
rect 3916 22356 3968 22362
rect 3916 22298 3968 22304
rect 3504 22188 3824 22208
rect 3504 22186 3516 22188
rect 3572 22186 3596 22188
rect 3652 22186 3676 22188
rect 3732 22186 3756 22188
rect 3812 22186 3824 22188
rect 3504 22134 3510 22186
rect 3572 22134 3574 22186
rect 3754 22134 3756 22186
rect 3818 22134 3824 22186
rect 3504 22132 3516 22134
rect 3572 22132 3596 22134
rect 3652 22132 3676 22134
rect 3732 22132 3756 22134
rect 3812 22132 3824 22134
rect 3504 22112 3824 22132
rect 3272 22084 3324 22090
rect 3272 22026 3324 22032
rect 4020 21886 4048 22774
rect 4100 22492 4152 22498
rect 4100 22434 4152 22440
rect 4112 22090 4140 22434
rect 4192 22356 4244 22362
rect 4192 22298 4244 22304
rect 4204 22090 4232 22298
rect 4100 22084 4152 22090
rect 4100 22026 4152 22032
rect 4192 22084 4244 22090
rect 4192 22026 4244 22032
rect 4296 21954 4324 23862
rect 4560 23172 4612 23178
rect 4560 23114 4612 23120
rect 4376 22900 4428 22906
rect 4376 22842 4428 22848
rect 4284 21948 4336 21954
rect 4284 21890 4336 21896
rect 4008 21880 4060 21886
rect 4008 21822 4060 21828
rect 4100 21880 4152 21886
rect 4100 21822 4152 21828
rect 2720 21744 2772 21750
rect 2720 21686 2772 21692
rect 3180 21744 3232 21750
rect 3180 21686 3232 21692
rect 2732 21206 2760 21686
rect 3916 21404 3968 21410
rect 3916 21346 3968 21352
rect 3364 21336 3416 21342
rect 3364 21278 3416 21284
rect 2720 21200 2772 21206
rect 2720 21142 2772 21148
rect 2732 20866 2760 21142
rect 3376 21002 3404 21278
rect 3504 21100 3824 21120
rect 3504 21098 3516 21100
rect 3572 21098 3596 21100
rect 3652 21098 3676 21100
rect 3732 21098 3756 21100
rect 3812 21098 3824 21100
rect 3504 21046 3510 21098
rect 3572 21046 3574 21098
rect 3754 21046 3756 21098
rect 3818 21046 3824 21098
rect 3504 21044 3516 21046
rect 3572 21044 3596 21046
rect 3652 21044 3676 21046
rect 3732 21044 3756 21046
rect 3812 21044 3824 21046
rect 3504 21024 3824 21044
rect 3928 21002 3956 21346
rect 4008 21200 4060 21206
rect 4008 21142 4060 21148
rect 3364 20996 3416 21002
rect 3364 20938 3416 20944
rect 3916 20996 3968 21002
rect 3916 20938 3968 20944
rect 2720 20860 2772 20866
rect 2720 20802 2772 20808
rect 2628 20452 2680 20458
rect 2628 20394 2680 20400
rect 2640 19930 2668 20394
rect 2732 20322 2760 20802
rect 2720 20316 2772 20322
rect 2720 20258 2772 20264
rect 3180 20316 3232 20322
rect 3180 20258 3232 20264
rect 2640 19902 2760 19930
rect 3192 19914 3220 20258
rect 3272 20112 3324 20118
rect 3272 20054 3324 20060
rect 2732 19710 2760 19902
rect 3180 19908 3232 19914
rect 3180 19850 3232 19856
rect 2628 19704 2680 19710
rect 2628 19646 2680 19652
rect 2720 19704 2772 19710
rect 3284 19681 3312 20054
rect 3376 19710 3404 20938
rect 4020 20866 4048 21142
rect 4008 20860 4060 20866
rect 4008 20802 4060 20808
rect 4112 20798 4140 21822
rect 4296 21478 4324 21890
rect 4284 21472 4336 21478
rect 4284 21414 4336 21420
rect 4388 21410 4416 22842
rect 4572 22498 4600 23114
rect 4650 22800 4706 22809
rect 4650 22735 4706 22744
rect 4560 22492 4612 22498
rect 4560 22434 4612 22440
rect 4572 21546 4600 22434
rect 4560 21540 4612 21546
rect 4560 21482 4612 21488
rect 4376 21404 4428 21410
rect 4376 21346 4428 21352
rect 4560 21336 4612 21342
rect 4560 21278 4612 21284
rect 4192 21268 4244 21274
rect 4192 21210 4244 21216
rect 4204 20866 4232 21210
rect 4572 21206 4600 21278
rect 4560 21200 4612 21206
rect 4560 21142 4612 21148
rect 4376 20996 4428 21002
rect 4376 20938 4428 20944
rect 4192 20860 4244 20866
rect 4388 20848 4416 20938
rect 4468 20860 4520 20866
rect 4388 20820 4468 20848
rect 4192 20802 4244 20808
rect 4468 20802 4520 20808
rect 4100 20792 4152 20798
rect 4100 20734 4152 20740
rect 3504 20012 3824 20032
rect 3504 20010 3516 20012
rect 3572 20010 3596 20012
rect 3652 20010 3676 20012
rect 3732 20010 3756 20012
rect 3812 20010 3824 20012
rect 3504 19958 3510 20010
rect 3572 19958 3574 20010
rect 3754 19958 3756 20010
rect 3818 19958 3824 20010
rect 3504 19956 3516 19958
rect 3572 19956 3596 19958
rect 3652 19956 3676 19958
rect 3732 19956 3756 19958
rect 3812 19956 3824 19958
rect 3504 19936 3824 19956
rect 3364 19704 3416 19710
rect 2720 19646 2772 19652
rect 3270 19672 3326 19681
rect 2640 19370 2668 19646
rect 1892 19364 1944 19370
rect 1892 19306 1944 19312
rect 2628 19364 2680 19370
rect 2628 19306 2680 19312
rect 1616 18480 1668 18486
rect 1616 18422 1668 18428
rect 1616 17460 1668 17466
rect 1616 17402 1668 17408
rect 1248 17392 1300 17398
rect 1248 17334 1300 17340
rect 1260 17194 1288 17334
rect 1248 17188 1300 17194
rect 1248 17130 1300 17136
rect 1628 17058 1656 17402
rect 1800 17392 1852 17398
rect 1800 17334 1852 17340
rect 1616 17052 1668 17058
rect 1616 16994 1668 17000
rect 1154 16544 1210 16553
rect 1154 16479 1210 16488
rect 972 16304 1024 16310
rect 972 16246 1024 16252
rect 696 14264 748 14270
rect 696 14206 748 14212
rect 708 13590 736 14206
rect 984 14202 1012 16246
rect 1168 15970 1196 16479
rect 1628 16038 1656 16994
rect 1708 16984 1760 16990
rect 1708 16926 1760 16932
rect 1720 16378 1748 16926
rect 1812 16446 1840 17334
rect 1904 16446 1932 19306
rect 2732 19302 2760 19646
rect 3364 19646 3416 19652
rect 3270 19607 3272 19616
rect 3324 19607 3326 19616
rect 3272 19578 3324 19584
rect 3284 19547 3312 19578
rect 2720 19296 2772 19302
rect 2720 19238 2772 19244
rect 3272 19296 3324 19302
rect 3272 19238 3324 19244
rect 3284 18758 3312 19238
rect 3364 19228 3416 19234
rect 3364 19170 3416 19176
rect 3376 18826 3404 19170
rect 3504 18924 3824 18944
rect 3504 18922 3516 18924
rect 3572 18922 3596 18924
rect 3652 18922 3676 18924
rect 3732 18922 3756 18924
rect 3812 18922 3824 18924
rect 3504 18870 3510 18922
rect 3572 18870 3574 18922
rect 3754 18870 3756 18922
rect 3818 18870 3824 18922
rect 3504 18868 3516 18870
rect 3572 18868 3596 18870
rect 3652 18868 3676 18870
rect 3732 18868 3756 18870
rect 3812 18868 3824 18870
rect 3504 18848 3824 18868
rect 3364 18820 3416 18826
rect 3364 18762 3416 18768
rect 3272 18752 3324 18758
rect 3272 18694 3324 18700
rect 4008 18276 4060 18282
rect 4008 18218 4060 18224
rect 3504 17836 3824 17856
rect 3504 17834 3516 17836
rect 3572 17834 3596 17836
rect 3652 17834 3676 17836
rect 3732 17834 3756 17836
rect 3812 17834 3824 17836
rect 3504 17782 3510 17834
rect 3572 17782 3574 17834
rect 3754 17782 3756 17834
rect 3818 17782 3824 17834
rect 3504 17780 3516 17782
rect 3572 17780 3596 17782
rect 3652 17780 3676 17782
rect 3732 17780 3756 17782
rect 3812 17780 3824 17782
rect 3504 17760 3824 17780
rect 2352 17528 2404 17534
rect 2352 17470 2404 17476
rect 2364 17398 2392 17470
rect 2352 17392 2404 17398
rect 2352 17334 2404 17340
rect 3916 17392 3968 17398
rect 3916 17334 3968 17340
rect 2364 17058 2392 17334
rect 2352 17052 2404 17058
rect 2352 16994 2404 17000
rect 3928 16990 3956 17334
rect 3916 16984 3968 16990
rect 3916 16926 3968 16932
rect 2536 16848 2588 16854
rect 2536 16790 2588 16796
rect 2548 16446 2576 16790
rect 3504 16748 3824 16768
rect 3504 16746 3516 16748
rect 3572 16746 3596 16748
rect 3652 16746 3676 16748
rect 3732 16746 3756 16748
rect 3812 16746 3824 16748
rect 3504 16694 3510 16746
rect 3572 16694 3574 16746
rect 3754 16694 3756 16746
rect 3818 16694 3824 16746
rect 3504 16692 3516 16694
rect 3572 16692 3596 16694
rect 3652 16692 3676 16694
rect 3732 16692 3756 16694
rect 3812 16692 3824 16694
rect 3504 16672 3824 16692
rect 3928 16650 3956 16926
rect 3916 16644 3968 16650
rect 3916 16586 3968 16592
rect 1800 16440 1852 16446
rect 1800 16382 1852 16388
rect 1892 16440 1944 16446
rect 1892 16382 1944 16388
rect 2536 16440 2588 16446
rect 2536 16382 2588 16388
rect 3272 16440 3324 16446
rect 3272 16382 3324 16388
rect 1708 16372 1760 16378
rect 1708 16314 1760 16320
rect 1720 16106 1748 16314
rect 1708 16100 1760 16106
rect 1708 16042 1760 16048
rect 1616 16032 1668 16038
rect 1616 15974 1668 15980
rect 3284 15970 3312 16382
rect 3364 16372 3416 16378
rect 3364 16314 3416 16320
rect 1156 15964 1208 15970
rect 1156 15906 1208 15912
rect 1984 15964 2036 15970
rect 1984 15906 2036 15912
rect 3272 15964 3324 15970
rect 3272 15906 3324 15912
rect 1168 15562 1196 15906
rect 1996 15562 2024 15906
rect 2260 15896 2312 15902
rect 2260 15838 2312 15844
rect 1156 15556 1208 15562
rect 1156 15498 1208 15504
rect 1984 15556 2036 15562
rect 1984 15498 2036 15504
rect 1996 15018 2024 15498
rect 2272 15358 2300 15838
rect 2260 15352 2312 15358
rect 2260 15294 2312 15300
rect 3284 15290 3312 15906
rect 3376 15766 3404 16314
rect 4020 15970 4048 18218
rect 4376 18208 4428 18214
rect 4376 18150 4428 18156
rect 4284 17052 4336 17058
rect 4284 16994 4336 17000
rect 4100 16984 4152 16990
rect 4100 16926 4152 16932
rect 4112 16650 4140 16926
rect 4296 16650 4324 16994
rect 4388 16990 4416 18150
rect 4468 17460 4520 17466
rect 4468 17402 4520 17408
rect 4560 17460 4612 17466
rect 4560 17402 4612 17408
rect 4480 17058 4508 17402
rect 4572 17369 4600 17402
rect 4558 17360 4614 17369
rect 4558 17295 4614 17304
rect 4468 17052 4520 17058
rect 4468 16994 4520 17000
rect 4376 16984 4428 16990
rect 4376 16926 4428 16932
rect 4468 16916 4520 16922
rect 4468 16858 4520 16864
rect 4480 16650 4508 16858
rect 4100 16644 4152 16650
rect 4100 16586 4152 16592
rect 4284 16644 4336 16650
rect 4284 16586 4336 16592
rect 4468 16644 4520 16650
rect 4468 16586 4520 16592
rect 4008 15964 4060 15970
rect 4008 15906 4060 15912
rect 3364 15760 3416 15766
rect 3364 15702 3416 15708
rect 3272 15284 3324 15290
rect 3272 15226 3324 15232
rect 3376 15018 3404 15702
rect 3504 15660 3824 15680
rect 3504 15658 3516 15660
rect 3572 15658 3596 15660
rect 3652 15658 3676 15660
rect 3732 15658 3756 15660
rect 3812 15658 3824 15660
rect 3504 15606 3510 15658
rect 3572 15606 3574 15658
rect 3754 15606 3756 15658
rect 3818 15606 3824 15658
rect 3504 15604 3516 15606
rect 3572 15604 3596 15606
rect 3652 15604 3676 15606
rect 3732 15604 3756 15606
rect 3812 15604 3824 15606
rect 3504 15584 3824 15604
rect 4020 15494 4048 15906
rect 4112 15494 4140 16586
rect 4296 16446 4324 16586
rect 4376 16508 4428 16514
rect 4376 16450 4428 16456
rect 4284 16440 4336 16446
rect 4284 16382 4336 16388
rect 4008 15488 4060 15494
rect 3928 15448 4008 15476
rect 1984 15012 2036 15018
rect 1984 14954 2036 14960
rect 3364 15012 3416 15018
rect 3364 14954 3416 14960
rect 1432 14672 1484 14678
rect 1432 14614 1484 14620
rect 972 14196 1024 14202
rect 1444 14184 1472 14614
rect 1996 14338 2024 14954
rect 2626 14640 2682 14649
rect 2626 14575 2682 14584
rect 1984 14332 2036 14338
rect 1984 14274 2036 14280
rect 1708 14196 1760 14202
rect 1444 14156 1708 14184
rect 972 14138 1024 14144
rect 1708 14138 1760 14144
rect 984 13930 1012 14138
rect 972 13924 1024 13930
rect 972 13866 1024 13872
rect 696 13584 748 13590
rect 696 13526 748 13532
rect 972 13584 1024 13590
rect 972 13526 1024 13532
rect 984 12745 1012 13526
rect 970 12736 1026 12745
rect 970 12671 1026 12680
rect 1156 12700 1208 12706
rect 1156 12642 1208 12648
rect 1168 11958 1196 12642
rect 1720 12638 1748 14138
rect 2640 13930 2668 14575
rect 3504 14572 3824 14592
rect 3504 14570 3516 14572
rect 3572 14570 3596 14572
rect 3652 14570 3676 14572
rect 3732 14570 3756 14572
rect 3812 14570 3824 14572
rect 3504 14518 3510 14570
rect 3572 14518 3574 14570
rect 3754 14518 3756 14570
rect 3818 14518 3824 14570
rect 3504 14516 3516 14518
rect 3572 14516 3596 14518
rect 3652 14516 3676 14518
rect 3732 14516 3756 14518
rect 3812 14516 3824 14518
rect 3504 14496 3824 14516
rect 3928 14134 3956 15448
rect 4008 15430 4060 15436
rect 4100 15488 4152 15494
rect 4100 15430 4152 15436
rect 4296 15426 4324 16382
rect 4284 15420 4336 15426
rect 4284 15362 4336 15368
rect 4008 14808 4060 14814
rect 4008 14750 4060 14756
rect 4100 14808 4152 14814
rect 4100 14750 4152 14756
rect 4020 14474 4048 14750
rect 4008 14468 4060 14474
rect 4008 14410 4060 14416
rect 3916 14128 3968 14134
rect 3916 14070 3968 14076
rect 2628 13924 2680 13930
rect 2628 13866 2680 13872
rect 4020 13726 4048 14410
rect 4112 14338 4140 14750
rect 4100 14332 4152 14338
rect 4100 14274 4152 14280
rect 4388 14214 4416 16450
rect 4468 15556 4520 15562
rect 4468 15498 4520 15504
rect 4480 14882 4508 15498
rect 4468 14876 4520 14882
rect 4468 14818 4520 14824
rect 4560 14876 4612 14882
rect 4560 14818 4612 14824
rect 4572 14270 4600 14818
rect 4560 14264 4612 14270
rect 4388 14186 4508 14214
rect 4560 14206 4612 14212
rect 4664 14214 4692 22735
rect 4928 22492 4980 22498
rect 4928 22434 4980 22440
rect 4940 22022 4968 22434
rect 4744 22016 4796 22022
rect 4744 21958 4796 21964
rect 4928 22016 4980 22022
rect 4928 21958 4980 21964
rect 4756 21886 4784 21958
rect 4744 21880 4796 21886
rect 4744 21822 4796 21828
rect 4836 21744 4888 21750
rect 4836 21686 4888 21692
rect 4744 21404 4796 21410
rect 4744 21346 4796 21352
rect 4756 20866 4784 21346
rect 4744 20860 4796 20866
rect 4744 20802 4796 20808
rect 4848 20118 4876 21686
rect 4928 20996 4980 21002
rect 4928 20938 4980 20944
rect 4940 20798 4968 20938
rect 4928 20792 4980 20798
rect 4928 20734 4980 20740
rect 4836 20112 4888 20118
rect 4836 20054 4888 20060
rect 4940 19681 4968 20734
rect 4926 19672 4982 19681
rect 4926 19607 4982 19616
rect 5400 19302 5428 24610
rect 5756 24056 5808 24062
rect 5756 23998 5808 24004
rect 5768 23178 5796 23998
rect 6044 23874 6072 25290
rect 5952 23846 6072 23874
rect 5756 23172 5808 23178
rect 5756 23114 5808 23120
rect 5952 22430 5980 23846
rect 6136 22498 6164 26174
rect 6216 24600 6268 24606
rect 6216 24542 6268 24548
rect 6124 22492 6176 22498
rect 6124 22434 6176 22440
rect 5940 22424 5992 22430
rect 5940 22366 5992 22372
rect 5572 22356 5624 22362
rect 5572 22298 5624 22304
rect 5584 21342 5612 22298
rect 5952 22090 5980 22366
rect 5940 22084 5992 22090
rect 5940 22026 5992 22032
rect 6124 21880 6176 21886
rect 6124 21822 6176 21828
rect 5848 21404 5900 21410
rect 5848 21346 5900 21352
rect 5572 21336 5624 21342
rect 5572 21278 5624 21284
rect 5756 21336 5808 21342
rect 5756 21278 5808 21284
rect 5768 20458 5796 21278
rect 5860 21002 5888 21346
rect 5848 20996 5900 21002
rect 5848 20938 5900 20944
rect 6136 20769 6164 21822
rect 6228 20798 6256 24542
rect 6320 24062 6348 29302
rect 6504 25626 6532 30186
rect 6860 30040 6912 30046
rect 6860 29982 6912 29988
rect 6872 29026 6900 29982
rect 7320 29496 7372 29502
rect 7320 29438 7372 29444
rect 6860 29020 6912 29026
rect 6860 28962 6912 28968
rect 6872 28618 6900 28962
rect 7332 28890 7360 29438
rect 7320 28884 7372 28890
rect 7320 28826 7372 28832
rect 6952 28816 7004 28822
rect 6952 28758 7004 28764
rect 6860 28612 6912 28618
rect 6860 28554 6912 28560
rect 6872 27462 6900 28554
rect 6964 28414 6992 28758
rect 6952 28408 7004 28414
rect 6952 28350 7004 28356
rect 6860 27456 6912 27462
rect 6860 27398 6912 27404
rect 6584 26844 6636 26850
rect 6584 26786 6636 26792
rect 6596 25830 6624 26786
rect 6872 26714 6900 27398
rect 6952 27184 7004 27190
rect 6952 27126 7004 27132
rect 6964 26782 6992 27126
rect 6952 26776 7004 26782
rect 6952 26718 7004 26724
rect 6860 26708 6912 26714
rect 6860 26650 6912 26656
rect 6768 26640 6820 26646
rect 6768 26582 6820 26588
rect 6780 26442 6808 26582
rect 6768 26436 6820 26442
rect 6768 26378 6820 26384
rect 6872 26306 6900 26650
rect 6964 26374 6992 26718
rect 7228 26640 7280 26646
rect 7228 26582 7280 26588
rect 6952 26368 7004 26374
rect 6952 26310 7004 26316
rect 6860 26300 6912 26306
rect 6860 26242 6912 26248
rect 6584 25824 6636 25830
rect 6584 25766 6636 25772
rect 7240 25694 7268 26582
rect 7228 25688 7280 25694
rect 7228 25630 7280 25636
rect 6492 25620 6544 25626
rect 6492 25562 6544 25568
rect 6400 25076 6452 25082
rect 6400 25018 6452 25024
rect 6308 24056 6360 24062
rect 6308 23998 6360 24004
rect 6308 23036 6360 23042
rect 6308 22978 6360 22984
rect 6320 22634 6348 22978
rect 6308 22628 6360 22634
rect 6308 22570 6360 22576
rect 6308 22288 6360 22294
rect 6308 22230 6360 22236
rect 6320 21342 6348 22230
rect 6412 21886 6440 25018
rect 7044 25008 7096 25014
rect 7044 24950 7096 24956
rect 6952 24056 7004 24062
rect 6952 23998 7004 24004
rect 6584 23988 6636 23994
rect 6584 23930 6636 23936
rect 6596 23110 6624 23930
rect 6584 23104 6636 23110
rect 6584 23046 6636 23052
rect 6492 22968 6544 22974
rect 6492 22910 6544 22916
rect 6504 22634 6532 22910
rect 6492 22628 6544 22634
rect 6492 22570 6544 22576
rect 6504 22022 6532 22570
rect 6964 22566 6992 23998
rect 7056 23518 7084 24950
rect 7136 23580 7188 23586
rect 7136 23522 7188 23528
rect 7044 23512 7096 23518
rect 7044 23454 7096 23460
rect 6952 22560 7004 22566
rect 6872 22520 6952 22548
rect 6492 22016 6544 22022
rect 6492 21958 6544 21964
rect 6400 21880 6452 21886
rect 6400 21822 6452 21828
rect 6412 21342 6440 21822
rect 6308 21336 6360 21342
rect 6308 21278 6360 21284
rect 6400 21336 6452 21342
rect 6400 21278 6452 21284
rect 6320 20934 6348 21278
rect 6308 20928 6360 20934
rect 6308 20870 6360 20876
rect 6216 20792 6268 20798
rect 6122 20760 6178 20769
rect 6216 20734 6268 20740
rect 6122 20695 6178 20704
rect 5756 20452 5808 20458
rect 5756 20394 5808 20400
rect 5388 19296 5440 19302
rect 5388 19238 5440 19244
rect 4836 19228 4888 19234
rect 4836 19170 4888 19176
rect 4848 18486 4876 19170
rect 5296 19160 5348 19166
rect 5296 19102 5348 19108
rect 5308 18826 5336 19102
rect 5296 18820 5348 18826
rect 5296 18762 5348 18768
rect 5110 18720 5166 18729
rect 5110 18655 5166 18664
rect 4836 18480 4888 18486
rect 4836 18422 4888 18428
rect 4744 18140 4796 18146
rect 4744 18082 4796 18088
rect 4756 17670 4784 18082
rect 4744 17664 4796 17670
rect 4744 17606 4796 17612
rect 4756 17194 4784 17606
rect 4848 17466 4876 18422
rect 4836 17460 4888 17466
rect 4836 17402 4888 17408
rect 4744 17188 4796 17194
rect 4744 17130 4796 17136
rect 4744 15760 4796 15766
rect 4744 15702 4796 15708
rect 4756 15562 4784 15702
rect 4744 15556 4796 15562
rect 4744 15498 4796 15504
rect 4756 14882 4784 15498
rect 4848 15494 4876 17402
rect 4836 15488 4888 15494
rect 4836 15430 4888 15436
rect 4848 14882 4876 15430
rect 4744 14876 4796 14882
rect 4744 14818 4796 14824
rect 4836 14876 4888 14882
rect 4836 14818 4888 14824
rect 4756 14474 4784 14818
rect 4744 14468 4796 14474
rect 4744 14410 4796 14416
rect 4848 14338 4876 14818
rect 4836 14332 4888 14338
rect 4836 14274 4888 14280
rect 4664 14186 4784 14214
rect 4284 14128 4336 14134
rect 4284 14070 4336 14076
rect 4100 13856 4152 13862
rect 4100 13798 4152 13804
rect 3364 13720 3416 13726
rect 3364 13662 3416 13668
rect 4008 13720 4060 13726
rect 4008 13662 4060 13668
rect 3376 13318 3404 13662
rect 3504 13484 3824 13504
rect 3504 13482 3516 13484
rect 3572 13482 3596 13484
rect 3652 13482 3676 13484
rect 3732 13482 3756 13484
rect 3812 13482 3824 13484
rect 3504 13430 3510 13482
rect 3572 13430 3574 13482
rect 3754 13430 3756 13482
rect 3818 13430 3824 13482
rect 3504 13428 3516 13430
rect 3572 13428 3596 13430
rect 3652 13428 3676 13430
rect 3732 13428 3756 13430
rect 3812 13428 3824 13430
rect 3504 13408 3824 13428
rect 4020 13386 4048 13662
rect 4008 13380 4060 13386
rect 4008 13322 4060 13328
rect 3364 13312 3416 13318
rect 3364 13254 3416 13260
rect 3916 13312 3968 13318
rect 3916 13254 3968 13260
rect 3928 13182 3956 13254
rect 3916 13176 3968 13182
rect 3916 13118 3968 13124
rect 4112 13114 4140 13798
rect 4100 13108 4152 13114
rect 4100 13050 4152 13056
rect 2074 12736 2130 12745
rect 2074 12671 2130 12680
rect 1708 12632 1760 12638
rect 1708 12574 1760 12580
rect 1246 12464 1302 12473
rect 1246 12399 1302 12408
rect 1260 12162 1288 12399
rect 1720 12298 1748 12574
rect 1708 12292 1760 12298
rect 1708 12234 1760 12240
rect 1248 12156 1300 12162
rect 1248 12098 1300 12104
rect 1156 11952 1208 11958
rect 1156 11894 1208 11900
rect 1338 11648 1394 11657
rect 1338 11583 1340 11592
rect 1392 11583 1394 11592
rect 1340 11554 1392 11560
rect 1352 11210 1380 11554
rect 1432 11408 1484 11414
rect 1432 11350 1484 11356
rect 1340 11204 1392 11210
rect 1340 11146 1392 11152
rect 1444 10870 1472 11350
rect 1432 10864 1484 10870
rect 1432 10806 1484 10812
rect 1444 10569 1472 10806
rect 1430 10560 1486 10569
rect 1430 10495 1486 10504
rect 1984 10456 2036 10462
rect 1984 10398 2036 10404
rect 1996 10122 2024 10398
rect 1984 10116 2036 10122
rect 1984 10058 2036 10064
rect 2088 9986 2116 12671
rect 3272 12632 3324 12638
rect 3272 12574 3324 12580
rect 3284 12094 3312 12574
rect 3504 12396 3824 12416
rect 3504 12394 3516 12396
rect 3572 12394 3596 12396
rect 3652 12394 3676 12396
rect 3732 12394 3756 12396
rect 3812 12394 3824 12396
rect 3504 12342 3510 12394
rect 3572 12342 3574 12394
rect 3754 12342 3756 12394
rect 3818 12342 3824 12394
rect 3504 12340 3516 12342
rect 3572 12340 3596 12342
rect 3652 12340 3676 12342
rect 3732 12340 3756 12342
rect 3812 12340 3824 12342
rect 3504 12320 3824 12340
rect 4112 12298 4140 13050
rect 4100 12292 4152 12298
rect 4100 12234 4152 12240
rect 3272 12088 3324 12094
rect 3272 12030 3324 12036
rect 2444 11952 2496 11958
rect 2444 11894 2496 11900
rect 2456 11006 2484 11894
rect 3504 11308 3824 11328
rect 3504 11306 3516 11308
rect 3572 11306 3596 11308
rect 3652 11306 3676 11308
rect 3732 11306 3756 11308
rect 3812 11306 3824 11308
rect 3504 11254 3510 11306
rect 3572 11254 3574 11306
rect 3754 11254 3756 11306
rect 3818 11254 3824 11306
rect 3504 11252 3516 11254
rect 3572 11252 3596 11254
rect 3652 11252 3676 11254
rect 3732 11252 3756 11254
rect 3812 11252 3824 11254
rect 3504 11232 3824 11252
rect 2444 11000 2496 11006
rect 2444 10942 2496 10948
rect 2076 9980 2128 9986
rect 2076 9922 2128 9928
rect 2088 9578 2116 9922
rect 2352 9844 2404 9850
rect 2352 9786 2404 9792
rect 2076 9572 2128 9578
rect 2076 9514 2128 9520
rect 1156 9436 1208 9442
rect 1156 9378 1208 9384
rect 696 8892 748 8898
rect 696 8834 748 8840
rect 708 8490 736 8834
rect 972 8756 1024 8762
rect 972 8698 1024 8704
rect 696 8484 748 8490
rect 696 8426 748 8432
rect 708 6246 736 8426
rect 984 8218 1012 8698
rect 972 8212 1024 8218
rect 972 8154 1024 8160
rect 1168 7742 1196 9378
rect 1432 9368 1484 9374
rect 1432 9310 1484 9316
rect 1444 8762 1472 9310
rect 1616 9232 1668 9238
rect 1616 9174 1668 9180
rect 1628 8898 1656 9174
rect 2088 9034 2116 9514
rect 2364 9510 2392 9786
rect 2352 9504 2404 9510
rect 2352 9446 2404 9452
rect 2456 9442 2484 10942
rect 2996 10864 3048 10870
rect 2996 10806 3048 10812
rect 3008 10530 3036 10806
rect 2996 10524 3048 10530
rect 2996 10466 3048 10472
rect 3008 9850 3036 10466
rect 4100 10456 4152 10462
rect 4100 10398 4152 10404
rect 3916 10320 3968 10326
rect 3916 10262 3968 10268
rect 3504 10220 3824 10240
rect 3504 10218 3516 10220
rect 3572 10218 3596 10220
rect 3652 10218 3676 10220
rect 3732 10218 3756 10220
rect 3812 10218 3824 10220
rect 3504 10166 3510 10218
rect 3572 10166 3574 10218
rect 3754 10166 3756 10218
rect 3818 10166 3824 10218
rect 3504 10164 3516 10166
rect 3572 10164 3596 10166
rect 3652 10164 3676 10166
rect 3732 10164 3756 10166
rect 3812 10164 3824 10166
rect 3504 10144 3824 10164
rect 2996 9844 3048 9850
rect 2996 9786 3048 9792
rect 3180 9504 3232 9510
rect 3180 9446 3232 9452
rect 2444 9436 2496 9442
rect 2444 9378 2496 9384
rect 3192 9034 3220 9446
rect 3928 9442 3956 10262
rect 4112 9986 4140 10398
rect 4100 9980 4152 9986
rect 4100 9922 4152 9928
rect 4112 9510 4140 9922
rect 4100 9504 4152 9510
rect 4100 9446 4152 9452
rect 3916 9436 3968 9442
rect 3916 9378 3968 9384
rect 4008 9436 4060 9442
rect 4008 9378 4060 9384
rect 4192 9436 4244 9442
rect 4192 9378 4244 9384
rect 3504 9132 3824 9152
rect 3504 9130 3516 9132
rect 3572 9130 3596 9132
rect 3652 9130 3676 9132
rect 3732 9130 3756 9132
rect 3812 9130 3824 9132
rect 3504 9078 3510 9130
rect 3572 9078 3574 9130
rect 3754 9078 3756 9130
rect 3818 9078 3824 9130
rect 3504 9076 3516 9078
rect 3572 9076 3596 9078
rect 3652 9076 3676 9078
rect 3732 9076 3756 9078
rect 3812 9076 3824 9078
rect 3504 9056 3824 9076
rect 2076 9028 2128 9034
rect 2076 8970 2128 8976
rect 3180 9028 3232 9034
rect 3180 8970 3232 8976
rect 1616 8892 1668 8898
rect 1616 8834 1668 8840
rect 3640 8824 3692 8830
rect 3640 8766 3692 8772
rect 1432 8756 1484 8762
rect 1432 8698 1484 8704
rect 2904 8756 2956 8762
rect 2904 8698 2956 8704
rect 1444 8490 1472 8698
rect 1432 8484 1484 8490
rect 1432 8426 1484 8432
rect 2916 8422 2944 8698
rect 2904 8416 2956 8422
rect 2904 8358 2956 8364
rect 2352 8348 2404 8354
rect 2352 8290 2404 8296
rect 1800 8280 1852 8286
rect 1800 8222 1852 8228
rect 1708 8212 1760 8218
rect 1708 8154 1760 8160
rect 1720 7946 1748 8154
rect 1708 7940 1760 7946
rect 1708 7882 1760 7888
rect 1156 7736 1208 7742
rect 1156 7678 1208 7684
rect 1432 7668 1484 7674
rect 1432 7610 1484 7616
rect 878 6480 934 6489
rect 878 6415 934 6424
rect 892 6314 920 6415
rect 880 6308 932 6314
rect 880 6250 932 6256
rect 696 6240 748 6246
rect 696 6182 748 6188
rect 708 5634 736 6182
rect 696 5628 748 5634
rect 696 5570 748 5576
rect 892 5226 920 6250
rect 1444 5498 1472 7610
rect 1812 7606 1840 8222
rect 2364 7810 2392 8290
rect 2916 7946 2944 8358
rect 3652 8354 3680 8766
rect 3928 8490 3956 9378
rect 4020 8694 4048 9378
rect 4204 8898 4232 9378
rect 4192 8892 4244 8898
rect 4192 8834 4244 8840
rect 4008 8688 4060 8694
rect 4008 8630 4060 8636
rect 3916 8484 3968 8490
rect 3916 8426 3968 8432
rect 4020 8422 4048 8630
rect 4204 8422 4232 8834
rect 4008 8416 4060 8422
rect 4008 8358 4060 8364
rect 4192 8416 4244 8422
rect 4192 8358 4244 8364
rect 3364 8348 3416 8354
rect 3364 8290 3416 8296
rect 3640 8348 3692 8354
rect 3640 8290 3692 8296
rect 3376 7946 3404 8290
rect 3504 8044 3824 8064
rect 3504 8042 3516 8044
rect 3572 8042 3596 8044
rect 3652 8042 3676 8044
rect 3732 8042 3756 8044
rect 3812 8042 3824 8044
rect 3504 7990 3510 8042
rect 3572 7990 3574 8042
rect 3754 7990 3756 8042
rect 3818 7990 3824 8042
rect 3504 7988 3516 7990
rect 3572 7988 3596 7990
rect 3652 7988 3676 7990
rect 3732 7988 3756 7990
rect 3812 7988 3824 7990
rect 3504 7968 3824 7988
rect 4020 7946 4048 8358
rect 2904 7940 2956 7946
rect 2904 7882 2956 7888
rect 3364 7940 3416 7946
rect 3364 7882 3416 7888
rect 4008 7940 4060 7946
rect 4008 7882 4060 7888
rect 2352 7804 2404 7810
rect 2352 7746 2404 7752
rect 1800 7600 1852 7606
rect 1800 7542 1852 7548
rect 1812 6110 1840 7542
rect 3376 7266 3404 7882
rect 3364 7260 3416 7266
rect 3364 7202 3416 7208
rect 3376 6858 3404 7202
rect 3916 7192 3968 7198
rect 3916 7134 3968 7140
rect 3504 6956 3824 6976
rect 3504 6954 3516 6956
rect 3572 6954 3596 6956
rect 3652 6954 3676 6956
rect 3732 6954 3756 6956
rect 3812 6954 3824 6956
rect 3504 6902 3510 6954
rect 3572 6902 3574 6954
rect 3754 6902 3756 6954
rect 3818 6902 3824 6954
rect 3504 6900 3516 6902
rect 3572 6900 3596 6902
rect 3652 6900 3676 6902
rect 3732 6900 3756 6902
rect 3812 6900 3824 6902
rect 3504 6880 3824 6900
rect 3364 6852 3416 6858
rect 3364 6794 3416 6800
rect 3928 6518 3956 7134
rect 4020 6858 4048 7882
rect 4008 6852 4060 6858
rect 4008 6794 4060 6800
rect 4296 6625 4324 14070
rect 4480 10530 4508 14186
rect 4652 12700 4704 12706
rect 4652 12642 4704 12648
rect 4664 12298 4692 12642
rect 4652 12292 4704 12298
rect 4652 12234 4704 12240
rect 4468 10524 4520 10530
rect 4468 10466 4520 10472
rect 4480 10122 4508 10466
rect 4560 10320 4612 10326
rect 4560 10262 4612 10268
rect 4572 10122 4600 10262
rect 4468 10116 4520 10122
rect 4468 10058 4520 10064
rect 4560 10116 4612 10122
rect 4560 10058 4612 10064
rect 4480 9034 4508 10058
rect 4468 9028 4520 9034
rect 4468 8970 4520 8976
rect 4480 8830 4508 8970
rect 4756 8898 4784 14186
rect 4836 12632 4888 12638
rect 4836 12574 4888 12580
rect 4848 11958 4876 12574
rect 5124 12162 5152 18655
rect 5400 18010 5428 19238
rect 5480 18684 5532 18690
rect 5480 18626 5532 18632
rect 5492 18078 5520 18626
rect 5940 18548 5992 18554
rect 5940 18490 5992 18496
rect 5480 18072 5532 18078
rect 5480 18014 5532 18020
rect 5388 18004 5440 18010
rect 5388 17946 5440 17952
rect 5296 17936 5348 17942
rect 5296 17878 5348 17884
rect 5308 17738 5336 17878
rect 5296 17732 5348 17738
rect 5296 17674 5348 17680
rect 5204 17392 5256 17398
rect 5204 17334 5256 17340
rect 5216 17058 5244 17334
rect 5400 17058 5428 17946
rect 5492 17534 5520 18014
rect 5480 17528 5532 17534
rect 5480 17470 5532 17476
rect 5492 17058 5520 17470
rect 5204 17052 5256 17058
rect 5204 16994 5256 17000
rect 5388 17052 5440 17058
rect 5388 16994 5440 17000
rect 5480 17052 5532 17058
rect 5480 16994 5532 17000
rect 5216 16650 5244 16994
rect 5400 16650 5428 16994
rect 5204 16644 5256 16650
rect 5204 16586 5256 16592
rect 5388 16644 5440 16650
rect 5388 16586 5440 16592
rect 5492 16582 5520 16994
rect 5756 16984 5808 16990
rect 5756 16926 5808 16932
rect 5768 16650 5796 16926
rect 5756 16644 5808 16650
rect 5756 16586 5808 16592
rect 5480 16576 5532 16582
rect 5480 16518 5532 16524
rect 5756 15964 5808 15970
rect 5756 15906 5808 15912
rect 5388 15760 5440 15766
rect 5388 15702 5440 15708
rect 5296 15216 5348 15222
rect 5296 15158 5348 15164
rect 5308 14134 5336 15158
rect 5400 15018 5428 15702
rect 5768 15562 5796 15906
rect 5848 15896 5900 15902
rect 5848 15838 5900 15844
rect 5756 15556 5808 15562
rect 5756 15498 5808 15504
rect 5860 15494 5888 15838
rect 5848 15488 5900 15494
rect 5848 15430 5900 15436
rect 5388 15012 5440 15018
rect 5440 14972 5520 15000
rect 5388 14954 5440 14960
rect 5388 14808 5440 14814
rect 5388 14750 5440 14756
rect 5400 14406 5428 14750
rect 5388 14400 5440 14406
rect 5388 14342 5440 14348
rect 5492 14270 5520 14972
rect 5848 14332 5900 14338
rect 5848 14274 5900 14280
rect 5480 14264 5532 14270
rect 5480 14206 5532 14212
rect 5296 14128 5348 14134
rect 5296 14070 5348 14076
rect 5308 13708 5336 14070
rect 5388 13720 5440 13726
rect 5308 13680 5388 13708
rect 5388 13662 5440 13668
rect 5400 13250 5428 13662
rect 5388 13244 5440 13250
rect 5388 13186 5440 13192
rect 5860 12638 5888 14274
rect 5848 12632 5900 12638
rect 5848 12574 5900 12580
rect 5112 12156 5164 12162
rect 5112 12098 5164 12104
rect 5952 11958 5980 18490
rect 6136 18282 6164 20695
rect 6320 19914 6348 20870
rect 6412 20322 6440 21278
rect 6400 20316 6452 20322
rect 6400 20258 6452 20264
rect 6676 20248 6728 20254
rect 6676 20190 6728 20196
rect 6308 19908 6360 19914
rect 6308 19850 6360 19856
rect 6688 19710 6716 20190
rect 6872 20186 6900 22520
rect 6952 22502 7004 22508
rect 7056 22362 7084 23454
rect 7148 23178 7176 23522
rect 7320 23376 7372 23382
rect 7320 23318 7372 23324
rect 7136 23172 7188 23178
rect 7136 23114 7188 23120
rect 7332 22974 7360 23318
rect 7320 22968 7372 22974
rect 7320 22910 7372 22916
rect 7044 22356 7096 22362
rect 7044 22298 7096 22304
rect 7228 21540 7280 21546
rect 7228 21482 7280 21488
rect 7044 21472 7096 21478
rect 7044 21414 7096 21420
rect 6952 21200 7004 21206
rect 6952 21142 7004 21148
rect 6964 20662 6992 21142
rect 7056 20730 7084 21414
rect 7240 20866 7268 21482
rect 7228 20860 7280 20866
rect 7280 20820 7452 20848
rect 7228 20802 7280 20808
rect 7044 20724 7096 20730
rect 7044 20666 7096 20672
rect 6952 20656 7004 20662
rect 6952 20598 7004 20604
rect 6860 20180 6912 20186
rect 6860 20122 6912 20128
rect 6676 19704 6728 19710
rect 6676 19646 6728 19652
rect 6492 19296 6544 19302
rect 6492 19238 6544 19244
rect 6308 19228 6360 19234
rect 6308 19170 6360 19176
rect 6320 18826 6348 19170
rect 6504 18826 6532 19238
rect 6308 18820 6360 18826
rect 6308 18762 6360 18768
rect 6492 18820 6544 18826
rect 6492 18762 6544 18768
rect 6124 18276 6176 18282
rect 6124 18218 6176 18224
rect 6320 18010 6348 18762
rect 6688 18622 6716 19646
rect 6676 18616 6728 18622
rect 6676 18558 6728 18564
rect 6492 18140 6544 18146
rect 6492 18082 6544 18088
rect 6308 18004 6360 18010
rect 6308 17946 6360 17952
rect 6504 17738 6532 18082
rect 6688 18078 6716 18558
rect 6676 18072 6728 18078
rect 6676 18014 6728 18020
rect 6688 17738 6716 18014
rect 6768 17936 6820 17942
rect 6768 17878 6820 17884
rect 6780 17738 6808 17878
rect 6492 17732 6544 17738
rect 6492 17674 6544 17680
rect 6676 17732 6728 17738
rect 6676 17674 6728 17680
rect 6768 17732 6820 17738
rect 6768 17674 6820 17680
rect 6768 16984 6820 16990
rect 6768 16926 6820 16932
rect 6780 16310 6808 16926
rect 6872 16514 6900 20122
rect 6964 18298 6992 20598
rect 7056 20322 7084 20666
rect 7136 20656 7188 20662
rect 7136 20598 7188 20604
rect 7044 20316 7096 20322
rect 7044 20258 7096 20264
rect 7056 19370 7084 20258
rect 7148 19642 7176 20598
rect 7320 20316 7372 20322
rect 7240 20276 7320 20304
rect 7240 19914 7268 20276
rect 7320 20258 7372 20264
rect 7320 20180 7372 20186
rect 7320 20122 7372 20128
rect 7228 19908 7280 19914
rect 7228 19850 7280 19856
rect 7332 19846 7360 20122
rect 7320 19840 7372 19846
rect 7320 19782 7372 19788
rect 7136 19636 7188 19642
rect 7136 19578 7188 19584
rect 7044 19364 7096 19370
rect 7044 19306 7096 19312
rect 6964 18270 7084 18298
rect 6952 18208 7004 18214
rect 6952 18150 7004 18156
rect 6964 17738 6992 18150
rect 6952 17732 7004 17738
rect 6952 17674 7004 17680
rect 6860 16508 6912 16514
rect 6860 16450 6912 16456
rect 6768 16304 6820 16310
rect 6768 16246 6820 16252
rect 6780 16038 6808 16246
rect 6768 16032 6820 16038
rect 6768 15974 6820 15980
rect 6308 15964 6360 15970
rect 6492 15964 6544 15970
rect 6360 15924 6440 15952
rect 6308 15906 6360 15912
rect 6412 15290 6440 15924
rect 6492 15906 6544 15912
rect 6504 15562 6532 15906
rect 6952 15896 7004 15902
rect 6952 15838 7004 15844
rect 6964 15562 6992 15838
rect 7056 15834 7084 18270
rect 7148 16990 7176 19578
rect 7332 18146 7360 19782
rect 7424 19710 7452 20820
rect 7412 19704 7464 19710
rect 7412 19646 7464 19652
rect 7424 19302 7452 19646
rect 7412 19296 7464 19302
rect 7412 19238 7464 19244
rect 7320 18140 7372 18146
rect 7320 18082 7372 18088
rect 7228 17936 7280 17942
rect 7228 17878 7280 17884
rect 7240 17398 7268 17878
rect 7228 17392 7280 17398
rect 7228 17334 7280 17340
rect 7136 16984 7188 16990
rect 7136 16926 7188 16932
rect 7240 16446 7268 17334
rect 7412 17052 7464 17058
rect 7412 16994 7464 17000
rect 7424 16650 7452 16994
rect 7412 16644 7464 16650
rect 7412 16586 7464 16592
rect 7228 16440 7280 16446
rect 7228 16382 7280 16388
rect 7320 16372 7372 16378
rect 7320 16314 7372 16320
rect 7332 16106 7360 16314
rect 7320 16100 7372 16106
rect 7320 16042 7372 16048
rect 7424 15902 7452 16586
rect 7412 15896 7464 15902
rect 7412 15838 7464 15844
rect 7044 15828 7096 15834
rect 7044 15770 7096 15776
rect 6492 15556 6544 15562
rect 6492 15498 6544 15504
rect 6952 15556 7004 15562
rect 6952 15498 7004 15504
rect 6400 15284 6452 15290
rect 6400 15226 6452 15232
rect 6412 14882 6440 15226
rect 6504 15018 6532 15498
rect 6492 15012 6544 15018
rect 6492 14954 6544 14960
rect 6400 14876 6452 14882
rect 6400 14818 6452 14824
rect 6412 14134 6440 14818
rect 6504 14474 6532 14954
rect 6676 14672 6728 14678
rect 6676 14614 6728 14620
rect 6688 14474 6716 14614
rect 6492 14468 6544 14474
rect 6492 14410 6544 14416
rect 6676 14468 6728 14474
rect 6676 14410 6728 14416
rect 6400 14128 6452 14134
rect 6400 14070 6452 14076
rect 7412 12700 7464 12706
rect 7412 12642 7464 12648
rect 6124 12632 6176 12638
rect 6124 12574 6176 12580
rect 6308 12632 6360 12638
rect 6308 12574 6360 12580
rect 6136 12094 6164 12574
rect 6320 12298 6348 12574
rect 6308 12292 6360 12298
rect 6308 12234 6360 12240
rect 6124 12088 6176 12094
rect 6124 12030 6176 12036
rect 4836 11952 4888 11958
rect 4836 11894 4888 11900
rect 5940 11952 5992 11958
rect 5940 11894 5992 11900
rect 4744 8892 4796 8898
rect 4744 8834 4796 8840
rect 4468 8824 4520 8830
rect 4468 8766 4520 8772
rect 4848 6858 4876 11894
rect 5952 10870 5980 11894
rect 6136 11006 6164 12030
rect 6320 11754 6348 12234
rect 6584 12088 6636 12094
rect 6584 12030 6636 12036
rect 6768 12088 6820 12094
rect 6768 12030 6820 12036
rect 6308 11748 6360 11754
rect 6308 11690 6360 11696
rect 6596 11482 6624 12030
rect 6780 11550 6808 12030
rect 6768 11544 6820 11550
rect 6768 11486 6820 11492
rect 6584 11476 6636 11482
rect 6584 11418 6636 11424
rect 6400 11408 6452 11414
rect 6400 11350 6452 11356
rect 6412 11074 6440 11350
rect 6400 11068 6452 11074
rect 6400 11010 6452 11016
rect 6124 11000 6176 11006
rect 6124 10942 6176 10948
rect 5664 10864 5716 10870
rect 5664 10806 5716 10812
rect 5940 10864 5992 10870
rect 5940 10806 5992 10812
rect 5676 9782 5704 10806
rect 6136 10326 6164 10942
rect 6412 10598 6440 11010
rect 7424 10938 7452 12642
rect 7412 10932 7464 10938
rect 7332 10892 7412 10920
rect 6400 10592 6452 10598
rect 6400 10534 6452 10540
rect 7044 10592 7096 10598
rect 7044 10534 7096 10540
rect 6124 10320 6176 10326
rect 6124 10262 6176 10268
rect 7056 10122 7084 10534
rect 7044 10116 7096 10122
rect 7044 10058 7096 10064
rect 5664 9776 5716 9782
rect 5664 9718 5716 9724
rect 5480 9504 5532 9510
rect 5480 9446 5532 9452
rect 5492 9034 5520 9446
rect 5572 9436 5624 9442
rect 5572 9378 5624 9384
rect 5480 9028 5532 9034
rect 5480 8970 5532 8976
rect 5480 8688 5532 8694
rect 5584 8676 5612 9378
rect 5532 8648 5612 8676
rect 5480 8630 5532 8636
rect 5296 8416 5348 8422
rect 5296 8358 5348 8364
rect 5308 7946 5336 8358
rect 5492 8354 5520 8630
rect 5676 8506 5704 9718
rect 6032 9368 6084 9374
rect 6032 9310 6084 9316
rect 6044 9209 6072 9310
rect 6492 9232 6544 9238
rect 6030 9200 6086 9209
rect 6492 9174 6544 9180
rect 6030 9135 6086 9144
rect 6044 8966 6072 9135
rect 6032 8960 6084 8966
rect 6032 8902 6084 8908
rect 6504 8898 6532 9174
rect 6492 8892 6544 8898
rect 6492 8834 6544 8840
rect 6124 8824 6176 8830
rect 6124 8766 6176 8772
rect 5584 8478 5704 8506
rect 5480 8348 5532 8354
rect 5480 8290 5532 8296
rect 5296 7940 5348 7946
rect 5296 7882 5348 7888
rect 5492 7606 5520 8290
rect 5480 7600 5532 7606
rect 5480 7542 5532 7548
rect 5492 7266 5520 7542
rect 5296 7260 5348 7266
rect 5296 7202 5348 7208
rect 5480 7260 5532 7266
rect 5480 7202 5532 7208
rect 5308 6858 5336 7202
rect 4836 6852 4888 6858
rect 4836 6794 4888 6800
rect 5296 6852 5348 6858
rect 5296 6794 5348 6800
rect 4282 6616 4338 6625
rect 4834 6616 4890 6625
rect 4282 6551 4338 6560
rect 4376 6580 4428 6586
rect 4834 6551 4890 6560
rect 4376 6522 4428 6528
rect 2904 6512 2956 6518
rect 2904 6454 2956 6460
rect 3088 6512 3140 6518
rect 3088 6454 3140 6460
rect 3916 6512 3968 6518
rect 4100 6512 4152 6518
rect 3968 6472 4048 6500
rect 3916 6454 3968 6460
rect 1800 6104 1852 6110
rect 1800 6046 1852 6052
rect 2168 6104 2220 6110
rect 2168 6046 2220 6052
rect 972 5492 1024 5498
rect 972 5434 1024 5440
rect 1432 5492 1484 5498
rect 1432 5434 1484 5440
rect 880 5220 932 5226
rect 880 5162 932 5168
rect 984 5158 1012 5434
rect 1444 5226 1472 5434
rect 1432 5220 1484 5226
rect 1432 5162 1484 5168
rect 972 5152 1024 5158
rect 972 5094 1024 5100
rect 2180 5090 2208 6046
rect 1616 5084 1668 5090
rect 1616 5026 1668 5032
rect 2168 5084 2220 5090
rect 2168 5026 2220 5032
rect 1628 4682 1656 5026
rect 1984 5016 2036 5022
rect 1984 4958 2036 4964
rect 1996 4682 2024 4958
rect 2180 4682 2208 5026
rect 2916 5022 2944 6454
rect 3100 6178 3128 6454
rect 3364 6240 3416 6246
rect 3364 6182 3416 6188
rect 3088 6172 3140 6178
rect 3088 6114 3140 6120
rect 2996 5968 3048 5974
rect 2996 5910 3048 5916
rect 3008 5770 3036 5910
rect 3100 5770 3128 6114
rect 2996 5764 3048 5770
rect 2996 5706 3048 5712
rect 3088 5764 3140 5770
rect 3088 5706 3140 5712
rect 3272 5084 3324 5090
rect 3272 5026 3324 5032
rect 2352 5016 2404 5022
rect 2352 4958 2404 4964
rect 2904 5016 2956 5022
rect 2904 4958 2956 4964
rect 1616 4676 1668 4682
rect 1616 4618 1668 4624
rect 1984 4676 2036 4682
rect 1984 4618 2036 4624
rect 2168 4676 2220 4682
rect 2168 4618 2220 4624
rect 1246 4304 1302 4313
rect 1246 4239 1302 4248
rect 1260 4138 1288 4239
rect 1248 4132 1300 4138
rect 1248 4074 1300 4080
rect 1260 3594 1288 4074
rect 2364 3798 2392 4958
rect 3284 4342 3312 5026
rect 3376 4954 3404 6182
rect 3916 6104 3968 6110
rect 3916 6046 3968 6052
rect 3504 5868 3824 5888
rect 3504 5866 3516 5868
rect 3572 5866 3596 5868
rect 3652 5866 3676 5868
rect 3732 5866 3756 5868
rect 3812 5866 3824 5868
rect 3504 5814 3510 5866
rect 3572 5814 3574 5866
rect 3754 5814 3756 5866
rect 3818 5814 3824 5866
rect 3504 5812 3516 5814
rect 3572 5812 3596 5814
rect 3652 5812 3676 5814
rect 3732 5812 3756 5814
rect 3812 5812 3824 5814
rect 3504 5792 3824 5812
rect 3928 5770 3956 6046
rect 3916 5764 3968 5770
rect 3916 5706 3968 5712
rect 4020 5090 4048 6472
rect 4100 6454 4152 6460
rect 4008 5084 4060 5090
rect 3928 5044 4008 5072
rect 3364 4948 3416 4954
rect 3364 4890 3416 4896
rect 3504 4780 3824 4800
rect 3504 4778 3516 4780
rect 3572 4778 3596 4780
rect 3652 4778 3676 4780
rect 3732 4778 3756 4780
rect 3812 4778 3824 4780
rect 3504 4726 3510 4778
rect 3572 4726 3574 4778
rect 3754 4726 3756 4778
rect 3818 4726 3824 4778
rect 3504 4724 3516 4726
rect 3572 4724 3596 4726
rect 3652 4724 3676 4726
rect 3732 4724 3756 4726
rect 3812 4724 3824 4726
rect 3504 4704 3824 4724
rect 3272 4336 3324 4342
rect 3272 4278 3324 4284
rect 3284 3934 3312 4278
rect 3928 4002 3956 5044
rect 4008 5026 4060 5032
rect 4008 4948 4060 4954
rect 4008 4890 4060 4896
rect 3916 3996 3968 4002
rect 3916 3938 3968 3944
rect 3272 3928 3324 3934
rect 3272 3870 3324 3876
rect 2352 3792 2404 3798
rect 2352 3734 2404 3740
rect 2904 3792 2956 3798
rect 2904 3734 2956 3740
rect 1248 3588 1300 3594
rect 1248 3530 1300 3536
rect 2916 3390 2944 3734
rect 2904 3384 2956 3390
rect 2904 3326 2956 3332
rect 1064 3316 1116 3322
rect 1064 3258 1116 3264
rect 1076 3050 1104 3258
rect 3284 3254 3312 3870
rect 3364 3792 3416 3798
rect 3364 3734 3416 3740
rect 3376 3458 3404 3734
rect 3504 3692 3824 3712
rect 3504 3690 3516 3692
rect 3572 3690 3596 3692
rect 3652 3690 3676 3692
rect 3732 3690 3756 3692
rect 3812 3690 3824 3692
rect 3504 3638 3510 3690
rect 3572 3638 3574 3690
rect 3754 3638 3756 3690
rect 3818 3638 3824 3690
rect 3504 3636 3516 3638
rect 3572 3636 3596 3638
rect 3652 3636 3676 3638
rect 3732 3636 3756 3638
rect 3812 3636 3824 3638
rect 3504 3616 3824 3636
rect 3928 3594 3956 3938
rect 3916 3588 3968 3594
rect 3916 3530 3968 3536
rect 3364 3452 3416 3458
rect 3364 3394 3416 3400
rect 3272 3248 3324 3254
rect 3272 3190 3324 3196
rect 1064 3044 1116 3050
rect 1064 2986 1116 2992
rect 1076 2506 1104 2986
rect 1708 2704 1760 2710
rect 1708 2646 1760 2652
rect 1064 2500 1116 2506
rect 1064 2442 1116 2448
rect 1154 2400 1210 2409
rect 1720 2370 1748 2646
rect 1154 2335 1210 2344
rect 1708 2364 1760 2370
rect 972 2296 1024 2302
rect 972 2238 1024 2244
rect 984 1962 1012 2238
rect 972 1956 1024 1962
rect 972 1898 1024 1904
rect 1168 1826 1196 2335
rect 1708 2306 1760 2312
rect 1720 2234 1748 2306
rect 1708 2228 1760 2234
rect 1708 2170 1760 2176
rect 3284 2166 3312 3190
rect 3376 3050 3404 3394
rect 3916 3248 3968 3254
rect 3916 3190 3968 3196
rect 3364 3044 3416 3050
rect 3364 2986 3416 2992
rect 3928 2914 3956 3190
rect 3364 2908 3416 2914
rect 3364 2850 3416 2856
rect 3916 2908 3968 2914
rect 3916 2850 3968 2856
rect 3376 2506 3404 2850
rect 4020 2846 4048 4890
rect 4008 2840 4060 2846
rect 4008 2782 4060 2788
rect 3916 2772 3968 2778
rect 3916 2714 3968 2720
rect 3504 2604 3824 2624
rect 3504 2602 3516 2604
rect 3572 2602 3596 2604
rect 3652 2602 3676 2604
rect 3732 2602 3756 2604
rect 3812 2602 3824 2604
rect 3504 2550 3510 2602
rect 3572 2550 3574 2602
rect 3754 2550 3756 2602
rect 3818 2550 3824 2602
rect 3504 2548 3516 2550
rect 3572 2548 3596 2550
rect 3652 2548 3676 2550
rect 3732 2548 3756 2550
rect 3812 2548 3824 2550
rect 3504 2528 3824 2548
rect 3928 2506 3956 2714
rect 3364 2500 3416 2506
rect 3364 2442 3416 2448
rect 3916 2500 3968 2506
rect 4112 2488 4140 6454
rect 4388 6246 4416 6522
rect 4376 6240 4428 6246
rect 4376 6182 4428 6188
rect 4388 5226 4416 6182
rect 4848 5566 4876 6551
rect 5308 5974 5336 6794
rect 5492 6586 5520 7202
rect 5480 6580 5532 6586
rect 5480 6522 5532 6528
rect 5296 5968 5348 5974
rect 5296 5910 5348 5916
rect 4468 5560 4520 5566
rect 4468 5502 4520 5508
rect 4652 5560 4704 5566
rect 4652 5502 4704 5508
rect 4836 5560 4888 5566
rect 4836 5502 4888 5508
rect 4376 5220 4428 5226
rect 4376 5162 4428 5168
rect 4480 4886 4508 5502
rect 4560 5424 4612 5430
rect 4560 5366 4612 5372
rect 4572 5022 4600 5366
rect 4560 5016 4612 5022
rect 4560 4958 4612 4964
rect 4468 4880 4520 4886
rect 4468 4822 4520 4828
rect 4572 4614 4600 4958
rect 4664 4954 4692 5502
rect 4848 5158 4876 5502
rect 4836 5152 4888 5158
rect 4836 5094 4888 5100
rect 4744 5084 4796 5090
rect 4744 5026 4796 5032
rect 4652 4948 4704 4954
rect 4652 4890 4704 4896
rect 4560 4608 4612 4614
rect 4560 4550 4612 4556
rect 4664 4070 4692 4890
rect 4756 4682 4784 5026
rect 4928 4880 4980 4886
rect 4928 4822 4980 4828
rect 4940 4682 4968 4822
rect 4744 4676 4796 4682
rect 4744 4618 4796 4624
rect 4928 4676 4980 4682
rect 4928 4618 4980 4624
rect 4652 4064 4704 4070
rect 4652 4006 4704 4012
rect 5480 4064 5532 4070
rect 5480 4006 5532 4012
rect 4376 3588 4428 3594
rect 4376 3530 4428 3536
rect 4388 3390 4416 3530
rect 4376 3384 4428 3390
rect 4376 3326 4428 3332
rect 4664 2914 4692 4006
rect 5388 3860 5440 3866
rect 5388 3802 5440 3808
rect 5400 3594 5428 3802
rect 5492 3594 5520 4006
rect 5388 3588 5440 3594
rect 5388 3530 5440 3536
rect 5480 3588 5532 3594
rect 5480 3530 5532 3536
rect 5400 2982 5428 3530
rect 5388 2976 5440 2982
rect 5388 2918 5440 2924
rect 4468 2908 4520 2914
rect 4468 2850 4520 2856
rect 4652 2908 4704 2914
rect 4652 2850 4704 2856
rect 3916 2442 3968 2448
rect 4020 2460 4324 2488
rect 3272 2160 3324 2166
rect 3272 2102 3324 2108
rect 1708 1956 1760 1962
rect 1708 1898 1760 1904
rect 1156 1820 1208 1826
rect 1156 1762 1208 1768
rect 1168 1418 1196 1762
rect 1156 1412 1208 1418
rect 1156 1354 1208 1360
rect 418 632 474 641
rect 418 567 474 576
rect 432 424 460 567
rect 1720 424 1748 1898
rect 3928 1894 3956 2442
rect 4020 2302 4048 2460
rect 4192 2364 4244 2370
rect 4192 2306 4244 2312
rect 4008 2296 4060 2302
rect 4008 2238 4060 2244
rect 4100 2228 4152 2234
rect 4204 2216 4232 2306
rect 4296 2302 4324 2460
rect 4480 2438 4508 2850
rect 4560 2704 4612 2710
rect 4560 2646 4612 2652
rect 4468 2432 4520 2438
rect 4468 2374 4520 2380
rect 4284 2296 4336 2302
rect 4284 2238 4336 2244
rect 4152 2188 4232 2216
rect 4100 2170 4152 2176
rect 3916 1888 3968 1894
rect 3916 1830 3968 1836
rect 2168 1616 2220 1622
rect 2168 1558 2220 1564
rect 2180 1078 2208 1558
rect 3504 1516 3824 1536
rect 3504 1514 3516 1516
rect 3572 1514 3596 1516
rect 3652 1514 3676 1516
rect 3732 1514 3756 1516
rect 3812 1514 3824 1516
rect 3504 1462 3510 1514
rect 3572 1462 3574 1514
rect 3754 1462 3756 1514
rect 3818 1462 3824 1514
rect 3504 1460 3516 1462
rect 3572 1460 3596 1462
rect 3652 1460 3676 1462
rect 3732 1460 3756 1462
rect 3812 1460 3824 1462
rect 3504 1440 3824 1460
rect 3928 1418 3956 1830
rect 4572 1758 4600 2646
rect 4664 2234 4692 2850
rect 5400 2506 5428 2918
rect 5388 2500 5440 2506
rect 5388 2442 5440 2448
rect 4652 2228 4704 2234
rect 4652 2170 4704 2176
rect 5584 1962 5612 8478
rect 5848 8280 5900 8286
rect 5848 8222 5900 8228
rect 5860 8121 5888 8222
rect 6136 8150 6164 8766
rect 6216 8348 6268 8354
rect 6216 8290 6268 8296
rect 6124 8144 6176 8150
rect 5846 8112 5902 8121
rect 6124 8086 6176 8092
rect 5846 8047 5902 8056
rect 5860 7946 5888 8047
rect 5938 7976 5994 7985
rect 5848 7940 5900 7946
rect 6228 7946 6256 8290
rect 6400 8212 6452 8218
rect 6400 8154 6452 8160
rect 6412 7946 6440 8154
rect 5938 7911 5994 7920
rect 6216 7940 6268 7946
rect 5848 7882 5900 7888
rect 5952 7334 5980 7911
rect 6216 7882 6268 7888
rect 6400 7940 6452 7946
rect 6400 7882 6452 7888
rect 5940 7328 5992 7334
rect 5940 7270 5992 7276
rect 5952 6858 5980 7270
rect 6504 6858 6532 8834
rect 7332 8762 7360 10892
rect 7412 10874 7464 10880
rect 7410 10560 7466 10569
rect 7410 10495 7466 10504
rect 7424 10462 7452 10495
rect 7412 10456 7464 10462
rect 7412 10398 7464 10404
rect 7424 9986 7452 10398
rect 7412 9980 7464 9986
rect 7412 9922 7464 9928
rect 7516 9918 7544 31662
rect 8608 30720 8660 30726
rect 8608 30662 8660 30668
rect 7688 30244 7740 30250
rect 7688 30186 7740 30192
rect 7700 29706 7728 30186
rect 7688 29700 7740 29706
rect 7688 29642 7740 29648
rect 7688 28476 7740 28482
rect 7688 28418 7740 28424
rect 7596 28408 7648 28414
rect 7596 28350 7648 28356
rect 7608 27462 7636 28350
rect 7700 28278 7728 28418
rect 7688 28272 7740 28278
rect 7688 28214 7740 28220
rect 7700 28074 7728 28214
rect 7688 28068 7740 28074
rect 7688 28010 7740 28016
rect 7596 27456 7648 27462
rect 7596 27398 7648 27404
rect 7608 26986 7636 27398
rect 7596 26980 7648 26986
rect 7596 26922 7648 26928
rect 7700 25762 7728 28010
rect 7872 27728 7924 27734
rect 7872 27670 7924 27676
rect 7884 27326 7912 27670
rect 7872 27320 7924 27326
rect 7872 27262 7924 27268
rect 7884 26102 7912 27262
rect 7872 26096 7924 26102
rect 7872 26038 7924 26044
rect 8240 26096 8292 26102
rect 8240 26038 8292 26044
rect 7688 25756 7740 25762
rect 7688 25698 7740 25704
rect 8252 25082 8280 26038
rect 8240 25076 8292 25082
rect 8240 25018 8292 25024
rect 7780 24736 7832 24742
rect 7780 24678 7832 24684
rect 7688 24600 7740 24606
rect 7688 24542 7740 24548
rect 7700 23994 7728 24542
rect 7688 23988 7740 23994
rect 7688 23930 7740 23936
rect 7700 23722 7728 23930
rect 7792 23722 7820 24678
rect 7688 23716 7740 23722
rect 7688 23658 7740 23664
rect 7780 23716 7832 23722
rect 7780 23658 7832 23664
rect 7872 23172 7924 23178
rect 7872 23114 7924 23120
rect 7596 22424 7648 22430
rect 7596 22366 7648 22372
rect 7608 21546 7636 22366
rect 7780 21880 7832 21886
rect 7780 21822 7832 21828
rect 7596 21540 7648 21546
rect 7596 21482 7648 21488
rect 7596 21404 7648 21410
rect 7596 21346 7648 21352
rect 7608 19370 7636 21346
rect 7792 21274 7820 21822
rect 7780 21268 7832 21274
rect 7780 21210 7832 21216
rect 7688 20792 7740 20798
rect 7688 20734 7740 20740
rect 7700 20118 7728 20734
rect 7792 20390 7820 21210
rect 7884 21002 7912 23114
rect 8148 22968 8200 22974
rect 8148 22910 8200 22916
rect 8160 22498 8188 22910
rect 8148 22492 8200 22498
rect 8148 22434 8200 22440
rect 8160 22090 8188 22434
rect 8148 22084 8200 22090
rect 8148 22026 8200 22032
rect 7872 20996 7924 21002
rect 7872 20938 7924 20944
rect 7884 20798 7912 20938
rect 7872 20792 7924 20798
rect 7872 20734 7924 20740
rect 7780 20384 7832 20390
rect 7780 20326 7832 20332
rect 7688 20112 7740 20118
rect 7688 20054 7740 20060
rect 7884 19846 7912 20734
rect 8148 20112 8200 20118
rect 8148 20054 8200 20060
rect 7872 19840 7924 19846
rect 7872 19782 7924 19788
rect 8160 19752 8188 20054
rect 8148 19746 8200 19752
rect 8148 19688 8200 19694
rect 8516 19704 8568 19710
rect 8516 19646 8568 19652
rect 7872 19568 7924 19574
rect 7872 19510 7924 19516
rect 7596 19364 7648 19370
rect 7596 19306 7648 19312
rect 7884 19234 7912 19510
rect 8528 19370 8556 19646
rect 8516 19364 8568 19370
rect 8516 19306 8568 19312
rect 7872 19228 7924 19234
rect 7872 19170 7924 19176
rect 8424 17528 8476 17534
rect 8424 17470 8476 17476
rect 8436 17369 8464 17470
rect 8422 17360 8478 17369
rect 8422 17295 8478 17304
rect 7596 16984 7648 16990
rect 7596 16926 7648 16932
rect 7608 16650 7636 16926
rect 7596 16644 7648 16650
rect 7596 16586 7648 16592
rect 8240 16508 8292 16514
rect 8240 16450 8292 16456
rect 7964 16372 8016 16378
rect 7964 16314 8016 16320
rect 7688 15964 7740 15970
rect 7688 15906 7740 15912
rect 7700 15290 7728 15906
rect 7976 15562 8004 16314
rect 8252 16038 8280 16450
rect 8424 16440 8476 16446
rect 8424 16382 8476 16388
rect 8436 16038 8464 16382
rect 8240 16032 8292 16038
rect 8240 15974 8292 15980
rect 8424 16032 8476 16038
rect 8424 15974 8476 15980
rect 7964 15556 8016 15562
rect 7964 15498 8016 15504
rect 7780 15420 7832 15426
rect 7780 15362 7832 15368
rect 7688 15284 7740 15290
rect 7688 15226 7740 15232
rect 7792 15018 7820 15362
rect 7976 15018 8004 15498
rect 8252 15426 8280 15974
rect 8332 15828 8384 15834
rect 8332 15770 8384 15776
rect 8240 15420 8292 15426
rect 8240 15362 8292 15368
rect 8344 15358 8372 15770
rect 8332 15352 8384 15358
rect 8332 15294 8384 15300
rect 8344 15018 8372 15294
rect 7780 15012 7832 15018
rect 7780 14954 7832 14960
rect 7964 15012 8016 15018
rect 7964 14954 8016 14960
rect 8332 15012 8384 15018
rect 8332 14954 8384 14960
rect 8238 14232 8294 14241
rect 8238 14167 8240 14176
rect 8292 14167 8294 14176
rect 8240 14138 8292 14144
rect 8054 13688 8110 13697
rect 8054 13623 8110 13632
rect 8068 12774 8096 13623
rect 8056 12768 8108 12774
rect 8056 12710 8108 12716
rect 7964 12700 8016 12706
rect 7964 12642 8016 12648
rect 7872 12020 7924 12026
rect 7872 11962 7924 11968
rect 7688 11952 7740 11958
rect 7688 11894 7740 11900
rect 7596 11476 7648 11482
rect 7596 11418 7648 11424
rect 7608 11142 7636 11418
rect 7700 11210 7728 11894
rect 7688 11204 7740 11210
rect 7688 11146 7740 11152
rect 7596 11136 7648 11142
rect 7596 11078 7648 11084
rect 7608 10462 7636 11078
rect 7596 10456 7648 10462
rect 7596 10398 7648 10404
rect 7608 10122 7636 10398
rect 7596 10116 7648 10122
rect 7596 10058 7648 10064
rect 7596 9980 7648 9986
rect 7596 9922 7648 9928
rect 7504 9912 7556 9918
rect 7504 9854 7556 9860
rect 7412 8892 7464 8898
rect 7412 8834 7464 8840
rect 7320 8756 7372 8762
rect 7320 8698 7372 8704
rect 7136 8348 7188 8354
rect 7136 8290 7188 8296
rect 6860 8280 6912 8286
rect 6860 8222 6912 8228
rect 6952 8280 7004 8286
rect 6952 8222 7004 8228
rect 6872 7946 6900 8222
rect 6860 7940 6912 7946
rect 6860 7882 6912 7888
rect 6768 7600 6820 7606
rect 6768 7542 6820 7548
rect 6780 7334 6808 7542
rect 6964 7402 6992 8222
rect 7044 8144 7096 8150
rect 7044 8086 7096 8092
rect 7056 7742 7084 8086
rect 7044 7736 7096 7742
rect 7044 7678 7096 7684
rect 6952 7396 7004 7402
rect 6952 7338 7004 7344
rect 6768 7328 6820 7334
rect 6768 7270 6820 7276
rect 5940 6852 5992 6858
rect 5940 6794 5992 6800
rect 6492 6852 6544 6858
rect 6492 6794 6544 6800
rect 6584 6580 6636 6586
rect 6584 6522 6636 6528
rect 6676 6580 6728 6586
rect 6676 6522 6728 6528
rect 6596 6110 6624 6522
rect 5664 6104 5716 6110
rect 5664 6046 5716 6052
rect 6584 6104 6636 6110
rect 6584 6046 6636 6052
rect 5676 5498 5704 6046
rect 5664 5492 5716 5498
rect 5664 5434 5716 5440
rect 5940 5492 5992 5498
rect 5940 5434 5992 5440
rect 5952 4614 5980 5434
rect 6596 5430 6624 6046
rect 6688 5566 6716 6522
rect 6768 6172 6820 6178
rect 6768 6114 6820 6120
rect 6780 5566 6808 6114
rect 6964 5770 6992 7338
rect 7148 6790 7176 8290
rect 7228 7804 7280 7810
rect 7228 7746 7280 7752
rect 7240 7402 7268 7746
rect 7228 7396 7280 7402
rect 7228 7338 7280 7344
rect 7424 6790 7452 8834
rect 7504 7736 7556 7742
rect 7504 7678 7556 7684
rect 7516 7402 7544 7678
rect 7504 7396 7556 7402
rect 7504 7338 7556 7344
rect 7136 6784 7188 6790
rect 7136 6726 7188 6732
rect 7412 6784 7464 6790
rect 7412 6726 7464 6732
rect 6952 5764 7004 5770
rect 6952 5706 7004 5712
rect 6676 5560 6728 5566
rect 6676 5502 6728 5508
rect 6768 5560 6820 5566
rect 6768 5502 6820 5508
rect 7504 5560 7556 5566
rect 7504 5502 7556 5508
rect 6584 5424 6636 5430
rect 6584 5366 6636 5372
rect 5940 4608 5992 4614
rect 5940 4550 5992 4556
rect 5952 4002 5980 4550
rect 6596 4478 6624 5366
rect 7516 5090 7544 5502
rect 7320 5084 7372 5090
rect 7320 5026 7372 5032
rect 7504 5084 7556 5090
rect 7504 5026 7556 5032
rect 6584 4472 6636 4478
rect 6584 4414 6636 4420
rect 6596 4342 6624 4414
rect 7332 4342 7360 5026
rect 7516 4682 7544 5026
rect 7504 4676 7556 4682
rect 7504 4618 7556 4624
rect 6400 4336 6452 4342
rect 6400 4278 6452 4284
rect 6584 4336 6636 4342
rect 6584 4278 6636 4284
rect 7136 4336 7188 4342
rect 7136 4278 7188 4284
rect 7320 4336 7372 4342
rect 7320 4278 7372 4284
rect 7504 4336 7556 4342
rect 7504 4278 7556 4284
rect 6412 4138 6440 4278
rect 6400 4132 6452 4138
rect 6400 4074 6452 4080
rect 7148 4002 7176 4278
rect 5664 3996 5716 4002
rect 5664 3938 5716 3944
rect 5940 3996 5992 4002
rect 5940 3938 5992 3944
rect 6952 3996 7004 4002
rect 6952 3938 7004 3944
rect 7136 3996 7188 4002
rect 7136 3938 7188 3944
rect 5676 3594 5704 3938
rect 5664 3588 5716 3594
rect 5664 3530 5716 3536
rect 5676 3254 5704 3530
rect 5952 3526 5980 3938
rect 6964 3594 6992 3938
rect 7148 3594 7176 3938
rect 6952 3588 7004 3594
rect 6952 3530 7004 3536
rect 7136 3588 7188 3594
rect 7136 3530 7188 3536
rect 5940 3520 5992 3526
rect 5940 3462 5992 3468
rect 5848 3452 5900 3458
rect 5848 3394 5900 3400
rect 5664 3248 5716 3254
rect 5664 3190 5716 3196
rect 5676 3050 5704 3190
rect 5664 3044 5716 3050
rect 5664 2986 5716 2992
rect 5572 1956 5624 1962
rect 5572 1898 5624 1904
rect 5860 1894 5888 3394
rect 6032 3384 6084 3390
rect 6032 3326 6084 3332
rect 6044 3254 6072 3326
rect 7516 3254 7544 4278
rect 7608 4070 7636 9922
rect 7700 8393 7728 11146
rect 7884 11074 7912 11962
rect 7976 11958 8004 12642
rect 8068 12094 8096 12710
rect 8516 12496 8568 12502
rect 8516 12438 8568 12444
rect 8528 12162 8556 12438
rect 8148 12156 8200 12162
rect 8148 12098 8200 12104
rect 8516 12156 8568 12162
rect 8516 12098 8568 12104
rect 8056 12088 8108 12094
rect 8056 12030 8108 12036
rect 7964 11952 8016 11958
rect 7964 11894 8016 11900
rect 8160 11754 8188 12098
rect 8148 11748 8200 11754
rect 8148 11690 8200 11696
rect 7872 11068 7924 11074
rect 7872 11010 7924 11016
rect 7780 10864 7832 10870
rect 7780 10806 7832 10812
rect 7792 10462 7820 10806
rect 7884 10530 7912 11010
rect 7872 10524 7924 10530
rect 7872 10466 7924 10472
rect 7780 10456 7832 10462
rect 7780 10398 7832 10404
rect 7792 9850 7820 10398
rect 7884 10054 7912 10466
rect 8160 10326 8188 11690
rect 8528 11686 8556 12098
rect 8516 11680 8568 11686
rect 8516 11622 8568 11628
rect 8148 10320 8200 10326
rect 8148 10262 8200 10268
rect 7872 10048 7924 10054
rect 7872 9990 7924 9996
rect 8160 9986 8188 10262
rect 8148 9980 8200 9986
rect 8148 9922 8200 9928
rect 8424 9912 8476 9918
rect 8424 9854 8476 9860
rect 7780 9844 7832 9850
rect 7780 9786 7832 9792
rect 7872 8960 7924 8966
rect 7872 8902 7924 8908
rect 7780 8688 7832 8694
rect 7780 8630 7832 8636
rect 7686 8384 7742 8393
rect 7686 8319 7742 8328
rect 7792 7674 7820 8630
rect 7884 8354 7912 8902
rect 8436 8898 8464 9854
rect 8620 9481 8648 30662
rect 9448 30522 9476 31664
rect 9988 30584 10040 30590
rect 9988 30526 10040 30532
rect 9436 30516 9488 30522
rect 9436 30458 9488 30464
rect 9896 30516 9948 30522
rect 9896 30458 9948 30464
rect 9160 30176 9212 30182
rect 9160 30118 9212 30124
rect 8976 30108 9028 30114
rect 8976 30050 9028 30056
rect 8988 29706 9016 30050
rect 8976 29700 9028 29706
rect 8976 29642 9028 29648
rect 8976 29496 9028 29502
rect 8976 29438 9028 29444
rect 8792 29428 8844 29434
rect 8792 29370 8844 29376
rect 8804 28006 8832 29370
rect 8988 29026 9016 29438
rect 9068 29428 9120 29434
rect 9068 29370 9120 29376
rect 9080 29026 9108 29370
rect 9172 29366 9200 30118
rect 9160 29360 9212 29366
rect 9160 29302 9212 29308
rect 8976 29020 9028 29026
rect 8976 28962 9028 28968
rect 9068 29020 9120 29026
rect 9068 28962 9120 28968
rect 8884 28816 8936 28822
rect 8884 28758 8936 28764
rect 8792 28000 8844 28006
rect 8792 27942 8844 27948
rect 8896 27802 8924 28758
rect 8988 28618 9016 28962
rect 8976 28612 9028 28618
rect 8976 28554 9028 28560
rect 9172 28550 9200 29302
rect 9528 28884 9580 28890
rect 9528 28826 9580 28832
rect 9160 28544 9212 28550
rect 9160 28486 9212 28492
rect 9540 28482 9568 28826
rect 9528 28476 9580 28482
rect 9580 28436 9660 28464
rect 9528 28418 9580 28424
rect 9068 28408 9120 28414
rect 9068 28350 9120 28356
rect 9080 28074 9108 28350
rect 9436 28340 9488 28346
rect 9436 28282 9488 28288
rect 9068 28068 9120 28074
rect 9068 28010 9120 28016
rect 9252 28068 9304 28074
rect 9252 28010 9304 28016
rect 8884 27796 8936 27802
rect 8884 27738 8936 27744
rect 8896 27326 8924 27738
rect 9264 27326 9292 28010
rect 9448 27938 9476 28282
rect 9344 27932 9396 27938
rect 9344 27874 9396 27880
rect 9436 27932 9488 27938
rect 9436 27874 9488 27880
rect 9356 27394 9384 27874
rect 9448 27530 9476 27874
rect 9436 27524 9488 27530
rect 9436 27466 9488 27472
rect 9344 27388 9396 27394
rect 9344 27330 9396 27336
rect 8700 27320 8752 27326
rect 8700 27262 8752 27268
rect 8884 27320 8936 27326
rect 8884 27262 8936 27268
rect 9252 27320 9304 27326
rect 9252 27262 9304 27268
rect 8712 26986 8740 27262
rect 8700 26980 8752 26986
rect 8700 26922 8752 26928
rect 9264 26238 9292 27262
rect 9632 26782 9660 28436
rect 9804 26844 9856 26850
rect 9804 26786 9856 26792
rect 9620 26776 9672 26782
rect 9620 26718 9672 26724
rect 8700 26232 8752 26238
rect 8700 26174 8752 26180
rect 9252 26232 9304 26238
rect 9252 26174 9304 26180
rect 8712 25898 8740 26174
rect 8700 25892 8752 25898
rect 8700 25834 8752 25840
rect 9632 25558 9660 26718
rect 9816 26442 9844 26786
rect 9804 26436 9856 26442
rect 9804 26378 9856 26384
rect 9804 25756 9856 25762
rect 9804 25698 9856 25704
rect 9620 25552 9672 25558
rect 9620 25494 9672 25500
rect 9632 25257 9660 25494
rect 9618 25248 9674 25257
rect 9618 25183 9674 25192
rect 9252 24668 9304 24674
rect 9252 24610 9304 24616
rect 9068 24260 9120 24266
rect 9068 24202 9120 24208
rect 9080 23586 9108 24202
rect 9264 24130 9292 24610
rect 9528 24464 9580 24470
rect 9528 24406 9580 24412
rect 9540 24266 9568 24406
rect 9528 24260 9580 24266
rect 9528 24202 9580 24208
rect 9632 24130 9660 25183
rect 9252 24124 9304 24130
rect 9252 24066 9304 24072
rect 9620 24124 9672 24130
rect 9620 24066 9672 24072
rect 9068 23580 9120 23586
rect 9068 23522 9120 23528
rect 9080 22906 9108 23522
rect 9528 23512 9580 23518
rect 9528 23454 9580 23460
rect 9068 22900 9120 22906
rect 9068 22842 9120 22848
rect 9540 22838 9568 23454
rect 9528 22832 9580 22838
rect 9528 22774 9580 22780
rect 8700 21744 8752 21750
rect 8700 21686 8752 21692
rect 8712 20934 8740 21686
rect 9068 21200 9120 21206
rect 9068 21142 9120 21148
rect 8700 20928 8752 20934
rect 8700 20870 8752 20876
rect 8712 20458 8740 20870
rect 9080 20798 9108 21142
rect 9540 20798 9568 22774
rect 9068 20792 9120 20798
rect 9068 20734 9120 20740
rect 9528 20792 9580 20798
rect 9528 20734 9580 20740
rect 9080 20458 9108 20734
rect 8700 20452 8752 20458
rect 8700 20394 8752 20400
rect 9068 20452 9120 20458
rect 9068 20394 9120 20400
rect 8976 20248 9028 20254
rect 8976 20190 9028 20196
rect 8988 19574 9016 20190
rect 8976 19568 9028 19574
rect 8976 19510 9028 19516
rect 8988 18690 9016 19510
rect 9080 19370 9108 20394
rect 9252 20316 9304 20322
rect 9252 20258 9304 20264
rect 9264 19914 9292 20258
rect 9252 19908 9304 19914
rect 9252 19850 9304 19856
rect 9540 19846 9568 20734
rect 9816 20662 9844 25698
rect 9804 20656 9856 20662
rect 9804 20598 9856 20604
rect 9804 20112 9856 20118
rect 9804 20054 9856 20060
rect 9816 19914 9844 20054
rect 9804 19908 9856 19914
rect 9804 19850 9856 19856
rect 9528 19840 9580 19846
rect 9528 19782 9580 19788
rect 9528 19704 9580 19710
rect 9528 19646 9580 19652
rect 9540 19574 9568 19646
rect 9528 19568 9580 19574
rect 9528 19510 9580 19516
rect 9068 19364 9120 19370
rect 9068 19306 9120 19312
rect 9816 18758 9844 19850
rect 9804 18752 9856 18758
rect 9804 18694 9856 18700
rect 8976 18684 9028 18690
rect 8976 18626 9028 18632
rect 9068 17460 9120 17466
rect 9068 17402 9120 17408
rect 9080 17058 9108 17402
rect 9068 17052 9120 17058
rect 9068 16994 9120 17000
rect 9160 17052 9212 17058
rect 9160 16994 9212 17000
rect 8792 16032 8844 16038
rect 8792 15974 8844 15980
rect 8804 13182 8832 15974
rect 9080 15834 9108 16994
rect 9172 16038 9200 16994
rect 9804 16984 9856 16990
rect 9804 16926 9856 16932
rect 9528 16916 9580 16922
rect 9528 16858 9580 16864
rect 9160 16032 9212 16038
rect 9160 15974 9212 15980
rect 9068 15828 9120 15834
rect 9068 15770 9120 15776
rect 9540 15766 9568 16858
rect 9712 16848 9764 16854
rect 9712 16790 9764 16796
rect 9724 16446 9752 16790
rect 9712 16440 9764 16446
rect 9712 16382 9764 16388
rect 9816 16106 9844 16926
rect 9804 16100 9856 16106
rect 9804 16042 9856 16048
rect 9528 15760 9580 15766
rect 9528 15702 9580 15708
rect 9540 15494 9568 15702
rect 9528 15488 9580 15494
rect 9528 15430 9580 15436
rect 8792 13176 8844 13182
rect 8792 13118 8844 13124
rect 9908 13046 9936 30458
rect 10000 29502 10028 30526
rect 10172 30448 10224 30454
rect 10172 30390 10224 30396
rect 9988 29496 10040 29502
rect 9988 29438 10040 29444
rect 10080 28612 10132 28618
rect 10080 28554 10132 28560
rect 9988 27252 10040 27258
rect 9988 27194 10040 27200
rect 10000 26850 10028 27194
rect 9988 26844 10040 26850
rect 9988 26786 10040 26792
rect 10000 25898 10028 26786
rect 9988 25892 10040 25898
rect 9988 25834 10040 25840
rect 10092 23874 10120 28554
rect 10184 25642 10212 30390
rect 10264 30176 10316 30182
rect 10264 30118 10316 30124
rect 10276 29570 10304 30118
rect 10356 29700 10408 29706
rect 10356 29642 10408 29648
rect 10264 29564 10316 29570
rect 10264 29506 10316 29512
rect 10368 29434 10396 29642
rect 10920 29570 10948 31664
rect 11000 30040 11052 30046
rect 11000 29982 11052 29988
rect 10908 29564 10960 29570
rect 10908 29506 10960 29512
rect 10356 29428 10408 29434
rect 10356 29370 10408 29376
rect 10368 27938 10396 29370
rect 11012 29026 11040 29982
rect 11828 29496 11880 29502
rect 11828 29438 11880 29444
rect 11840 29026 11868 29438
rect 12208 29394 12236 31664
rect 13392 30652 13444 30658
rect 13392 30594 13444 30600
rect 12564 30108 12616 30114
rect 12564 30050 12616 30056
rect 12288 30040 12340 30046
rect 12288 29982 12340 29988
rect 12300 29502 12328 29982
rect 12576 29570 12604 30050
rect 13024 29972 13076 29978
rect 13024 29914 13076 29920
rect 12564 29564 12616 29570
rect 12564 29506 12616 29512
rect 13036 29502 13064 29914
rect 13208 29904 13260 29910
rect 13208 29846 13260 29852
rect 12288 29496 12340 29502
rect 12288 29438 12340 29444
rect 13024 29496 13076 29502
rect 13024 29438 13076 29444
rect 12208 29366 12512 29394
rect 13220 29366 13248 29846
rect 13300 29428 13352 29434
rect 13300 29370 13352 29376
rect 11000 29020 11052 29026
rect 11000 28962 11052 28968
rect 11828 29020 11880 29026
rect 11828 28962 11880 28968
rect 10448 28816 10500 28822
rect 10448 28758 10500 28764
rect 10460 28414 10488 28758
rect 11012 28550 11040 28962
rect 11840 28550 11868 28962
rect 11920 28952 11972 28958
rect 11920 28894 11972 28900
rect 11000 28544 11052 28550
rect 11000 28486 11052 28492
rect 11828 28544 11880 28550
rect 11828 28486 11880 28492
rect 10448 28408 10500 28414
rect 10448 28350 10500 28356
rect 11012 28278 11040 28486
rect 10540 28272 10592 28278
rect 10540 28214 10592 28220
rect 11000 28272 11052 28278
rect 11000 28214 11052 28220
rect 11276 28272 11328 28278
rect 11276 28214 11328 28220
rect 10552 28074 10580 28214
rect 10540 28068 10592 28074
rect 10540 28010 10592 28016
rect 10356 27932 10408 27938
rect 10356 27874 10408 27880
rect 10368 27530 10396 27874
rect 10356 27524 10408 27530
rect 10356 27466 10408 27472
rect 10552 26986 10580 28010
rect 10816 27864 10868 27870
rect 10816 27806 10868 27812
rect 10828 27530 10856 27806
rect 10816 27524 10868 27530
rect 10816 27466 10868 27472
rect 10632 27388 10684 27394
rect 10632 27330 10684 27336
rect 10540 26980 10592 26986
rect 10540 26922 10592 26928
rect 10356 26776 10408 26782
rect 10356 26718 10408 26724
rect 10368 25762 10396 26718
rect 10552 26238 10580 26922
rect 10644 26850 10672 27330
rect 10828 26918 10856 27466
rect 11012 27326 11040 28214
rect 11288 28006 11316 28214
rect 11276 28000 11328 28006
rect 11276 27942 11328 27948
rect 11288 27530 11316 27942
rect 11276 27524 11328 27530
rect 11276 27466 11328 27472
rect 11000 27320 11052 27326
rect 11000 27262 11052 27268
rect 10816 26912 10868 26918
rect 10816 26854 10868 26860
rect 10632 26844 10684 26850
rect 10632 26786 10684 26792
rect 10644 26306 10672 26786
rect 10828 26374 10856 26854
rect 11840 26442 11868 28486
rect 11932 28278 11960 28894
rect 11920 28272 11972 28278
rect 11920 28214 11972 28220
rect 12288 27184 12340 27190
rect 12288 27126 12340 27132
rect 11828 26436 11880 26442
rect 11828 26378 11880 26384
rect 10816 26368 10868 26374
rect 10816 26310 10868 26316
rect 10632 26300 10684 26306
rect 10632 26242 10684 26248
rect 11840 26238 11868 26378
rect 10540 26232 10592 26238
rect 10540 26174 10592 26180
rect 11828 26232 11880 26238
rect 11828 26174 11880 26180
rect 10724 26164 10776 26170
rect 10724 26106 10776 26112
rect 10356 25756 10408 25762
rect 10356 25698 10408 25704
rect 10184 25614 10396 25642
rect 10000 23846 10120 23874
rect 10262 23888 10318 23897
rect 10000 23722 10028 23846
rect 10368 23874 10396 25614
rect 10632 25620 10684 25626
rect 10632 25562 10684 25568
rect 10448 25212 10500 25218
rect 10448 25154 10500 25160
rect 10460 24266 10488 25154
rect 10448 24260 10500 24266
rect 10448 24202 10500 24208
rect 10460 24062 10488 24202
rect 10448 24056 10500 24062
rect 10448 23998 10500 24004
rect 10368 23846 10488 23874
rect 10262 23823 10318 23832
rect 9988 23716 10040 23722
rect 9988 23658 10040 23664
rect 10276 23178 10304 23823
rect 10264 23172 10316 23178
rect 10264 23114 10316 23120
rect 9988 22492 10040 22498
rect 9988 22434 10040 22440
rect 10000 21886 10028 22434
rect 9988 21880 10040 21886
rect 9988 21822 10040 21828
rect 10264 20656 10316 20662
rect 10264 20598 10316 20604
rect 9988 19704 10040 19710
rect 9988 19646 10040 19652
rect 10172 19704 10224 19710
rect 10172 19646 10224 19652
rect 10000 19302 10028 19646
rect 10184 19370 10212 19646
rect 10172 19364 10224 19370
rect 10172 19306 10224 19312
rect 9988 19296 10040 19302
rect 9988 19238 10040 19244
rect 10276 19098 10304 20598
rect 10356 19908 10408 19914
rect 10356 19850 10408 19856
rect 10368 19778 10396 19850
rect 10356 19772 10408 19778
rect 10356 19714 10408 19720
rect 10368 19574 10396 19714
rect 10356 19568 10408 19574
rect 10356 19510 10408 19516
rect 10264 19092 10316 19098
rect 10264 19034 10316 19040
rect 10356 19024 10408 19030
rect 10356 18966 10408 18972
rect 10368 18622 10396 18966
rect 10356 18616 10408 18622
rect 10356 18558 10408 18564
rect 9252 13040 9304 13046
rect 9252 12982 9304 12988
rect 9896 13040 9948 13046
rect 9896 12982 9948 12988
rect 8792 11952 8844 11958
rect 8792 11894 8844 11900
rect 8804 10122 8832 11894
rect 9160 11680 9212 11686
rect 9160 11622 9212 11628
rect 9068 11612 9120 11618
rect 8988 11572 9068 11600
rect 8884 11476 8936 11482
rect 8884 11418 8936 11424
rect 8896 11210 8924 11418
rect 8884 11204 8936 11210
rect 8884 11146 8936 11152
rect 8988 10326 9016 11572
rect 9068 11554 9120 11560
rect 9172 11210 9200 11622
rect 9160 11204 9212 11210
rect 9160 11146 9212 11152
rect 8976 10320 9028 10326
rect 8976 10262 9028 10268
rect 8792 10116 8844 10122
rect 8792 10058 8844 10064
rect 8792 9980 8844 9986
rect 8792 9922 8844 9928
rect 8804 9578 8832 9922
rect 8792 9572 8844 9578
rect 8792 9514 8844 9520
rect 8606 9472 8662 9481
rect 8606 9407 8662 9416
rect 8424 8892 8476 8898
rect 8424 8834 8476 8840
rect 7872 8348 7924 8354
rect 7872 8290 7924 8296
rect 8620 8218 8648 9407
rect 8700 8960 8752 8966
rect 8700 8902 8752 8908
rect 8608 8212 8660 8218
rect 8608 8154 8660 8160
rect 8620 7810 8648 8154
rect 8608 7804 8660 7810
rect 8608 7746 8660 7752
rect 7780 7668 7832 7674
rect 7780 7610 7832 7616
rect 8620 7334 8648 7746
rect 8608 7328 8660 7334
rect 8608 7270 8660 7276
rect 8148 7056 8200 7062
rect 8148 6998 8200 7004
rect 8160 6722 8188 6998
rect 8148 6716 8200 6722
rect 8148 6658 8200 6664
rect 8160 5158 8188 6658
rect 8712 6654 8740 8902
rect 8804 8354 8832 9514
rect 8792 8348 8844 8354
rect 8844 8308 8924 8336
rect 8792 8290 8844 8296
rect 8792 7668 8844 7674
rect 8792 7610 8844 7616
rect 8700 6648 8752 6654
rect 8700 6590 8752 6596
rect 8712 6314 8740 6590
rect 8700 6308 8752 6314
rect 8700 6250 8752 6256
rect 8424 6104 8476 6110
rect 8424 6046 8476 6052
rect 8436 5702 8464 6046
rect 8424 5696 8476 5702
rect 8424 5638 8476 5644
rect 8148 5152 8200 5158
rect 8148 5094 8200 5100
rect 8160 4682 8188 5094
rect 8148 4676 8200 4682
rect 8148 4618 8200 4624
rect 8804 4554 8832 7610
rect 8896 7402 8924 8308
rect 8884 7396 8936 7402
rect 8884 7338 8936 7344
rect 8882 7296 8938 7305
rect 8882 7231 8938 7240
rect 8896 6858 8924 7231
rect 8884 6852 8936 6858
rect 8884 6794 8936 6800
rect 8712 4526 8832 4554
rect 7596 4064 7648 4070
rect 7596 4006 7648 4012
rect 7608 3594 7636 4006
rect 7596 3588 7648 3594
rect 7596 3530 7648 3536
rect 8148 3316 8200 3322
rect 8148 3258 8200 3264
rect 6032 3248 6084 3254
rect 6032 3190 6084 3196
rect 7504 3248 7556 3254
rect 7504 3190 7556 3196
rect 6044 2438 6072 3190
rect 7516 2982 7544 3190
rect 8160 3050 8188 3258
rect 8148 3044 8200 3050
rect 8148 2986 8200 2992
rect 7504 2976 7556 2982
rect 7504 2918 7556 2924
rect 6860 2908 6912 2914
rect 6860 2850 6912 2856
rect 6124 2840 6176 2846
rect 6124 2782 6176 2788
rect 6136 2506 6164 2782
rect 6872 2506 6900 2850
rect 6124 2500 6176 2506
rect 6124 2442 6176 2448
rect 6860 2500 6912 2506
rect 6860 2442 6912 2448
rect 6032 2432 6084 2438
rect 6032 2374 6084 2380
rect 8160 2302 8188 2986
rect 6768 2296 6820 2302
rect 6768 2238 6820 2244
rect 8056 2296 8108 2302
rect 8056 2238 8108 2244
rect 8148 2296 8200 2302
rect 8148 2238 8200 2244
rect 4652 1888 4704 1894
rect 4652 1830 4704 1836
rect 5848 1888 5900 1894
rect 5848 1830 5900 1836
rect 4560 1752 4612 1758
rect 4560 1694 4612 1700
rect 3916 1412 3968 1418
rect 3916 1354 3968 1360
rect 4572 1282 4600 1694
rect 4664 1418 4692 1830
rect 4652 1412 4704 1418
rect 4652 1354 4704 1360
rect 5860 1350 5888 1830
rect 6780 1826 6808 2238
rect 7228 2160 7280 2166
rect 7228 2102 7280 2108
rect 6768 1820 6820 1826
rect 6768 1762 6820 1768
rect 5848 1344 5900 1350
rect 5848 1286 5900 1292
rect 6780 1282 6808 1762
rect 6952 1752 7004 1758
rect 6952 1694 7004 1700
rect 6964 1418 6992 1694
rect 6952 1412 7004 1418
rect 6952 1354 7004 1360
rect 4560 1276 4612 1282
rect 4560 1218 4612 1224
rect 6768 1276 6820 1282
rect 6768 1218 6820 1224
rect 4468 1140 4520 1146
rect 4468 1082 4520 1088
rect 2168 1072 2220 1078
rect 2168 1014 2220 1020
rect 3180 1072 3232 1078
rect 3180 1014 3232 1020
rect 3192 424 3220 1014
rect 3504 428 3824 448
rect 3504 426 3516 428
rect 3572 426 3596 428
rect 3652 426 3676 428
rect 3732 426 3756 428
rect 3812 426 3824 428
rect 390 0 502 424
rect 1678 0 1790 424
rect 3150 0 3262 424
rect 3504 374 3510 426
rect 3572 374 3574 426
rect 3754 374 3756 426
rect 3818 374 3824 426
rect 4480 424 4508 1082
rect 5938 768 5994 777
rect 5938 703 5994 712
rect 5952 424 5980 703
rect 7240 424 7268 2102
rect 8068 1962 8096 2238
rect 8056 1956 8108 1962
rect 8056 1898 8108 1904
rect 8712 424 8740 4526
rect 8988 4410 9016 10262
rect 9160 6308 9212 6314
rect 9160 6250 9212 6256
rect 9172 5430 9200 6250
rect 9264 5566 9292 12982
rect 9894 12736 9950 12745
rect 9894 12671 9950 12680
rect 9908 12638 9936 12671
rect 9896 12632 9948 12638
rect 9896 12574 9948 12580
rect 9804 12156 9856 12162
rect 9804 12098 9856 12104
rect 9528 11544 9580 11550
rect 9712 11544 9764 11550
rect 9580 11504 9660 11532
rect 9528 11486 9580 11492
rect 9528 10116 9580 10122
rect 9528 10058 9580 10064
rect 9540 9850 9568 10058
rect 9344 9844 9396 9850
rect 9344 9786 9396 9792
rect 9528 9844 9580 9850
rect 9528 9786 9580 9792
rect 9356 9510 9384 9786
rect 9344 9504 9396 9510
rect 9344 9446 9396 9452
rect 9356 9034 9384 9446
rect 9632 9374 9660 11504
rect 9712 11486 9764 11492
rect 9724 11385 9752 11486
rect 9816 11482 9844 12098
rect 9908 11754 9936 12574
rect 9986 12056 10042 12065
rect 9986 11991 10042 12000
rect 9896 11748 9948 11754
rect 9896 11690 9948 11696
rect 10000 11618 10028 11991
rect 9988 11612 10040 11618
rect 9988 11554 10040 11560
rect 9804 11476 9856 11482
rect 9804 11418 9856 11424
rect 9710 11376 9766 11385
rect 9710 11311 9766 11320
rect 9724 11142 9752 11311
rect 9712 11136 9764 11142
rect 9712 11078 9764 11084
rect 10000 11074 10028 11554
rect 9988 11068 10040 11074
rect 9988 11010 10040 11016
rect 10170 10968 10226 10977
rect 10170 10903 10226 10912
rect 10184 10870 10212 10903
rect 10172 10864 10224 10870
rect 10172 10806 10224 10812
rect 10264 10864 10316 10870
rect 10264 10806 10316 10812
rect 9988 9436 10040 9442
rect 9988 9378 10040 9384
rect 9436 9368 9488 9374
rect 9436 9310 9488 9316
rect 9620 9368 9672 9374
rect 9620 9310 9672 9316
rect 9344 9028 9396 9034
rect 9344 8970 9396 8976
rect 9448 8694 9476 9310
rect 9712 9300 9764 9306
rect 9712 9242 9764 9248
rect 9724 8898 9752 9242
rect 10000 8898 10028 9378
rect 9712 8892 9764 8898
rect 9712 8834 9764 8840
rect 9988 8892 10040 8898
rect 9988 8834 10040 8840
rect 9436 8688 9488 8694
rect 9436 8630 9488 8636
rect 9252 5560 9304 5566
rect 9252 5502 9304 5508
rect 9160 5424 9212 5430
rect 9160 5366 9212 5372
rect 9160 5016 9212 5022
rect 9160 4958 9212 4964
rect 9172 4682 9200 4958
rect 9160 4676 9212 4682
rect 9160 4618 9212 4624
rect 8976 4404 9028 4410
rect 8976 4346 9028 4352
rect 9172 3866 9200 4618
rect 9448 4138 9476 8630
rect 10000 8422 10028 8834
rect 9988 8416 10040 8422
rect 9988 8358 10040 8364
rect 9528 6172 9580 6178
rect 9528 6114 9580 6120
rect 9540 5498 9568 6114
rect 9712 5628 9764 5634
rect 9712 5570 9764 5576
rect 9528 5492 9580 5498
rect 9528 5434 9580 5440
rect 9540 5226 9568 5434
rect 9724 5226 9752 5570
rect 10080 5560 10132 5566
rect 10080 5502 10132 5508
rect 9528 5220 9580 5226
rect 9528 5162 9580 5168
rect 9712 5220 9764 5226
rect 9712 5162 9764 5168
rect 9724 4682 9752 5162
rect 9804 5084 9856 5090
rect 9804 5026 9856 5032
rect 9712 4676 9764 4682
rect 9712 4618 9764 4624
rect 9816 4614 9844 5026
rect 10092 4886 10120 5502
rect 10080 4880 10132 4886
rect 10080 4822 10132 4828
rect 9804 4608 9856 4614
rect 9804 4550 9856 4556
rect 10092 4426 10120 4822
rect 9908 4398 10120 4426
rect 10172 4472 10224 4478
rect 10172 4414 10224 4420
rect 9436 4132 9488 4138
rect 9436 4074 9488 4080
rect 9160 3860 9212 3866
rect 9160 3802 9212 3808
rect 9908 3458 9936 4398
rect 10184 3866 10212 4414
rect 10172 3860 10224 3866
rect 10172 3802 10224 3808
rect 10184 3458 10212 3802
rect 9896 3452 9948 3458
rect 9896 3394 9948 3400
rect 10172 3452 10224 3458
rect 10172 3394 10224 3400
rect 9252 3248 9304 3254
rect 9252 3190 9304 3196
rect 9264 2370 9292 3190
rect 9712 2840 9764 2846
rect 9712 2782 9764 2788
rect 9988 2840 10040 2846
rect 9988 2782 10040 2788
rect 9252 2364 9304 2370
rect 9252 2306 9304 2312
rect 9724 1962 9752 2782
rect 10000 2506 10028 2782
rect 9988 2500 10040 2506
rect 9988 2442 10040 2448
rect 9804 2228 9856 2234
rect 9804 2170 9856 2176
rect 9712 1956 9764 1962
rect 9712 1898 9764 1904
rect 9816 1418 9844 2170
rect 10080 1752 10132 1758
rect 10080 1694 10132 1700
rect 10092 1418 10120 1694
rect 9804 1412 9856 1418
rect 9804 1354 9856 1360
rect 10080 1412 10132 1418
rect 10080 1354 10132 1360
rect 10276 618 10304 10806
rect 10356 9436 10408 9442
rect 10356 9378 10408 9384
rect 10368 8966 10396 9378
rect 10356 8960 10408 8966
rect 10356 8902 10408 8908
rect 10356 7804 10408 7810
rect 10356 7746 10408 7752
rect 10368 6246 10396 7746
rect 10356 6240 10408 6246
rect 10356 6182 10408 6188
rect 10460 5684 10488 23846
rect 10540 20792 10592 20798
rect 10540 20734 10592 20740
rect 10552 19234 10580 20734
rect 10540 19228 10592 19234
rect 10540 19170 10592 19176
rect 10552 18826 10580 19170
rect 10540 18820 10592 18826
rect 10540 18762 10592 18768
rect 10540 16304 10592 16310
rect 10540 16246 10592 16252
rect 10552 12298 10580 16246
rect 10540 12292 10592 12298
rect 10540 12234 10592 12240
rect 10540 5696 10592 5702
rect 10460 5656 10540 5684
rect 10356 5560 10408 5566
rect 10356 5502 10408 5508
rect 10368 3390 10396 5502
rect 10460 4682 10488 5656
rect 10540 5638 10592 5644
rect 10448 4676 10500 4682
rect 10448 4618 10500 4624
rect 10540 4608 10592 4614
rect 10540 4550 10592 4556
rect 10552 3390 10580 4550
rect 10644 3866 10672 25562
rect 10736 22566 10764 26106
rect 11460 25008 11512 25014
rect 11460 24950 11512 24956
rect 11276 24056 11328 24062
rect 11276 23998 11328 24004
rect 11092 23580 11144 23586
rect 11092 23522 11144 23528
rect 11184 23580 11236 23586
rect 11184 23522 11236 23528
rect 10908 23512 10960 23518
rect 10908 23454 10960 23460
rect 10920 22838 10948 23454
rect 11104 23042 11132 23522
rect 11092 23036 11144 23042
rect 11092 22978 11144 22984
rect 10908 22832 10960 22838
rect 10960 22792 11040 22820
rect 10908 22774 10960 22780
rect 10724 22560 10776 22566
rect 10776 22520 10856 22548
rect 10724 22502 10776 22508
rect 10724 22424 10776 22430
rect 10724 22366 10776 22372
rect 10736 21818 10764 22366
rect 10828 22090 10856 22520
rect 10908 22424 10960 22430
rect 10908 22366 10960 22372
rect 10816 22084 10868 22090
rect 10816 22026 10868 22032
rect 10920 22022 10948 22366
rect 10908 22016 10960 22022
rect 10908 21958 10960 21964
rect 11012 21954 11040 22792
rect 11000 21948 11052 21954
rect 11000 21890 11052 21896
rect 10724 21812 10776 21818
rect 10724 21754 10776 21760
rect 10736 21342 10764 21754
rect 10908 21404 10960 21410
rect 10908 21346 10960 21352
rect 10724 21336 10776 21342
rect 10724 21278 10776 21284
rect 10816 21336 10868 21342
rect 10816 21278 10868 21284
rect 10736 21002 10764 21278
rect 10724 20996 10776 21002
rect 10724 20938 10776 20944
rect 10828 20662 10856 21278
rect 10920 20730 10948 21346
rect 10908 20724 10960 20730
rect 10908 20666 10960 20672
rect 10816 20656 10868 20662
rect 10816 20598 10868 20604
rect 11012 20236 11040 21890
rect 11104 21410 11132 22978
rect 11196 22838 11224 23522
rect 11184 22832 11236 22838
rect 11184 22774 11236 22780
rect 11092 21404 11144 21410
rect 11092 21346 11144 21352
rect 11104 21002 11132 21346
rect 11196 21274 11224 22774
rect 11184 21268 11236 21274
rect 11184 21210 11236 21216
rect 11092 20996 11144 21002
rect 11092 20938 11144 20944
rect 11196 20662 11224 21210
rect 11184 20656 11236 20662
rect 11184 20598 11236 20604
rect 11196 20322 11224 20598
rect 11184 20316 11236 20322
rect 11184 20258 11236 20264
rect 11092 20248 11144 20254
rect 11012 20208 11092 20236
rect 11092 20190 11144 20196
rect 11104 19710 11132 20190
rect 11196 19846 11224 20258
rect 11184 19840 11236 19846
rect 11184 19782 11236 19788
rect 11092 19704 11144 19710
rect 11092 19646 11144 19652
rect 11288 18826 11316 23998
rect 11472 23518 11500 24950
rect 11920 24056 11972 24062
rect 11920 23998 11972 24004
rect 11460 23512 11512 23518
rect 11460 23454 11512 23460
rect 11472 23110 11500 23454
rect 11460 23104 11512 23110
rect 11460 23046 11512 23052
rect 11932 23042 11960 23998
rect 12012 23988 12064 23994
rect 12012 23930 12064 23936
rect 12104 23988 12156 23994
rect 12104 23930 12156 23936
rect 12024 23897 12052 23930
rect 12010 23888 12066 23897
rect 12010 23823 12066 23832
rect 12116 23450 12144 23930
rect 12104 23444 12156 23450
rect 12104 23386 12156 23392
rect 12116 23178 12144 23386
rect 12104 23172 12156 23178
rect 12104 23114 12156 23120
rect 11920 23036 11972 23042
rect 11920 22978 11972 22984
rect 11920 22832 11972 22838
rect 11920 22774 11972 22780
rect 11552 22424 11604 22430
rect 11552 22366 11604 22372
rect 11460 22016 11512 22022
rect 11460 21958 11512 21964
rect 11472 21410 11500 21958
rect 11460 21404 11512 21410
rect 11460 21346 11512 21352
rect 11368 20996 11420 21002
rect 11368 20938 11420 20944
rect 11380 20186 11408 20938
rect 11472 20798 11500 21346
rect 11460 20792 11512 20798
rect 11460 20734 11512 20740
rect 11368 20180 11420 20186
rect 11368 20122 11420 20128
rect 11564 19234 11592 22366
rect 11828 21336 11880 21342
rect 11828 21278 11880 21284
rect 11644 20656 11696 20662
rect 11644 20598 11696 20604
rect 11656 20322 11684 20598
rect 11644 20316 11696 20322
rect 11644 20258 11696 20264
rect 11656 19370 11684 20258
rect 11840 20254 11868 21278
rect 11736 20248 11788 20254
rect 11736 20190 11788 20196
rect 11828 20248 11880 20254
rect 11828 20190 11880 20196
rect 11748 19710 11776 20190
rect 11736 19704 11788 19710
rect 11736 19646 11788 19652
rect 11748 19370 11776 19646
rect 11644 19364 11696 19370
rect 11644 19306 11696 19312
rect 11736 19364 11788 19370
rect 11736 19306 11788 19312
rect 11552 19228 11604 19234
rect 11552 19170 11604 19176
rect 11564 18826 11592 19170
rect 11736 19160 11788 19166
rect 11736 19102 11788 19108
rect 11276 18820 11328 18826
rect 11276 18762 11328 18768
rect 11552 18820 11604 18826
rect 11552 18762 11604 18768
rect 11288 18690 11316 18762
rect 11276 18684 11328 18690
rect 11276 18626 11328 18632
rect 11288 17058 11316 18626
rect 11564 17738 11592 18762
rect 11552 17732 11604 17738
rect 11552 17674 11604 17680
rect 11276 17052 11328 17058
rect 11276 16994 11328 17000
rect 11748 16582 11776 19102
rect 11932 17670 11960 22774
rect 12196 21880 12248 21886
rect 12196 21822 12248 21828
rect 12012 21812 12064 21818
rect 12012 21754 12064 21760
rect 12024 20186 12052 21754
rect 12208 20186 12236 21822
rect 12012 20180 12064 20186
rect 12012 20122 12064 20128
rect 12196 20180 12248 20186
rect 12196 20122 12248 20128
rect 12024 19914 12052 20122
rect 12104 20112 12156 20118
rect 12104 20054 12156 20060
rect 12012 19908 12064 19914
rect 12012 19850 12064 19856
rect 12116 19710 12144 20054
rect 12300 19914 12328 27126
rect 12380 23376 12432 23382
rect 12380 23318 12432 23324
rect 12392 23178 12420 23318
rect 12380 23172 12432 23178
rect 12380 23114 12432 23120
rect 12288 19908 12340 19914
rect 12288 19850 12340 19856
rect 12104 19704 12156 19710
rect 12104 19646 12156 19652
rect 12116 19302 12144 19646
rect 12300 19370 12328 19850
rect 12392 19710 12420 23114
rect 12380 19704 12432 19710
rect 12380 19646 12432 19652
rect 12288 19364 12340 19370
rect 12288 19306 12340 19312
rect 12104 19296 12156 19302
rect 12104 19238 12156 19244
rect 12116 18826 12144 19238
rect 12104 18820 12156 18826
rect 12104 18762 12156 18768
rect 12116 18622 12144 18762
rect 12104 18616 12156 18622
rect 12104 18558 12156 18564
rect 11920 17664 11972 17670
rect 11920 17606 11972 17612
rect 11736 16576 11788 16582
rect 11736 16518 11788 16524
rect 11748 16446 11776 16518
rect 11736 16440 11788 16446
rect 11736 16382 11788 16388
rect 10724 15964 10776 15970
rect 10724 15906 10776 15912
rect 11000 15964 11052 15970
rect 11000 15906 11052 15912
rect 10736 15562 10764 15906
rect 11012 15766 11040 15906
rect 11000 15760 11052 15766
rect 11000 15702 11052 15708
rect 11012 15562 11040 15702
rect 10724 15556 10776 15562
rect 10724 15498 10776 15504
rect 11000 15556 11052 15562
rect 11000 15498 11052 15504
rect 10736 14950 10764 15498
rect 11748 15494 11776 16382
rect 12104 16372 12156 16378
rect 12104 16314 12156 16320
rect 12116 15970 12144 16314
rect 12104 15964 12156 15970
rect 12104 15906 12156 15912
rect 12116 15562 12144 15906
rect 12288 15896 12340 15902
rect 12288 15838 12340 15844
rect 12104 15556 12156 15562
rect 12104 15498 12156 15504
rect 11736 15488 11788 15494
rect 11736 15430 11788 15436
rect 11920 15488 11972 15494
rect 11920 15430 11972 15436
rect 10724 14944 10776 14950
rect 10724 14886 10776 14892
rect 11184 14944 11236 14950
rect 11184 14886 11236 14892
rect 11092 14808 11144 14814
rect 11092 14750 11144 14756
rect 10724 14740 10776 14746
rect 10724 14682 10776 14688
rect 10736 6110 10764 14682
rect 11104 14474 11132 14750
rect 11196 14474 11224 14886
rect 11748 14882 11776 15430
rect 11932 15358 11960 15430
rect 11920 15352 11972 15358
rect 11920 15294 11972 15300
rect 11736 14876 11788 14882
rect 11736 14818 11788 14824
rect 11748 14474 11776 14818
rect 12116 14474 12144 15498
rect 11092 14468 11144 14474
rect 11092 14410 11144 14416
rect 11184 14468 11236 14474
rect 11184 14410 11236 14416
rect 11736 14468 11788 14474
rect 11736 14410 11788 14416
rect 12104 14468 12156 14474
rect 12104 14410 12156 14416
rect 11196 14270 11224 14410
rect 12116 14270 12144 14410
rect 11184 14264 11236 14270
rect 11184 14206 11236 14212
rect 12104 14264 12156 14270
rect 12104 14206 12156 14212
rect 11828 14128 11880 14134
rect 11828 14070 11880 14076
rect 11840 13862 11868 14070
rect 11828 13856 11880 13862
rect 11828 13798 11880 13804
rect 12300 13318 12328 15838
rect 12380 13652 12432 13658
rect 12380 13594 12432 13600
rect 12288 13312 12340 13318
rect 12288 13254 12340 13260
rect 10816 13108 10868 13114
rect 10816 13050 10868 13056
rect 10828 12638 10856 13050
rect 11460 13040 11512 13046
rect 11460 12982 11512 12988
rect 11472 12774 11500 12982
rect 12300 12774 12328 13254
rect 12392 13182 12420 13594
rect 12380 13176 12432 13182
rect 12380 13118 12432 13124
rect 12392 12774 12420 13118
rect 11460 12768 11512 12774
rect 11460 12710 11512 12716
rect 12288 12768 12340 12774
rect 12288 12710 12340 12716
rect 12380 12768 12432 12774
rect 12380 12710 12432 12716
rect 11276 12700 11328 12706
rect 11276 12642 11328 12648
rect 10816 12632 10868 12638
rect 10816 12574 10868 12580
rect 10828 12298 10856 12574
rect 10816 12292 10868 12298
rect 10816 12234 10868 12240
rect 11288 12162 11316 12642
rect 11472 12230 11500 12710
rect 11460 12224 11512 12230
rect 11460 12166 11512 12172
rect 11276 12156 11328 12162
rect 11276 12098 11328 12104
rect 10814 10152 10870 10161
rect 10814 10087 10870 10096
rect 10828 9850 10856 10087
rect 10816 9844 10868 9850
rect 10816 9786 10868 9792
rect 10828 9374 10856 9786
rect 11552 9776 11604 9782
rect 11552 9718 11604 9724
rect 10816 9368 10868 9374
rect 10816 9310 10868 9316
rect 11184 8756 11236 8762
rect 11184 8698 11236 8704
rect 11196 8354 11224 8698
rect 11460 8688 11512 8694
rect 11460 8630 11512 8636
rect 10816 8348 10868 8354
rect 10816 8290 10868 8296
rect 11184 8348 11236 8354
rect 11184 8290 11236 8296
rect 10828 7878 10856 8290
rect 11196 7946 11224 8290
rect 11472 8286 11500 8630
rect 11564 8422 11592 9718
rect 12300 9578 12328 12710
rect 12392 12298 12420 12710
rect 12484 12706 12512 29366
rect 13116 29360 13168 29366
rect 13116 29302 13168 29308
rect 13208 29360 13260 29366
rect 13208 29302 13260 29308
rect 13128 28414 13156 29302
rect 13220 28482 13248 29302
rect 13312 29094 13340 29370
rect 13300 29088 13352 29094
rect 13300 29030 13352 29036
rect 13300 28952 13352 28958
rect 13300 28894 13352 28900
rect 13312 28618 13340 28894
rect 13300 28612 13352 28618
rect 13300 28554 13352 28560
rect 13208 28476 13260 28482
rect 13208 28418 13260 28424
rect 13116 28408 13168 28414
rect 13116 28350 13168 28356
rect 12656 27864 12708 27870
rect 12656 27806 12708 27812
rect 12668 27394 12696 27806
rect 12656 27388 12708 27394
rect 12656 27330 12708 27336
rect 12564 27320 12616 27326
rect 12564 27262 12616 27268
rect 12576 26986 12604 27262
rect 12564 26980 12616 26986
rect 12564 26922 12616 26928
rect 12576 25354 12604 26922
rect 12748 25688 12800 25694
rect 12748 25630 12800 25636
rect 12564 25348 12616 25354
rect 12564 25290 12616 25296
rect 12576 24266 12604 25290
rect 12656 25008 12708 25014
rect 12656 24950 12708 24956
rect 12564 24260 12616 24266
rect 12564 24202 12616 24208
rect 12668 23926 12696 24950
rect 12564 23920 12616 23926
rect 12562 23888 12564 23897
rect 12656 23920 12708 23926
rect 12616 23888 12618 23897
rect 12656 23862 12708 23868
rect 12562 23823 12618 23832
rect 12668 22974 12696 23862
rect 12656 22968 12708 22974
rect 12656 22910 12708 22916
rect 12656 22288 12708 22294
rect 12656 22230 12708 22236
rect 12668 21750 12696 22230
rect 12656 21744 12708 21750
rect 12656 21686 12708 21692
rect 12668 20866 12696 21686
rect 12656 20860 12708 20866
rect 12656 20802 12708 20808
rect 12760 19302 12788 25630
rect 13024 25552 13076 25558
rect 13024 25494 13076 25500
rect 12840 23444 12892 23450
rect 12840 23386 12892 23392
rect 12852 22974 12880 23386
rect 12840 22968 12892 22974
rect 12840 22910 12892 22916
rect 13036 22838 13064 25494
rect 13300 25008 13352 25014
rect 13300 24950 13352 24956
rect 13312 24713 13340 24950
rect 13298 24704 13354 24713
rect 13298 24639 13354 24648
rect 13208 24056 13260 24062
rect 13208 23998 13260 24004
rect 13220 23722 13248 23998
rect 13208 23716 13260 23722
rect 13208 23658 13260 23664
rect 13220 23178 13248 23658
rect 13208 23172 13260 23178
rect 13260 23132 13340 23160
rect 13208 23114 13260 23120
rect 13208 22968 13260 22974
rect 13208 22910 13260 22916
rect 13024 22832 13076 22838
rect 13024 22774 13076 22780
rect 13220 22634 13248 22910
rect 13208 22628 13260 22634
rect 13208 22570 13260 22576
rect 13024 22492 13076 22498
rect 13024 22434 13076 22440
rect 13036 21750 13064 22434
rect 13312 21954 13340 23132
rect 13300 21948 13352 21954
rect 13300 21890 13352 21896
rect 13024 21744 13076 21750
rect 13024 21686 13076 21692
rect 12840 21404 12892 21410
rect 12840 21346 12892 21352
rect 12852 21002 12880 21346
rect 13036 21342 13064 21686
rect 13312 21546 13340 21890
rect 13300 21540 13352 21546
rect 13300 21482 13352 21488
rect 13024 21336 13076 21342
rect 13024 21278 13076 21284
rect 13036 21002 13064 21278
rect 12840 20996 12892 21002
rect 12840 20938 12892 20944
rect 13024 20996 13076 21002
rect 13024 20938 13076 20944
rect 12840 19704 12892 19710
rect 12840 19646 12892 19652
rect 12748 19296 12800 19302
rect 12748 19238 12800 19244
rect 12760 18826 12788 19238
rect 12852 19234 12880 19646
rect 12932 19636 12984 19642
rect 12932 19578 12984 19584
rect 12840 19228 12892 19234
rect 12840 19170 12892 19176
rect 12748 18820 12800 18826
rect 12748 18762 12800 18768
rect 12760 18146 12788 18762
rect 12852 18690 12880 19170
rect 12840 18684 12892 18690
rect 12840 18626 12892 18632
rect 12944 18146 12972 19578
rect 13116 18616 13168 18622
rect 13116 18558 13168 18564
rect 13128 18146 13156 18558
rect 12748 18140 12800 18146
rect 12748 18082 12800 18088
rect 12932 18140 12984 18146
rect 12932 18082 12984 18088
rect 13116 18140 13168 18146
rect 13116 18082 13168 18088
rect 12760 17738 12788 18082
rect 12748 17732 12800 17738
rect 12748 17674 12800 17680
rect 12760 17534 12788 17674
rect 12944 17670 12972 18082
rect 13024 17732 13076 17738
rect 13128 17720 13156 18082
rect 13076 17692 13156 17720
rect 13024 17674 13076 17680
rect 12932 17664 12984 17670
rect 12932 17606 12984 17612
rect 12748 17528 12800 17534
rect 12748 17470 12800 17476
rect 12760 17126 12788 17470
rect 12748 17120 12800 17126
rect 12748 17062 12800 17068
rect 12944 17058 12972 17606
rect 12932 17052 12984 17058
rect 12932 16994 12984 17000
rect 12564 16440 12616 16446
rect 12564 16382 12616 16388
rect 12576 16038 12604 16382
rect 12564 16032 12616 16038
rect 12564 15974 12616 15980
rect 12576 15018 12604 15974
rect 13116 15284 13168 15290
rect 13116 15226 13168 15232
rect 12564 15012 12616 15018
rect 12564 14954 12616 14960
rect 13128 13794 13156 15226
rect 13404 14214 13432 30594
rect 13680 30250 13708 31664
rect 14968 30250 14996 31664
rect 13668 30244 13720 30250
rect 13668 30186 13720 30192
rect 14864 30244 14916 30250
rect 14864 30186 14916 30192
rect 14956 30244 15008 30250
rect 14956 30186 15008 30192
rect 13666 29736 13722 29745
rect 13666 29671 13722 29680
rect 13680 29570 13708 29671
rect 13668 29564 13720 29570
rect 13668 29506 13720 29512
rect 13680 29026 13708 29506
rect 13668 29020 13720 29026
rect 13668 28962 13720 28968
rect 13680 28618 13708 28962
rect 14588 28952 14640 28958
rect 14588 28894 14640 28900
rect 14680 28952 14732 28958
rect 14680 28894 14732 28900
rect 14600 28618 14628 28894
rect 13668 28612 13720 28618
rect 13668 28554 13720 28560
rect 14588 28612 14640 28618
rect 14588 28554 14640 28560
rect 14692 28278 14720 28894
rect 14680 28272 14732 28278
rect 14680 28214 14732 28220
rect 14692 26306 14720 28214
rect 14876 27802 14904 30186
rect 16440 30130 16468 31664
rect 16888 30516 16940 30522
rect 16888 30458 16940 30464
rect 16900 30182 16928 30458
rect 16888 30176 16940 30182
rect 16440 30102 16560 30130
rect 16888 30118 16940 30124
rect 16152 30040 16204 30046
rect 16152 29982 16204 29988
rect 16428 30040 16480 30046
rect 16428 29982 16480 29988
rect 15508 29564 15560 29570
rect 15508 29506 15560 29512
rect 15048 29428 15100 29434
rect 15048 29370 15100 29376
rect 15416 29428 15468 29434
rect 15416 29370 15468 29376
rect 15060 28890 15088 29370
rect 15232 29088 15284 29094
rect 15232 29030 15284 29036
rect 15048 28884 15100 28890
rect 15048 28826 15100 28832
rect 15060 28414 15088 28826
rect 15048 28408 15100 28414
rect 15048 28350 15100 28356
rect 14956 28000 15008 28006
rect 14956 27942 15008 27948
rect 14864 27796 14916 27802
rect 14864 27738 14916 27744
rect 14968 27462 14996 27942
rect 15060 27462 15088 28350
rect 15244 28278 15272 29030
rect 15324 29020 15376 29026
rect 15428 29008 15456 29370
rect 15520 29026 15548 29506
rect 15968 29496 16020 29502
rect 15968 29438 16020 29444
rect 15376 28980 15456 29008
rect 15324 28962 15376 28968
rect 15428 28618 15456 28980
rect 15508 29020 15560 29026
rect 15508 28962 15560 28968
rect 15416 28612 15468 28618
rect 15416 28554 15468 28560
rect 15980 28346 16008 29438
rect 16164 29366 16192 29982
rect 16244 29904 16296 29910
rect 16244 29846 16296 29852
rect 16256 29706 16284 29846
rect 16440 29706 16468 29982
rect 16244 29700 16296 29706
rect 16244 29642 16296 29648
rect 16428 29700 16480 29706
rect 16428 29642 16480 29648
rect 16532 29473 16560 30102
rect 16796 29496 16848 29502
rect 16518 29464 16574 29473
rect 16796 29438 16848 29444
rect 16518 29399 16574 29408
rect 16152 29360 16204 29366
rect 16152 29302 16204 29308
rect 16152 29020 16204 29026
rect 16152 28962 16204 28968
rect 16164 28482 16192 28962
rect 16152 28476 16204 28482
rect 16152 28418 16204 28424
rect 15416 28340 15468 28346
rect 15416 28282 15468 28288
rect 15968 28340 16020 28346
rect 15968 28282 16020 28288
rect 15232 28272 15284 28278
rect 15232 28214 15284 28220
rect 14956 27456 15008 27462
rect 14956 27398 15008 27404
rect 15048 27456 15100 27462
rect 15048 27398 15100 27404
rect 14968 27190 14996 27398
rect 14956 27184 15008 27190
rect 14956 27126 15008 27132
rect 14864 26844 14916 26850
rect 14864 26786 14916 26792
rect 14680 26300 14732 26306
rect 14680 26242 14732 26248
rect 14680 26096 14732 26102
rect 14680 26038 14732 26044
rect 14692 25898 14720 26038
rect 14876 25898 14904 26786
rect 15060 26730 15088 27398
rect 15244 27190 15272 28214
rect 15428 27734 15456 28282
rect 16164 28074 16192 28418
rect 16612 28272 16664 28278
rect 16612 28214 16664 28220
rect 16152 28068 16204 28074
rect 16152 28010 16204 28016
rect 15968 27932 16020 27938
rect 15968 27874 16020 27880
rect 15416 27728 15468 27734
rect 15416 27670 15468 27676
rect 15428 27530 15456 27670
rect 15980 27530 16008 27874
rect 16624 27734 16652 28214
rect 16808 27938 16836 29438
rect 16900 29162 16928 30118
rect 17728 30114 17756 31664
rect 19200 31626 19228 31664
rect 19200 31598 19320 31626
rect 18864 31436 19184 31456
rect 18864 31434 18876 31436
rect 18932 31434 18956 31436
rect 19012 31434 19036 31436
rect 19092 31434 19116 31436
rect 19172 31434 19184 31436
rect 18864 31382 18870 31434
rect 18932 31382 18934 31434
rect 19114 31382 19116 31434
rect 19178 31382 19184 31434
rect 18864 31380 18876 31382
rect 18932 31380 18956 31382
rect 19012 31380 19036 31382
rect 19092 31380 19116 31382
rect 19172 31380 19184 31382
rect 18864 31360 19184 31380
rect 19292 30658 19320 31598
rect 19280 30652 19332 30658
rect 19280 30594 19332 30600
rect 18360 30448 18412 30454
rect 18360 30390 18412 30396
rect 17716 30108 17768 30114
rect 17716 30050 17768 30056
rect 18268 30040 18320 30046
rect 18268 29982 18320 29988
rect 18280 29638 18308 29982
rect 18268 29632 18320 29638
rect 18268 29574 18320 29580
rect 17624 29564 17676 29570
rect 17624 29506 17676 29512
rect 17636 29434 17664 29506
rect 18280 29502 18308 29574
rect 17900 29496 17952 29502
rect 17900 29438 17952 29444
rect 18268 29496 18320 29502
rect 18268 29438 18320 29444
rect 17624 29428 17676 29434
rect 17624 29370 17676 29376
rect 17348 29360 17400 29366
rect 17348 29302 17400 29308
rect 16888 29156 16940 29162
rect 16888 29098 16940 29104
rect 16980 28884 17032 28890
rect 16980 28826 17032 28832
rect 17164 28884 17216 28890
rect 17164 28826 17216 28832
rect 16992 28618 17020 28826
rect 16980 28612 17032 28618
rect 16980 28554 17032 28560
rect 17176 28550 17204 28826
rect 17164 28544 17216 28550
rect 17164 28486 17216 28492
rect 16796 27932 16848 27938
rect 16796 27874 16848 27880
rect 16612 27728 16664 27734
rect 16612 27670 16664 27676
rect 15416 27524 15468 27530
rect 15416 27466 15468 27472
rect 15968 27524 16020 27530
rect 15968 27466 16020 27472
rect 16428 27524 16480 27530
rect 16428 27466 16480 27472
rect 15968 27252 16020 27258
rect 15968 27194 16020 27200
rect 15232 27184 15284 27190
rect 15232 27126 15284 27132
rect 15244 26850 15272 27126
rect 15232 26844 15284 26850
rect 15232 26786 15284 26792
rect 14968 26702 15088 26730
rect 15140 26708 15192 26714
rect 14968 26442 14996 26702
rect 15140 26650 15192 26656
rect 15048 26640 15100 26646
rect 15048 26582 15100 26588
rect 14956 26436 15008 26442
rect 14956 26378 15008 26384
rect 15060 26238 15088 26582
rect 15048 26232 15100 26238
rect 15048 26174 15100 26180
rect 14680 25892 14732 25898
rect 14680 25834 14732 25840
rect 14864 25892 14916 25898
rect 14864 25834 14916 25840
rect 14692 25558 14720 25834
rect 15060 25830 15088 26174
rect 15048 25824 15100 25830
rect 15048 25766 15100 25772
rect 15152 25762 15180 26650
rect 15244 26170 15272 26786
rect 15324 26776 15376 26782
rect 15324 26718 15376 26724
rect 15232 26164 15284 26170
rect 15232 26106 15284 26112
rect 15336 25898 15364 26718
rect 15508 26436 15560 26442
rect 15508 26378 15560 26384
rect 15520 26238 15548 26378
rect 15508 26232 15560 26238
rect 15508 26174 15560 26180
rect 15324 25892 15376 25898
rect 15324 25834 15376 25840
rect 15140 25756 15192 25762
rect 15140 25698 15192 25704
rect 14680 25552 14732 25558
rect 14680 25494 14732 25500
rect 14956 25280 15008 25286
rect 14956 25222 15008 25228
rect 14968 25014 14996 25222
rect 14956 25008 15008 25014
rect 14956 24950 15008 24956
rect 13944 24464 13996 24470
rect 13944 24406 13996 24412
rect 13956 24130 13984 24406
rect 13944 24124 13996 24130
rect 13944 24066 13996 24072
rect 13956 23994 13984 24066
rect 13944 23988 13996 23994
rect 13944 23930 13996 23936
rect 14968 23178 14996 24950
rect 14956 23172 15008 23178
rect 14956 23114 15008 23120
rect 14968 22906 14996 23114
rect 14956 22900 15008 22906
rect 14956 22842 15008 22848
rect 14772 22424 14824 22430
rect 14772 22366 14824 22372
rect 14784 21886 14812 22366
rect 14772 21880 14824 21886
rect 14772 21822 14824 21828
rect 14784 21546 14812 21822
rect 14772 21540 14824 21546
rect 14772 21482 14824 21488
rect 14968 20390 14996 22842
rect 15140 22492 15192 22498
rect 15140 22434 15192 22440
rect 15152 21750 15180 22434
rect 15140 21744 15192 21750
rect 15140 21686 15192 21692
rect 14956 20384 15008 20390
rect 14956 20326 15008 20332
rect 14680 20180 14732 20186
rect 14680 20122 14732 20128
rect 14692 19914 14720 20122
rect 14968 19914 14996 20326
rect 14680 19908 14732 19914
rect 14680 19850 14732 19856
rect 14956 19908 15008 19914
rect 14956 19850 15008 19856
rect 13484 19160 13536 19166
rect 13484 19102 13536 19108
rect 13496 18826 13524 19102
rect 13484 18820 13536 18826
rect 13484 18762 13536 18768
rect 14680 18752 14732 18758
rect 14680 18694 14732 18700
rect 13944 18684 13996 18690
rect 13944 18626 13996 18632
rect 13668 18548 13720 18554
rect 13668 18490 13720 18496
rect 13576 18072 13628 18078
rect 13576 18014 13628 18020
rect 13588 17194 13616 18014
rect 13680 17738 13708 18490
rect 13668 17732 13720 17738
rect 13668 17674 13720 17680
rect 13680 17534 13708 17674
rect 13668 17528 13720 17534
rect 13668 17470 13720 17476
rect 13760 17460 13812 17466
rect 13760 17402 13812 17408
rect 13576 17188 13628 17194
rect 13576 17130 13628 17136
rect 13772 16038 13800 17402
rect 13956 16514 13984 18626
rect 14588 18480 14640 18486
rect 14588 18422 14640 18428
rect 14600 18214 14628 18422
rect 14588 18208 14640 18214
rect 14588 18150 14640 18156
rect 14600 17670 14628 18150
rect 14588 17664 14640 17670
rect 14588 17606 14640 17612
rect 14600 17466 14628 17606
rect 14588 17460 14640 17466
rect 14588 17402 14640 17408
rect 14128 17392 14180 17398
rect 14128 17334 14180 17340
rect 14312 17392 14364 17398
rect 14312 17334 14364 17340
rect 14140 17194 14168 17334
rect 14128 17188 14180 17194
rect 14128 17130 14180 17136
rect 13944 16508 13996 16514
rect 13944 16450 13996 16456
rect 13760 16032 13812 16038
rect 13760 15974 13812 15980
rect 13404 14186 13524 14214
rect 12840 13788 12892 13794
rect 12840 13730 12892 13736
rect 13116 13788 13168 13794
rect 13116 13730 13168 13736
rect 12748 13584 12800 13590
rect 12748 13526 12800 13532
rect 12760 13182 12788 13526
rect 12852 13318 12880 13730
rect 13128 13386 13156 13730
rect 13392 13584 13444 13590
rect 13392 13526 13444 13532
rect 13404 13386 13432 13526
rect 13116 13380 13168 13386
rect 13116 13322 13168 13328
rect 13392 13380 13444 13386
rect 13392 13322 13444 13328
rect 12840 13312 12892 13318
rect 12840 13254 12892 13260
rect 12748 13176 12800 13182
rect 12748 13118 12800 13124
rect 12840 13176 12892 13182
rect 12840 13118 12892 13124
rect 12472 12700 12524 12706
rect 12472 12642 12524 12648
rect 12380 12292 12432 12298
rect 12380 12234 12432 12240
rect 12392 12094 12420 12234
rect 12380 12088 12432 12094
rect 12380 12030 12432 12036
rect 12564 11952 12616 11958
rect 12564 11894 12616 11900
rect 12576 11618 12604 11894
rect 12564 11612 12616 11618
rect 12564 11554 12616 11560
rect 12380 11544 12432 11550
rect 12380 11486 12432 11492
rect 12392 11142 12420 11486
rect 12576 11210 12604 11554
rect 12656 11476 12708 11482
rect 12656 11418 12708 11424
rect 12564 11204 12616 11210
rect 12564 11146 12616 11152
rect 12380 11136 12432 11142
rect 12380 11078 12432 11084
rect 12576 11074 12604 11146
rect 12668 11142 12696 11418
rect 12760 11414 12788 13118
rect 12852 12706 12880 13118
rect 12840 12700 12892 12706
rect 12840 12642 12892 12648
rect 13300 12632 13352 12638
rect 13300 12574 13352 12580
rect 13312 12298 13340 12574
rect 13300 12292 13352 12298
rect 13300 12234 13352 12240
rect 12748 11408 12800 11414
rect 12748 11350 12800 11356
rect 12656 11136 12708 11142
rect 12656 11078 12708 11084
rect 12564 11068 12616 11074
rect 12564 11010 12616 11016
rect 12576 10666 12604 11010
rect 12564 10660 12616 10666
rect 12564 10602 12616 10608
rect 12760 10530 12788 11350
rect 13116 11204 13168 11210
rect 13116 11146 13168 11152
rect 13128 10666 13156 11146
rect 13300 11000 13352 11006
rect 13300 10942 13352 10948
rect 13116 10660 13168 10666
rect 13116 10602 13168 10608
rect 12748 10524 12800 10530
rect 12748 10466 12800 10472
rect 13312 10394 13340 10942
rect 13300 10388 13352 10394
rect 13300 10330 13352 10336
rect 12746 9880 12802 9889
rect 12746 9815 12802 9824
rect 12288 9572 12340 9578
rect 12288 9514 12340 9520
rect 12010 9336 12066 9345
rect 12010 9271 12066 9280
rect 12024 9238 12052 9271
rect 12012 9232 12064 9238
rect 12012 9174 12064 9180
rect 12024 8898 12052 9174
rect 12012 8892 12064 8898
rect 12012 8834 12064 8840
rect 12300 8830 12328 9514
rect 12760 8966 12788 9815
rect 12748 8960 12800 8966
rect 12748 8902 12800 8908
rect 12656 8892 12708 8898
rect 12656 8834 12708 8840
rect 12288 8824 12340 8830
rect 12208 8784 12288 8812
rect 11552 8416 11604 8422
rect 11552 8358 11604 8364
rect 11460 8280 11512 8286
rect 11460 8222 11512 8228
rect 11184 7940 11236 7946
rect 11184 7882 11236 7888
rect 10816 7872 10868 7878
rect 10816 7814 10868 7820
rect 11472 7674 11500 8222
rect 11564 7810 11592 8358
rect 11552 7804 11604 7810
rect 11552 7746 11604 7752
rect 11460 7668 11512 7674
rect 11460 7610 11512 7616
rect 11552 7056 11604 7062
rect 11552 6998 11604 7004
rect 11564 6790 11592 6998
rect 11552 6784 11604 6790
rect 11552 6726 11604 6732
rect 11564 6586 11592 6726
rect 12208 6722 12236 8784
rect 12288 8766 12340 8772
rect 12668 8762 12696 8834
rect 12760 8830 12788 8902
rect 12748 8824 12800 8830
rect 12748 8766 12800 8772
rect 12656 8756 12708 8762
rect 12656 8698 12708 8704
rect 12668 8286 12696 8698
rect 12656 8280 12708 8286
rect 12656 8222 12708 8228
rect 12288 7736 12340 7742
rect 12288 7678 12340 7684
rect 12300 7266 12328 7678
rect 12288 7260 12340 7266
rect 12288 7202 12340 7208
rect 12300 6858 12328 7202
rect 12748 7056 12800 7062
rect 12748 6998 12800 7004
rect 13496 7010 13524 14186
rect 14220 14128 14272 14134
rect 14220 14070 14272 14076
rect 14232 13182 14260 14070
rect 14220 13176 14272 13182
rect 14220 13118 14272 13124
rect 14036 13040 14088 13046
rect 14036 12982 14088 12988
rect 14048 12162 14076 12982
rect 14232 12706 14260 13118
rect 14324 13114 14352 17334
rect 14692 16428 14720 18694
rect 14772 18140 14824 18146
rect 14772 18082 14824 18088
rect 14784 17738 14812 18082
rect 14772 17732 14824 17738
rect 14772 17674 14824 17680
rect 14968 17126 14996 19850
rect 15048 19160 15100 19166
rect 15048 19102 15100 19108
rect 15060 18826 15088 19102
rect 15048 18820 15100 18826
rect 15048 18762 15100 18768
rect 14956 17120 15008 17126
rect 14956 17062 15008 17068
rect 14772 16848 14824 16854
rect 14772 16790 14824 16796
rect 14600 16400 14720 16428
rect 14496 14808 14548 14814
rect 14496 14750 14548 14756
rect 14404 13720 14456 13726
rect 14404 13662 14456 13668
rect 14312 13108 14364 13114
rect 14312 13050 14364 13056
rect 14220 12700 14272 12706
rect 14220 12642 14272 12648
rect 14232 12230 14260 12642
rect 14220 12224 14272 12230
rect 14220 12166 14272 12172
rect 14036 12156 14088 12162
rect 14036 12098 14088 12104
rect 14036 12020 14088 12026
rect 14036 11962 14088 11968
rect 14048 11550 14076 11962
rect 14416 11686 14444 13662
rect 14404 11680 14456 11686
rect 14404 11622 14456 11628
rect 14036 11544 14088 11550
rect 14036 11486 14088 11492
rect 13760 11000 13812 11006
rect 13760 10942 13812 10948
rect 13576 10864 13628 10870
rect 13576 10806 13628 10812
rect 13588 10530 13616 10806
rect 13772 10598 13800 10942
rect 13760 10592 13812 10598
rect 13760 10534 13812 10540
rect 13576 10524 13628 10530
rect 13576 10466 13628 10472
rect 13588 9986 13616 10466
rect 13772 10122 13800 10534
rect 13760 10116 13812 10122
rect 13760 10058 13812 10064
rect 13576 9980 13628 9986
rect 13576 9922 13628 9928
rect 14048 7606 14076 11486
rect 14128 10320 14180 10326
rect 14128 10262 14180 10268
rect 14140 10122 14168 10262
rect 14508 10122 14536 14750
rect 14128 10116 14180 10122
rect 14128 10058 14180 10064
rect 14496 10116 14548 10122
rect 14496 10058 14548 10064
rect 14508 9850 14536 10058
rect 14496 9844 14548 9850
rect 14496 9786 14548 9792
rect 14600 9356 14628 16400
rect 14784 16310 14812 16790
rect 14968 16650 14996 17062
rect 14956 16644 15008 16650
rect 14956 16586 15008 16592
rect 14772 16304 14824 16310
rect 14772 16246 14824 16252
rect 14968 15562 14996 16586
rect 14956 15556 15008 15562
rect 14956 15498 15008 15504
rect 14864 15284 14916 15290
rect 14864 15226 14916 15232
rect 14680 14944 14732 14950
rect 14680 14886 14732 14892
rect 14692 13930 14720 14886
rect 14680 13924 14732 13930
rect 14680 13866 14732 13872
rect 14876 13726 14904 15226
rect 14968 15222 14996 15498
rect 14956 15216 15008 15222
rect 14956 15158 15008 15164
rect 14968 14950 14996 15158
rect 14956 14944 15008 14950
rect 14956 14886 15008 14892
rect 14956 14672 15008 14678
rect 14956 14614 15008 14620
rect 14968 14474 14996 14614
rect 14956 14468 15008 14474
rect 14956 14410 15008 14416
rect 15152 14214 15180 21686
rect 15336 21410 15364 25834
rect 15520 25694 15548 26174
rect 15508 25688 15560 25694
rect 15508 25630 15560 25636
rect 15600 25620 15652 25626
rect 15600 25562 15652 25568
rect 15612 25014 15640 25562
rect 15600 25008 15652 25014
rect 15600 24950 15652 24956
rect 15612 24674 15640 24950
rect 15600 24668 15652 24674
rect 15600 24610 15652 24616
rect 15784 24668 15836 24674
rect 15784 24610 15836 24616
rect 15612 24130 15640 24610
rect 15796 24266 15824 24610
rect 15784 24260 15836 24266
rect 15784 24202 15836 24208
rect 15600 24124 15652 24130
rect 15600 24066 15652 24072
rect 15796 23874 15824 24202
rect 15704 23846 15824 23874
rect 15704 22634 15732 23846
rect 15692 22628 15744 22634
rect 15692 22570 15744 22576
rect 15704 22362 15732 22570
rect 15980 22498 16008 27194
rect 16440 26850 16468 27466
rect 16624 27190 16652 27670
rect 16808 27462 16836 27874
rect 17176 27530 17204 28486
rect 17360 28414 17388 29302
rect 17636 29094 17664 29370
rect 17912 29162 17940 29438
rect 18372 29366 18400 30390
rect 18864 30348 19184 30368
rect 18864 30346 18876 30348
rect 18932 30346 18956 30348
rect 19012 30346 19036 30348
rect 19092 30346 19116 30348
rect 19172 30346 19184 30348
rect 18864 30294 18870 30346
rect 18932 30294 18934 30346
rect 19114 30294 19116 30346
rect 19178 30294 19184 30346
rect 18864 30292 18876 30294
rect 18932 30292 18956 30294
rect 19012 30292 19036 30294
rect 19092 30292 19116 30294
rect 19172 30292 19184 30294
rect 18864 30272 19184 30292
rect 18544 30244 18596 30250
rect 18544 30186 18596 30192
rect 18360 29360 18412 29366
rect 18360 29302 18412 29308
rect 17900 29156 17952 29162
rect 17900 29098 17952 29104
rect 17624 29088 17676 29094
rect 17624 29030 17676 29036
rect 17532 28952 17584 28958
rect 17532 28894 17584 28900
rect 17544 28482 17572 28894
rect 17636 28550 17664 29030
rect 18084 28816 18136 28822
rect 18084 28758 18136 28764
rect 17624 28544 17676 28550
rect 17624 28486 17676 28492
rect 17532 28476 17584 28482
rect 17532 28418 17584 28424
rect 17348 28408 17400 28414
rect 17348 28350 17400 28356
rect 17164 27524 17216 27530
rect 17164 27466 17216 27472
rect 16796 27456 16848 27462
rect 16796 27398 16848 27404
rect 16888 27388 16940 27394
rect 16888 27330 16940 27336
rect 16612 27184 16664 27190
rect 16612 27126 16664 27132
rect 16624 26850 16652 27126
rect 16428 26844 16480 26850
rect 16428 26786 16480 26792
rect 16612 26844 16664 26850
rect 16612 26786 16664 26792
rect 16440 26442 16468 26786
rect 16624 26442 16652 26786
rect 16796 26640 16848 26646
rect 16796 26582 16848 26588
rect 16808 26442 16836 26582
rect 16428 26436 16480 26442
rect 16428 26378 16480 26384
rect 16612 26436 16664 26442
rect 16612 26378 16664 26384
rect 16796 26436 16848 26442
rect 16796 26378 16848 26384
rect 16428 26300 16480 26306
rect 16428 26242 16480 26248
rect 16336 25688 16388 25694
rect 16336 25630 16388 25636
rect 16244 25552 16296 25558
rect 16244 25494 16296 25500
rect 16256 25218 16284 25494
rect 16348 25286 16376 25630
rect 16440 25558 16468 26242
rect 16808 25762 16836 26378
rect 16796 25756 16848 25762
rect 16796 25698 16848 25704
rect 16428 25552 16480 25558
rect 16428 25494 16480 25500
rect 16440 25354 16468 25494
rect 16428 25348 16480 25354
rect 16428 25290 16480 25296
rect 16808 25286 16836 25698
rect 16336 25280 16388 25286
rect 16336 25222 16388 25228
rect 16796 25280 16848 25286
rect 16796 25222 16848 25228
rect 16244 25212 16296 25218
rect 16244 25154 16296 25160
rect 16900 25082 16928 27330
rect 17360 25558 17388 28350
rect 17544 28006 17572 28418
rect 18096 28414 18124 28758
rect 18084 28408 18136 28414
rect 18084 28350 18136 28356
rect 17992 28272 18044 28278
rect 17992 28214 18044 28220
rect 18004 28074 18032 28214
rect 17992 28068 18044 28074
rect 17992 28010 18044 28016
rect 17532 28000 17584 28006
rect 17532 27942 17584 27948
rect 17808 26232 17860 26238
rect 17808 26174 17860 26180
rect 17716 26096 17768 26102
rect 17716 26038 17768 26044
rect 17728 25694 17756 26038
rect 17716 25688 17768 25694
rect 17716 25630 17768 25636
rect 17348 25552 17400 25558
rect 17348 25494 17400 25500
rect 17360 25150 17388 25494
rect 17348 25144 17400 25150
rect 17348 25086 17400 25092
rect 16888 25076 16940 25082
rect 16888 25018 16940 25024
rect 16980 25008 17032 25014
rect 16980 24950 17032 24956
rect 17072 25008 17124 25014
rect 17072 24950 17124 24956
rect 16992 24742 17020 24950
rect 16980 24736 17032 24742
rect 16980 24678 17032 24684
rect 16060 24600 16112 24606
rect 16060 24542 16112 24548
rect 16072 24266 16100 24542
rect 16992 24266 17020 24678
rect 16060 24260 16112 24266
rect 16060 24202 16112 24208
rect 16980 24260 17032 24266
rect 16980 24202 17032 24208
rect 17084 24198 17112 24950
rect 17072 24192 17124 24198
rect 17072 24134 17124 24140
rect 15968 22492 16020 22498
rect 15968 22434 16020 22440
rect 16336 22492 16388 22498
rect 16336 22434 16388 22440
rect 15692 22356 15744 22362
rect 15692 22298 15744 22304
rect 16348 21750 16376 22434
rect 16520 22288 16572 22294
rect 16520 22230 16572 22236
rect 16612 22288 16664 22294
rect 16612 22230 16664 22236
rect 16532 22090 16560 22230
rect 16520 22084 16572 22090
rect 16520 22026 16572 22032
rect 16624 22022 16652 22230
rect 16612 22016 16664 22022
rect 16612 21958 16664 21964
rect 16336 21744 16388 21750
rect 16336 21686 16388 21692
rect 15324 21404 15376 21410
rect 15324 21346 15376 21352
rect 16244 21268 16296 21274
rect 16244 21210 16296 21216
rect 16256 21002 16284 21210
rect 16244 20996 16296 21002
rect 16244 20938 16296 20944
rect 16348 20304 16376 21686
rect 17360 21546 17388 25086
rect 17716 24600 17768 24606
rect 17716 24542 17768 24548
rect 17728 24266 17756 24542
rect 17716 24260 17768 24266
rect 17716 24202 17768 24208
rect 17624 22288 17676 22294
rect 17624 22230 17676 22236
rect 17636 21886 17664 22230
rect 17624 21880 17676 21886
rect 17624 21822 17676 21828
rect 17348 21540 17400 21546
rect 17348 21482 17400 21488
rect 16428 21472 16480 21478
rect 16428 21414 16480 21420
rect 16440 21002 16468 21414
rect 16520 21404 16572 21410
rect 16520 21346 16572 21352
rect 16428 20996 16480 21002
rect 16428 20938 16480 20944
rect 16532 20769 16560 21346
rect 17072 21336 17124 21342
rect 17072 21278 17124 21284
rect 17084 21002 17112 21278
rect 17072 20996 17124 21002
rect 17072 20938 17124 20944
rect 17164 20996 17216 21002
rect 17164 20938 17216 20944
rect 16518 20760 16574 20769
rect 16518 20695 16574 20704
rect 16532 20662 16560 20695
rect 16520 20656 16572 20662
rect 16520 20598 16572 20604
rect 16532 20458 16560 20598
rect 17084 20458 17112 20938
rect 17176 20798 17204 20938
rect 17360 20798 17388 21482
rect 17440 21336 17492 21342
rect 17440 21278 17492 21284
rect 17164 20792 17216 20798
rect 17164 20734 17216 20740
rect 17348 20792 17400 20798
rect 17348 20734 17400 20740
rect 16520 20452 16572 20458
rect 16520 20394 16572 20400
rect 17072 20452 17124 20458
rect 17072 20394 17124 20400
rect 16428 20316 16480 20322
rect 16348 20276 16428 20304
rect 16428 20258 16480 20264
rect 16440 19574 16468 20258
rect 16532 19914 16560 20394
rect 17360 20186 17388 20734
rect 17452 20322 17480 21278
rect 17636 20848 17664 21822
rect 17716 20860 17768 20866
rect 17636 20820 17716 20848
rect 17716 20802 17768 20808
rect 17820 20322 17848 26174
rect 18268 26096 18320 26102
rect 18268 26038 18320 26044
rect 18176 25688 18228 25694
rect 18176 25630 18228 25636
rect 17900 25008 17952 25014
rect 17900 24950 17952 24956
rect 17912 24674 17940 24950
rect 18188 24810 18216 25630
rect 18280 25626 18308 26038
rect 18452 25756 18504 25762
rect 18452 25698 18504 25704
rect 18268 25620 18320 25626
rect 18268 25562 18320 25568
rect 18280 25082 18308 25562
rect 18360 25212 18412 25218
rect 18360 25154 18412 25160
rect 18268 25076 18320 25082
rect 18268 25018 18320 25024
rect 18176 24804 18228 24810
rect 18176 24746 18228 24752
rect 17900 24668 17952 24674
rect 17900 24610 17952 24616
rect 17992 24600 18044 24606
rect 17992 24542 18044 24548
rect 18004 24198 18032 24542
rect 17992 24192 18044 24198
rect 17992 24134 18044 24140
rect 18268 23512 18320 23518
rect 18268 23454 18320 23460
rect 17992 23376 18044 23382
rect 17992 23318 18044 23324
rect 18004 23178 18032 23318
rect 17992 23172 18044 23178
rect 17992 23114 18044 23120
rect 18084 22900 18136 22906
rect 18084 22842 18136 22848
rect 18096 21954 18124 22842
rect 18280 22838 18308 23454
rect 18268 22832 18320 22838
rect 18268 22774 18320 22780
rect 18084 21948 18136 21954
rect 18084 21890 18136 21896
rect 18280 21818 18308 22774
rect 18372 21886 18400 25154
rect 18464 24470 18492 25698
rect 18452 24464 18504 24470
rect 18452 24406 18504 24412
rect 18360 21880 18412 21886
rect 18360 21822 18412 21828
rect 18268 21812 18320 21818
rect 18268 21754 18320 21760
rect 18360 21404 18412 21410
rect 18360 21346 18412 21352
rect 18372 21002 18400 21346
rect 18360 20996 18412 21002
rect 18360 20938 18412 20944
rect 18084 20724 18136 20730
rect 18084 20666 18136 20672
rect 18096 20390 18124 20666
rect 18084 20384 18136 20390
rect 18084 20326 18136 20332
rect 17440 20316 17492 20322
rect 17440 20258 17492 20264
rect 17808 20316 17860 20322
rect 17808 20258 17860 20264
rect 17348 20180 17400 20186
rect 17348 20122 17400 20128
rect 16520 19908 16572 19914
rect 16520 19850 16572 19856
rect 17820 19846 17848 20258
rect 18096 19914 18124 20326
rect 18084 19908 18136 19914
rect 18084 19850 18136 19856
rect 18556 19846 18584 30186
rect 20488 30114 20516 31664
rect 21776 31662 21988 31664
rect 19004 30108 19056 30114
rect 19004 30050 19056 30056
rect 20476 30108 20528 30114
rect 20476 30050 20528 30056
rect 19016 29706 19044 30050
rect 19554 29736 19610 29745
rect 19004 29700 19056 29706
rect 20488 29706 20516 30050
rect 20660 29904 20712 29910
rect 20660 29846 20712 29852
rect 19554 29671 19610 29680
rect 20476 29700 20528 29706
rect 19004 29642 19056 29648
rect 19568 29502 19596 29671
rect 20476 29642 20528 29648
rect 20672 29502 20700 29846
rect 19556 29496 19608 29502
rect 19556 29438 19608 29444
rect 20660 29496 20712 29502
rect 20660 29438 20712 29444
rect 21120 29428 21172 29434
rect 21120 29370 21172 29376
rect 20108 29360 20160 29366
rect 20108 29302 20160 29308
rect 18864 29260 19184 29280
rect 18864 29258 18876 29260
rect 18932 29258 18956 29260
rect 19012 29258 19036 29260
rect 19092 29258 19116 29260
rect 19172 29258 19184 29260
rect 18864 29206 18870 29258
rect 18932 29206 18934 29258
rect 19114 29206 19116 29258
rect 19178 29206 19184 29258
rect 18864 29204 18876 29206
rect 18932 29204 18956 29206
rect 19012 29204 19036 29206
rect 19092 29204 19116 29206
rect 19172 29204 19184 29206
rect 18864 29184 19184 29204
rect 20120 29026 20148 29302
rect 21132 29026 21160 29370
rect 18728 29020 18780 29026
rect 18728 28962 18780 28968
rect 20108 29020 20160 29026
rect 20108 28962 20160 28968
rect 21120 29020 21172 29026
rect 21120 28962 21172 28968
rect 18740 28482 18768 28962
rect 19280 28816 19332 28822
rect 19280 28758 19332 28764
rect 18728 28476 18780 28482
rect 18728 28418 18780 28424
rect 18740 28074 18768 28418
rect 18864 28172 19184 28192
rect 18864 28170 18876 28172
rect 18932 28170 18956 28172
rect 19012 28170 19036 28172
rect 19092 28170 19116 28172
rect 19172 28170 19184 28172
rect 18864 28118 18870 28170
rect 18932 28118 18934 28170
rect 19114 28118 19116 28170
rect 19178 28118 19184 28170
rect 18864 28116 18876 28118
rect 18932 28116 18956 28118
rect 19012 28116 19036 28118
rect 19092 28116 19116 28118
rect 19172 28116 19184 28118
rect 18864 28096 19184 28116
rect 19292 28074 19320 28758
rect 20120 28346 20148 28962
rect 20292 28952 20344 28958
rect 20292 28894 20344 28900
rect 19372 28340 19424 28346
rect 19372 28282 19424 28288
rect 20108 28340 20160 28346
rect 20108 28282 20160 28288
rect 18728 28068 18780 28074
rect 18728 28010 18780 28016
rect 19280 28068 19332 28074
rect 19280 28010 19332 28016
rect 19384 28006 19412 28282
rect 19372 28000 19424 28006
rect 19372 27942 19424 27948
rect 18864 27084 19184 27104
rect 18864 27082 18876 27084
rect 18932 27082 18956 27084
rect 19012 27082 19036 27084
rect 19092 27082 19116 27084
rect 19172 27082 19184 27084
rect 18864 27030 18870 27082
rect 18932 27030 18934 27082
rect 19114 27030 19116 27082
rect 19178 27030 19184 27082
rect 18864 27028 18876 27030
rect 18932 27028 18956 27030
rect 19012 27028 19036 27030
rect 19092 27028 19116 27030
rect 19172 27028 19184 27030
rect 18864 27008 19184 27028
rect 20120 26238 20148 28282
rect 20304 28278 20332 28894
rect 20292 28272 20344 28278
rect 20292 28214 20344 28220
rect 20936 28000 20988 28006
rect 20936 27942 20988 27948
rect 20200 27932 20252 27938
rect 20200 27874 20252 27880
rect 20212 27394 20240 27874
rect 20948 27530 20976 27942
rect 20936 27524 20988 27530
rect 20936 27466 20988 27472
rect 20200 27388 20252 27394
rect 20200 27330 20252 27336
rect 21132 27326 21160 28962
rect 21120 27320 21172 27326
rect 21120 27262 21172 27268
rect 20660 27184 20712 27190
rect 20660 27126 20712 27132
rect 20108 26232 20160 26238
rect 20108 26174 20160 26180
rect 20200 26232 20252 26238
rect 20200 26174 20252 26180
rect 18864 25996 19184 26016
rect 18864 25994 18876 25996
rect 18932 25994 18956 25996
rect 19012 25994 19036 25996
rect 19092 25994 19116 25996
rect 19172 25994 19184 25996
rect 18864 25942 18870 25994
rect 18932 25942 18934 25994
rect 19114 25942 19116 25994
rect 19178 25942 19184 25994
rect 18864 25940 18876 25942
rect 18932 25940 18956 25942
rect 19012 25940 19036 25942
rect 19092 25940 19116 25942
rect 19172 25940 19184 25942
rect 18864 25920 19184 25940
rect 20212 25762 20240 26174
rect 20200 25756 20252 25762
rect 20200 25698 20252 25704
rect 20212 25354 20240 25698
rect 20384 25688 20436 25694
rect 20384 25630 20436 25636
rect 20200 25348 20252 25354
rect 20200 25290 20252 25296
rect 20396 25286 20424 25630
rect 18636 25280 18688 25286
rect 18636 25222 18688 25228
rect 20384 25280 20436 25286
rect 20384 25222 20436 25228
rect 18648 23042 18676 25222
rect 20672 25150 20700 27126
rect 21396 26776 21448 26782
rect 21396 26718 21448 26724
rect 21408 26442 21436 26718
rect 21396 26436 21448 26442
rect 21396 26378 21448 26384
rect 20936 26164 20988 26170
rect 20936 26106 20988 26112
rect 20292 25144 20344 25150
rect 20292 25086 20344 25092
rect 20660 25144 20712 25150
rect 20660 25086 20712 25092
rect 19372 25076 19424 25082
rect 19372 25018 19424 25024
rect 18864 24908 19184 24928
rect 18864 24906 18876 24908
rect 18932 24906 18956 24908
rect 19012 24906 19036 24908
rect 19092 24906 19116 24908
rect 19172 24906 19184 24908
rect 18864 24854 18870 24906
rect 18932 24854 18934 24906
rect 19114 24854 19116 24906
rect 19178 24854 19184 24906
rect 18864 24852 18876 24854
rect 18932 24852 18956 24854
rect 19012 24852 19036 24854
rect 19092 24852 19116 24854
rect 19172 24852 19184 24854
rect 18864 24832 19184 24852
rect 19384 24674 19412 25018
rect 18728 24668 18780 24674
rect 18728 24610 18780 24616
rect 19372 24668 19424 24674
rect 19372 24610 19424 24616
rect 18740 23586 18768 24610
rect 20304 24062 20332 25086
rect 20948 24674 20976 26106
rect 21408 25762 21436 26378
rect 21396 25756 21448 25762
rect 21396 25698 21448 25704
rect 21408 25354 21436 25698
rect 21396 25348 21448 25354
rect 21396 25290 21448 25296
rect 21672 25212 21724 25218
rect 21672 25154 21724 25160
rect 21684 24742 21712 25154
rect 21672 24736 21724 24742
rect 21672 24678 21724 24684
rect 20936 24668 20988 24674
rect 20936 24610 20988 24616
rect 20948 24266 20976 24610
rect 21212 24600 21264 24606
rect 21212 24542 21264 24548
rect 20936 24260 20988 24266
rect 20936 24202 20988 24208
rect 20292 24056 20344 24062
rect 20292 23998 20344 24004
rect 21224 23994 21252 24542
rect 21580 24464 21632 24470
rect 21580 24406 21632 24412
rect 19372 23988 19424 23994
rect 19372 23930 19424 23936
rect 21212 23988 21264 23994
rect 21212 23930 21264 23936
rect 18864 23820 19184 23840
rect 18864 23818 18876 23820
rect 18932 23818 18956 23820
rect 19012 23818 19036 23820
rect 19092 23818 19116 23820
rect 19172 23818 19184 23820
rect 18864 23766 18870 23818
rect 18932 23766 18934 23818
rect 19114 23766 19116 23818
rect 19178 23766 19184 23818
rect 18864 23764 18876 23766
rect 18932 23764 18956 23766
rect 19012 23764 19036 23766
rect 19092 23764 19116 23766
rect 19172 23764 19184 23766
rect 18864 23744 19184 23764
rect 19384 23722 19412 23930
rect 20016 23920 20068 23926
rect 20016 23862 20068 23868
rect 20028 23722 20056 23862
rect 19372 23716 19424 23722
rect 19372 23658 19424 23664
rect 20016 23716 20068 23722
rect 20016 23658 20068 23664
rect 18728 23580 18780 23586
rect 18728 23522 18780 23528
rect 18740 23178 18768 23522
rect 18728 23172 18780 23178
rect 18728 23114 18780 23120
rect 18636 23036 18688 23042
rect 18636 22978 18688 22984
rect 18648 22634 18676 22978
rect 19384 22906 19412 23658
rect 21592 23586 21620 24406
rect 21684 24266 21712 24678
rect 21672 24260 21724 24266
rect 21672 24202 21724 24208
rect 21580 23580 21632 23586
rect 21580 23522 21632 23528
rect 21488 23376 21540 23382
rect 21488 23318 21540 23324
rect 19372 22900 19424 22906
rect 19372 22842 19424 22848
rect 20660 22900 20712 22906
rect 20660 22842 20712 22848
rect 18864 22732 19184 22752
rect 18864 22730 18876 22732
rect 18932 22730 18956 22732
rect 19012 22730 19036 22732
rect 19092 22730 19116 22732
rect 19172 22730 19184 22732
rect 18864 22678 18870 22730
rect 18932 22678 18934 22730
rect 19114 22678 19116 22730
rect 19178 22678 19184 22730
rect 18864 22676 18876 22678
rect 18932 22676 18956 22678
rect 19012 22676 19036 22678
rect 19092 22676 19116 22678
rect 19172 22676 19184 22678
rect 18864 22656 19184 22676
rect 19384 22634 19412 22842
rect 18636 22628 18688 22634
rect 18636 22570 18688 22576
rect 19372 22628 19424 22634
rect 19372 22570 19424 22576
rect 20672 22294 20700 22842
rect 20660 22288 20712 22294
rect 20660 22230 20712 22236
rect 18728 21744 18780 21750
rect 18728 21686 18780 21692
rect 18740 21342 18768 21686
rect 18864 21644 19184 21664
rect 18864 21642 18876 21644
rect 18932 21642 18956 21644
rect 19012 21642 19036 21644
rect 19092 21642 19116 21644
rect 19172 21642 19184 21644
rect 18864 21590 18870 21642
rect 18932 21590 18934 21642
rect 19114 21590 19116 21642
rect 19178 21590 19184 21642
rect 18864 21588 18876 21590
rect 18932 21588 18956 21590
rect 19012 21588 19036 21590
rect 19092 21588 19116 21590
rect 19172 21588 19184 21590
rect 18864 21568 19184 21588
rect 19372 21404 19424 21410
rect 19372 21346 19424 21352
rect 18728 21336 18780 21342
rect 18728 21278 18780 21284
rect 19384 20730 19412 21346
rect 19372 20724 19424 20730
rect 19372 20666 19424 20672
rect 18864 20556 19184 20576
rect 18864 20554 18876 20556
rect 18932 20554 18956 20556
rect 19012 20554 19036 20556
rect 19092 20554 19116 20556
rect 19172 20554 19184 20556
rect 18864 20502 18870 20554
rect 18932 20502 18934 20554
rect 19114 20502 19116 20554
rect 19178 20502 19184 20554
rect 18864 20500 18876 20502
rect 18932 20500 18956 20502
rect 19012 20500 19036 20502
rect 19092 20500 19116 20502
rect 19172 20500 19184 20502
rect 18864 20480 19184 20500
rect 17808 19840 17860 19846
rect 17808 19782 17860 19788
rect 18544 19840 18596 19846
rect 18544 19782 18596 19788
rect 19924 19840 19976 19846
rect 19924 19782 19976 19788
rect 16428 19568 16480 19574
rect 16428 19510 16480 19516
rect 17820 19370 17848 19782
rect 18084 19568 18136 19574
rect 18084 19510 18136 19516
rect 19832 19568 19884 19574
rect 19832 19510 19884 19516
rect 17808 19364 17860 19370
rect 17808 19306 17860 19312
rect 15232 19296 15284 19302
rect 15232 19238 15284 19244
rect 16888 19296 16940 19302
rect 16888 19238 16940 19244
rect 15244 18826 15272 19238
rect 16152 19228 16204 19234
rect 16152 19170 16204 19176
rect 16612 19228 16664 19234
rect 16612 19170 16664 19176
rect 16164 18826 16192 19170
rect 15232 18820 15284 18826
rect 15232 18762 15284 18768
rect 16152 18820 16204 18826
rect 16152 18762 16204 18768
rect 15232 18616 15284 18622
rect 15232 18558 15284 18564
rect 15244 18146 15272 18558
rect 16164 18214 16192 18762
rect 16624 18486 16652 19170
rect 16900 18826 16928 19238
rect 16888 18820 16940 18826
rect 16888 18762 16940 18768
rect 16704 18616 16756 18622
rect 16704 18558 16756 18564
rect 16612 18480 16664 18486
rect 16612 18422 16664 18428
rect 16152 18208 16204 18214
rect 16152 18150 16204 18156
rect 15232 18140 15284 18146
rect 15232 18082 15284 18088
rect 16612 18140 16664 18146
rect 16612 18082 16664 18088
rect 15244 17194 15272 18082
rect 16428 17460 16480 17466
rect 16428 17402 16480 17408
rect 15968 17392 16020 17398
rect 15968 17334 16020 17340
rect 16060 17392 16112 17398
rect 16060 17334 16112 17340
rect 15232 17188 15284 17194
rect 15232 17130 15284 17136
rect 15980 17058 16008 17334
rect 15968 17052 16020 17058
rect 15968 16994 16020 17000
rect 15980 16650 16008 16994
rect 15968 16644 16020 16650
rect 15968 16586 16020 16592
rect 15232 16032 15284 16038
rect 15232 15974 15284 15980
rect 15968 16032 16020 16038
rect 15968 15974 16020 15980
rect 15244 15222 15272 15974
rect 15600 15964 15652 15970
rect 15652 15924 15732 15952
rect 15600 15906 15652 15912
rect 15704 15222 15732 15924
rect 15980 15562 16008 15974
rect 15968 15556 16020 15562
rect 15968 15498 16020 15504
rect 16072 15442 16100 17334
rect 16440 17058 16468 17402
rect 16624 17398 16652 18082
rect 16612 17392 16664 17398
rect 16612 17334 16664 17340
rect 16428 17052 16480 17058
rect 16428 16994 16480 17000
rect 16440 16514 16468 16994
rect 16520 16984 16572 16990
rect 16520 16926 16572 16932
rect 16532 16650 16560 16926
rect 16520 16644 16572 16650
rect 16520 16586 16572 16592
rect 16428 16508 16480 16514
rect 16428 16450 16480 16456
rect 15980 15414 16100 15442
rect 15232 15216 15284 15222
rect 15232 15158 15284 15164
rect 15692 15216 15744 15222
rect 15692 15158 15744 15164
rect 14968 14186 15180 14214
rect 14864 13720 14916 13726
rect 14864 13662 14916 13668
rect 14680 13108 14732 13114
rect 14680 13050 14732 13056
rect 14692 10530 14720 13050
rect 14864 13040 14916 13046
rect 14864 12982 14916 12988
rect 14772 12700 14824 12706
rect 14772 12642 14824 12648
rect 14784 12298 14812 12642
rect 14772 12292 14824 12298
rect 14772 12234 14824 12240
rect 14772 11000 14824 11006
rect 14772 10942 14824 10948
rect 14784 10530 14812 10942
rect 14876 10666 14904 12982
rect 14968 12842 14996 14186
rect 15048 14128 15100 14134
rect 15244 14116 15272 15158
rect 15600 14468 15652 14474
rect 15600 14410 15652 14416
rect 15416 14400 15468 14406
rect 15416 14342 15468 14348
rect 15100 14088 15272 14116
rect 15048 14070 15100 14076
rect 15060 13794 15088 14070
rect 15140 13856 15192 13862
rect 15140 13798 15192 13804
rect 15324 13856 15376 13862
rect 15324 13798 15376 13804
rect 15048 13788 15100 13794
rect 15048 13730 15100 13736
rect 15060 13114 15088 13730
rect 15048 13108 15100 13114
rect 15048 13050 15100 13056
rect 14956 12836 15008 12842
rect 14956 12778 15008 12784
rect 14956 12700 15008 12706
rect 14956 12642 15008 12648
rect 14968 11958 14996 12642
rect 14956 11952 15008 11958
rect 14956 11894 15008 11900
rect 14968 11210 14996 11894
rect 14956 11204 15008 11210
rect 14956 11146 15008 11152
rect 14864 10660 14916 10666
rect 14864 10602 14916 10608
rect 14680 10524 14732 10530
rect 14680 10466 14732 10472
rect 14772 10524 14824 10530
rect 14772 10466 14824 10472
rect 14692 9578 14720 10466
rect 14784 10122 14812 10466
rect 14864 10320 14916 10326
rect 14864 10262 14916 10268
rect 14772 10116 14824 10122
rect 14772 10058 14824 10064
rect 14772 9776 14824 9782
rect 14772 9718 14824 9724
rect 14680 9572 14732 9578
rect 14680 9514 14732 9520
rect 14784 9510 14812 9718
rect 14772 9504 14824 9510
rect 14772 9446 14824 9452
rect 14232 9328 14628 9356
rect 14036 7600 14088 7606
rect 14036 7542 14088 7548
rect 12760 6858 12788 6998
rect 13496 6982 13616 7010
rect 12288 6852 12340 6858
rect 12288 6794 12340 6800
rect 12748 6852 12800 6858
rect 12748 6794 12800 6800
rect 12196 6716 12248 6722
rect 12196 6658 12248 6664
rect 11552 6580 11604 6586
rect 11552 6522 11604 6528
rect 10816 6512 10868 6518
rect 10816 6454 10868 6460
rect 10828 6110 10856 6454
rect 11276 6308 11328 6314
rect 11276 6250 11328 6256
rect 10724 6104 10776 6110
rect 10724 6046 10776 6052
rect 10816 6104 10868 6110
rect 10816 6046 10868 6052
rect 10736 5022 10764 6046
rect 10828 5566 10856 6046
rect 10816 5560 10868 5566
rect 10816 5502 10868 5508
rect 10908 5492 10960 5498
rect 10908 5434 10960 5440
rect 10920 5090 10948 5434
rect 11288 5158 11316 6250
rect 11564 5770 11592 6522
rect 12208 6314 12236 6658
rect 13208 6648 13260 6654
rect 13208 6590 13260 6596
rect 12196 6308 12248 6314
rect 12196 6250 12248 6256
rect 11552 5764 11604 5770
rect 11552 5706 11604 5712
rect 11460 5696 11512 5702
rect 11460 5638 11512 5644
rect 11276 5152 11328 5158
rect 11276 5094 11328 5100
rect 10908 5084 10960 5090
rect 10908 5026 10960 5032
rect 10724 5016 10776 5022
rect 10724 4958 10776 4964
rect 10736 4342 10764 4958
rect 10920 4682 10948 5026
rect 11288 4682 11316 5094
rect 11472 5022 11500 5638
rect 12208 5566 12236 6250
rect 13220 6178 13248 6590
rect 13208 6172 13260 6178
rect 13208 6114 13260 6120
rect 12288 6036 12340 6042
rect 12288 5978 12340 5984
rect 12196 5560 12248 5566
rect 12196 5502 12248 5508
rect 11460 5016 11512 5022
rect 11460 4958 11512 4964
rect 10908 4676 10960 4682
rect 10908 4618 10960 4624
rect 11276 4676 11328 4682
rect 11276 4618 11328 4624
rect 11920 4676 11972 4682
rect 11920 4618 11972 4624
rect 11932 4546 11960 4618
rect 11092 4540 11144 4546
rect 11092 4482 11144 4488
rect 11920 4540 11972 4546
rect 11920 4482 11972 4488
rect 10724 4336 10776 4342
rect 10724 4278 10776 4284
rect 11000 4132 11052 4138
rect 11000 4074 11052 4080
rect 10632 3860 10684 3866
rect 10632 3802 10684 3808
rect 10356 3384 10408 3390
rect 10356 3326 10408 3332
rect 10540 3384 10592 3390
rect 11012 3361 11040 4074
rect 10540 3326 10592 3332
rect 10998 3352 11054 3361
rect 10368 3050 10396 3326
rect 10998 3287 11054 3296
rect 10356 3044 10408 3050
rect 10356 2986 10408 2992
rect 11104 2914 11132 4482
rect 12300 4478 12328 5978
rect 12380 5968 12432 5974
rect 12380 5910 12432 5916
rect 12392 5566 12420 5910
rect 13220 5770 13248 6114
rect 13484 6104 13536 6110
rect 13484 6046 13536 6052
rect 13208 5764 13260 5770
rect 13208 5706 13260 5712
rect 12932 5628 12984 5634
rect 12932 5570 12984 5576
rect 12380 5560 12432 5566
rect 12380 5502 12432 5508
rect 12392 4886 12420 5502
rect 12380 4880 12432 4886
rect 12380 4822 12432 4828
rect 12392 4554 12420 4822
rect 12392 4526 12604 4554
rect 12288 4472 12340 4478
rect 12288 4414 12340 4420
rect 11736 4404 11788 4410
rect 11736 4346 11788 4352
rect 11184 4336 11236 4342
rect 11184 4278 11236 4284
rect 11092 2908 11144 2914
rect 11092 2850 11144 2856
rect 10356 2296 10408 2302
rect 10356 2238 10408 2244
rect 10368 1962 10396 2238
rect 11104 2234 11132 2850
rect 11196 2302 11224 4278
rect 11748 3934 11776 4346
rect 12012 3996 12064 4002
rect 12012 3938 12064 3944
rect 11736 3928 11788 3934
rect 11736 3870 11788 3876
rect 11644 3860 11696 3866
rect 11644 3802 11696 3808
rect 11276 3792 11328 3798
rect 11276 3734 11328 3740
rect 11288 3594 11316 3734
rect 11276 3588 11328 3594
rect 11276 3530 11328 3536
rect 11184 2296 11236 2302
rect 11184 2238 11236 2244
rect 11092 2228 11144 2234
rect 11092 2170 11144 2176
rect 10356 1956 10408 1962
rect 10356 1898 10408 1904
rect 10368 1418 10396 1898
rect 11104 1826 11132 2170
rect 11092 1820 11144 1826
rect 11092 1762 11144 1768
rect 11288 1758 11316 3530
rect 11656 3254 11684 3802
rect 11748 3769 11776 3870
rect 11734 3760 11790 3769
rect 11734 3695 11790 3704
rect 11748 3458 11776 3695
rect 12024 3526 12052 3938
rect 12012 3520 12064 3526
rect 12012 3462 12064 3468
rect 11736 3452 11788 3458
rect 11736 3394 11788 3400
rect 11736 3316 11788 3322
rect 11736 3258 11788 3264
rect 11644 3248 11696 3254
rect 11644 3190 11696 3196
rect 11656 2914 11684 3190
rect 11748 2982 11776 3258
rect 11828 3248 11880 3254
rect 11828 3190 11880 3196
rect 11840 3050 11868 3190
rect 12024 3050 12052 3462
rect 12300 3390 12328 4414
rect 12380 4064 12432 4070
rect 12380 4006 12432 4012
rect 12392 3526 12420 4006
rect 12380 3520 12432 3526
rect 12576 3497 12604 4526
rect 12380 3462 12432 3468
rect 12562 3488 12618 3497
rect 12392 3390 12420 3462
rect 12562 3423 12618 3432
rect 12944 3390 12972 5570
rect 13496 5430 13524 6046
rect 13588 5634 13616 6982
rect 13944 6716 13996 6722
rect 13944 6658 13996 6664
rect 13576 5628 13628 5634
rect 13576 5570 13628 5576
rect 13484 5424 13536 5430
rect 13484 5366 13536 5372
rect 13852 5424 13904 5430
rect 13852 5366 13904 5372
rect 13392 4336 13444 4342
rect 13392 4278 13444 4284
rect 13116 3520 13168 3526
rect 13116 3462 13168 3468
rect 12104 3384 12156 3390
rect 12104 3326 12156 3332
rect 12288 3384 12340 3390
rect 12288 3326 12340 3332
rect 12380 3384 12432 3390
rect 12380 3326 12432 3332
rect 12932 3384 12984 3390
rect 12932 3326 12984 3332
rect 11828 3044 11880 3050
rect 11828 2986 11880 2992
rect 12012 3044 12064 3050
rect 12012 2986 12064 2992
rect 11736 2976 11788 2982
rect 11736 2918 11788 2924
rect 11644 2908 11696 2914
rect 11644 2850 11696 2856
rect 11656 2148 11684 2850
rect 11748 2438 11776 2918
rect 11840 2506 11868 2986
rect 12116 2982 12144 3326
rect 13128 2982 13156 3462
rect 13404 3050 13432 4278
rect 13864 4138 13892 5366
rect 13852 4132 13904 4138
rect 13852 4074 13904 4080
rect 13864 3526 13892 4074
rect 13852 3520 13904 3526
rect 13852 3462 13904 3468
rect 13484 3316 13536 3322
rect 13484 3258 13536 3264
rect 13392 3044 13444 3050
rect 13392 2986 13444 2992
rect 12104 2976 12156 2982
rect 12104 2918 12156 2924
rect 13116 2976 13168 2982
rect 13116 2918 13168 2924
rect 11828 2500 11880 2506
rect 11828 2442 11880 2448
rect 11736 2432 11788 2438
rect 11736 2374 11788 2380
rect 11736 2160 11788 2166
rect 11656 2120 11736 2148
rect 11736 2102 11788 2108
rect 11748 1758 11776 2102
rect 13128 1894 13156 2918
rect 13392 2704 13444 2710
rect 13392 2646 13444 2652
rect 13404 2506 13432 2646
rect 13392 2500 13444 2506
rect 13392 2442 13444 2448
rect 13496 2370 13524 3258
rect 13576 3248 13628 3254
rect 13576 3190 13628 3196
rect 13484 2364 13536 2370
rect 13484 2306 13536 2312
rect 13484 2228 13536 2234
rect 13484 2170 13536 2176
rect 13496 1894 13524 2170
rect 13588 1962 13616 3190
rect 13576 1956 13628 1962
rect 13576 1898 13628 1904
rect 13116 1888 13168 1894
rect 13116 1830 13168 1836
rect 13484 1888 13536 1894
rect 13484 1830 13536 1836
rect 13956 1758 13984 6658
rect 11276 1752 11328 1758
rect 11276 1694 11328 1700
rect 11736 1752 11788 1758
rect 11736 1694 11788 1700
rect 13944 1752 13996 1758
rect 13944 1694 13996 1700
rect 10356 1412 10408 1418
rect 10356 1354 10408 1360
rect 11748 1350 11776 1694
rect 12748 1616 12800 1622
rect 12748 1558 12800 1564
rect 11736 1344 11788 1350
rect 11736 1286 11788 1292
rect 12760 1078 12788 1558
rect 11460 1072 11512 1078
rect 11460 1014 11512 1020
rect 12748 1072 12800 1078
rect 12748 1014 12800 1020
rect 10184 590 10304 618
rect 10184 482 10212 590
rect 10000 454 10212 482
rect 10000 424 10028 454
rect 11472 424 11500 1014
rect 12760 449 12788 509
rect 12746 440 12802 449
rect 3504 372 3516 374
rect 3572 372 3596 374
rect 3652 372 3676 374
rect 3732 372 3756 374
rect 3812 372 3824 374
rect 3504 352 3824 372
rect 4438 0 4550 424
rect 5910 0 6022 424
rect 7198 0 7310 424
rect 8670 0 8782 424
rect 9958 0 10070 424
rect 11430 0 11542 424
rect 12718 384 12746 424
rect 14232 424 14260 9328
rect 14588 9028 14640 9034
rect 14588 8970 14640 8976
rect 14600 8762 14628 8970
rect 14784 8830 14812 9446
rect 14772 8824 14824 8830
rect 14772 8766 14824 8772
rect 14588 8756 14640 8762
rect 14588 8698 14640 8704
rect 14772 8688 14824 8694
rect 14772 8630 14824 8636
rect 14312 8144 14364 8150
rect 14312 8086 14364 8092
rect 14324 7946 14352 8086
rect 14312 7940 14364 7946
rect 14312 7882 14364 7888
rect 14324 7742 14352 7882
rect 14312 7736 14364 7742
rect 14312 7678 14364 7684
rect 14404 7600 14456 7606
rect 14404 7542 14456 7548
rect 14680 7600 14732 7606
rect 14680 7542 14732 7548
rect 14416 4546 14444 7542
rect 14692 7266 14720 7542
rect 14680 7260 14732 7266
rect 14680 7202 14732 7208
rect 14692 6586 14720 7202
rect 14680 6580 14732 6586
rect 14680 6522 14732 6528
rect 14784 6178 14812 8630
rect 14876 7742 14904 10262
rect 15152 10074 15180 13798
rect 15336 13386 15364 13798
rect 15324 13380 15376 13386
rect 15324 13322 15376 13328
rect 15232 12700 15284 12706
rect 15232 12642 15284 12648
rect 15244 12298 15272 12642
rect 15232 12292 15284 12298
rect 15232 12234 15284 12240
rect 15428 11210 15456 14342
rect 15612 14202 15640 14410
rect 15600 14196 15652 14202
rect 15600 14138 15652 14144
rect 15704 11210 15732 15158
rect 15876 14196 15928 14202
rect 15876 14138 15928 14144
rect 15784 13176 15836 13182
rect 15784 13118 15836 13124
rect 15796 12774 15824 13118
rect 15784 12768 15836 12774
rect 15784 12710 15836 12716
rect 15416 11204 15468 11210
rect 15416 11146 15468 11152
rect 15692 11204 15744 11210
rect 15692 11146 15744 11152
rect 15428 11006 15456 11146
rect 15704 11074 15732 11146
rect 15692 11068 15744 11074
rect 15692 11010 15744 11016
rect 15416 11000 15468 11006
rect 15416 10942 15468 10948
rect 15152 10046 15364 10074
rect 15048 9844 15100 9850
rect 15048 9786 15100 9792
rect 14864 7736 14916 7742
rect 14864 7678 14916 7684
rect 14956 7260 15008 7266
rect 14876 7220 14956 7248
rect 14876 6518 14904 7220
rect 14956 7202 15008 7208
rect 15060 7146 15088 9786
rect 15140 7736 15192 7742
rect 15140 7678 15192 7684
rect 14968 7118 15088 7146
rect 14864 6512 14916 6518
rect 14864 6454 14916 6460
rect 14772 6172 14824 6178
rect 14772 6114 14824 6120
rect 14680 5764 14732 5770
rect 14680 5706 14732 5712
rect 14588 5560 14640 5566
rect 14588 5502 14640 5508
rect 14600 4614 14628 5502
rect 14692 5022 14720 5706
rect 14876 5702 14904 6454
rect 14864 5696 14916 5702
rect 14864 5638 14916 5644
rect 14680 5016 14732 5022
rect 14680 4958 14732 4964
rect 14692 4614 14720 4958
rect 14588 4608 14640 4614
rect 14508 4568 14588 4596
rect 14404 4540 14456 4546
rect 14404 4482 14456 4488
rect 14416 4342 14444 4482
rect 14508 4478 14536 4568
rect 14588 4550 14640 4556
rect 14680 4608 14732 4614
rect 14680 4550 14732 4556
rect 14496 4472 14548 4478
rect 14496 4414 14548 4420
rect 14404 4336 14456 4342
rect 14404 4278 14456 4284
rect 14404 3928 14456 3934
rect 14404 3870 14456 3876
rect 14416 3390 14444 3870
rect 14508 3866 14536 4414
rect 14968 4002 14996 7118
rect 15152 7062 15180 7678
rect 15140 7056 15192 7062
rect 15140 6998 15192 7004
rect 15152 6858 15180 6998
rect 15140 6852 15192 6858
rect 15140 6794 15192 6800
rect 15232 6852 15284 6858
rect 15232 6794 15284 6800
rect 15244 6314 15272 6794
rect 15336 6568 15364 10046
rect 15704 9034 15732 11010
rect 15888 9918 15916 14138
rect 15980 14134 16008 15414
rect 16716 14474 16744 18558
rect 17072 18480 17124 18486
rect 17072 18422 17124 18428
rect 17084 18146 17112 18422
rect 17072 18140 17124 18146
rect 17072 18082 17124 18088
rect 17440 18140 17492 18146
rect 17440 18082 17492 18088
rect 17084 17466 17112 18082
rect 17164 18072 17216 18078
rect 17164 18014 17216 18020
rect 17176 17738 17204 18014
rect 17164 17732 17216 17738
rect 17164 17674 17216 17680
rect 17072 17460 17124 17466
rect 17072 17402 17124 17408
rect 17452 16446 17480 18082
rect 17808 18072 17860 18078
rect 17808 18014 17860 18020
rect 17820 17534 17848 18014
rect 17808 17528 17860 17534
rect 17808 17470 17860 17476
rect 17532 17392 17584 17398
rect 17532 17334 17584 17340
rect 17544 16582 17572 17334
rect 17716 17052 17768 17058
rect 17716 16994 17768 17000
rect 17728 16854 17756 16994
rect 17820 16922 17848 17470
rect 17808 16916 17860 16922
rect 17808 16858 17860 16864
rect 17716 16848 17768 16854
rect 17716 16790 17768 16796
rect 17532 16576 17584 16582
rect 17532 16518 17584 16524
rect 17728 16446 17756 16790
rect 17440 16440 17492 16446
rect 17440 16382 17492 16388
rect 17716 16440 17768 16446
rect 17716 16382 17768 16388
rect 17452 16038 17480 16382
rect 17728 16038 17756 16382
rect 17440 16032 17492 16038
rect 17440 15974 17492 15980
rect 17716 16032 17768 16038
rect 17716 15974 17768 15980
rect 17820 15426 17848 16858
rect 17808 15420 17860 15426
rect 17808 15362 17860 15368
rect 16704 14468 16756 14474
rect 16704 14410 16756 14416
rect 17532 14468 17584 14474
rect 17532 14410 17584 14416
rect 16060 14400 16112 14406
rect 16060 14342 16112 14348
rect 16072 14270 16100 14342
rect 16060 14264 16112 14270
rect 16060 14206 16112 14212
rect 15968 14128 16020 14134
rect 15968 14070 16020 14076
rect 15980 9918 16008 14070
rect 16060 13856 16112 13862
rect 16060 13798 16112 13804
rect 17346 13824 17402 13833
rect 16072 13318 16100 13798
rect 17346 13759 17402 13768
rect 17360 13726 17388 13759
rect 16336 13720 16388 13726
rect 16336 13662 16388 13668
rect 17348 13720 17400 13726
rect 17348 13662 17400 13668
rect 16348 13386 16376 13662
rect 16336 13380 16388 13386
rect 16336 13322 16388 13328
rect 16060 13312 16112 13318
rect 16060 13254 16112 13260
rect 16428 13312 16480 13318
rect 16428 13254 16480 13260
rect 16152 13176 16204 13182
rect 16152 13118 16204 13124
rect 16164 12842 16192 13118
rect 16152 12836 16204 12842
rect 16152 12778 16204 12784
rect 16164 12298 16192 12778
rect 16336 12700 16388 12706
rect 16336 12642 16388 12648
rect 16152 12292 16204 12298
rect 16152 12234 16204 12240
rect 16348 11754 16376 12642
rect 16440 12502 16468 13254
rect 16612 13244 16664 13250
rect 16612 13186 16664 13192
rect 17256 13244 17308 13250
rect 17360 13232 17388 13662
rect 17308 13204 17388 13232
rect 17256 13186 17308 13192
rect 16624 12638 16652 13186
rect 17360 12774 17388 13204
rect 17544 13182 17572 14410
rect 18096 14214 18124 19510
rect 18864 19468 19184 19488
rect 18864 19466 18876 19468
rect 18932 19466 18956 19468
rect 19012 19466 19036 19468
rect 19092 19466 19116 19468
rect 19172 19466 19184 19468
rect 18864 19414 18870 19466
rect 18932 19414 18934 19466
rect 19114 19414 19116 19466
rect 19178 19414 19184 19466
rect 18864 19412 18876 19414
rect 18932 19412 18956 19414
rect 19012 19412 19036 19414
rect 19092 19412 19116 19414
rect 19172 19412 19184 19414
rect 18864 19392 19184 19412
rect 18864 18380 19184 18400
rect 18864 18378 18876 18380
rect 18932 18378 18956 18380
rect 19012 18378 19036 18380
rect 19092 18378 19116 18380
rect 19172 18378 19184 18380
rect 18864 18326 18870 18378
rect 18932 18326 18934 18378
rect 19114 18326 19116 18378
rect 19178 18326 19184 18378
rect 18864 18324 18876 18326
rect 18932 18324 18956 18326
rect 19012 18324 19036 18326
rect 19092 18324 19116 18326
rect 19172 18324 19184 18326
rect 18864 18304 19184 18324
rect 19844 17942 19872 19510
rect 18176 17936 18228 17942
rect 18176 17878 18228 17884
rect 19832 17936 19884 17942
rect 19832 17878 19884 17884
rect 18188 17602 18216 17878
rect 18176 17596 18228 17602
rect 18176 17538 18228 17544
rect 18188 17194 18216 17538
rect 18864 17292 19184 17312
rect 18864 17290 18876 17292
rect 18932 17290 18956 17292
rect 19012 17290 19036 17292
rect 19092 17290 19116 17292
rect 19172 17290 19184 17292
rect 18864 17238 18870 17290
rect 18932 17238 18934 17290
rect 19114 17238 19116 17290
rect 19178 17238 19184 17290
rect 18864 17236 18876 17238
rect 18932 17236 18956 17238
rect 19012 17236 19036 17238
rect 19092 17236 19116 17238
rect 19172 17236 19184 17238
rect 18864 17216 19184 17236
rect 18176 17188 18228 17194
rect 18176 17130 18228 17136
rect 18188 16650 18216 17130
rect 19556 17120 19608 17126
rect 19556 17062 19608 17068
rect 18820 17052 18872 17058
rect 18740 17012 18820 17040
rect 18544 16984 18596 16990
rect 18544 16926 18596 16932
rect 18176 16644 18228 16650
rect 18176 16586 18228 16592
rect 18452 16304 18504 16310
rect 18452 16246 18504 16252
rect 18464 15290 18492 16246
rect 18556 15902 18584 16926
rect 18740 16106 18768 17012
rect 18820 16994 18872 17000
rect 19004 16984 19056 16990
rect 19004 16926 19056 16932
rect 19016 16582 19044 16926
rect 19372 16848 19424 16854
rect 19372 16790 19424 16796
rect 19004 16576 19056 16582
rect 19004 16518 19056 16524
rect 19280 16508 19332 16514
rect 19280 16450 19332 16456
rect 18864 16204 19184 16224
rect 18864 16202 18876 16204
rect 18932 16202 18956 16204
rect 19012 16202 19036 16204
rect 19092 16202 19116 16204
rect 19172 16202 19184 16204
rect 18864 16150 18870 16202
rect 18932 16150 18934 16202
rect 19114 16150 19116 16202
rect 19178 16150 19184 16202
rect 18864 16148 18876 16150
rect 18932 16148 18956 16150
rect 19012 16148 19036 16150
rect 19092 16148 19116 16150
rect 19172 16148 19184 16150
rect 18864 16128 19184 16148
rect 19292 16106 19320 16450
rect 19384 16446 19412 16790
rect 19372 16440 19424 16446
rect 19372 16382 19424 16388
rect 18728 16100 18780 16106
rect 18728 16042 18780 16048
rect 19280 16100 19332 16106
rect 19280 16042 19332 16048
rect 18544 15896 18596 15902
rect 18544 15838 18596 15844
rect 18544 15420 18596 15426
rect 18740 15408 18768 16042
rect 18912 15760 18964 15766
rect 18912 15702 18964 15708
rect 19004 15760 19056 15766
rect 19004 15702 19056 15708
rect 18544 15362 18596 15368
rect 18648 15380 18768 15408
rect 18452 15284 18504 15290
rect 18452 15226 18504 15232
rect 18268 15216 18320 15222
rect 18268 15158 18320 15164
rect 18096 14186 18216 14214
rect 17900 14128 17952 14134
rect 17900 14070 17952 14076
rect 17532 13176 17584 13182
rect 17532 13118 17584 13124
rect 17624 13040 17676 13046
rect 17624 12982 17676 12988
rect 17348 12768 17400 12774
rect 17348 12710 17400 12716
rect 16612 12632 16664 12638
rect 16612 12574 16664 12580
rect 16980 12632 17032 12638
rect 16980 12574 17032 12580
rect 17348 12632 17400 12638
rect 17348 12574 17400 12580
rect 16428 12496 16480 12502
rect 16428 12438 16480 12444
rect 16440 11754 16468 12438
rect 16624 12298 16652 12574
rect 16992 12298 17020 12574
rect 16612 12292 16664 12298
rect 16612 12234 16664 12240
rect 16980 12292 17032 12298
rect 16980 12234 17032 12240
rect 16992 11754 17020 12234
rect 17360 12162 17388 12574
rect 17636 12162 17664 12982
rect 17348 12156 17400 12162
rect 17348 12098 17400 12104
rect 17624 12156 17676 12162
rect 17624 12098 17676 12104
rect 17440 12088 17492 12094
rect 17440 12030 17492 12036
rect 16336 11748 16388 11754
rect 16336 11690 16388 11696
rect 16428 11748 16480 11754
rect 16428 11690 16480 11696
rect 16980 11748 17032 11754
rect 16980 11690 17032 11696
rect 17452 11142 17480 12030
rect 17532 11748 17584 11754
rect 17532 11690 17584 11696
rect 17544 11210 17572 11690
rect 17636 11618 17664 12098
rect 17808 12020 17860 12026
rect 17808 11962 17860 11968
rect 17624 11612 17676 11618
rect 17676 11572 17756 11600
rect 17624 11554 17676 11560
rect 17532 11204 17584 11210
rect 17532 11146 17584 11152
rect 17624 11204 17676 11210
rect 17624 11146 17676 11152
rect 17440 11136 17492 11142
rect 17440 11078 17492 11084
rect 16060 10932 16112 10938
rect 16060 10874 16112 10880
rect 16072 10326 16100 10874
rect 17636 10598 17664 11146
rect 17728 11142 17756 11572
rect 17820 11142 17848 11962
rect 17716 11136 17768 11142
rect 17716 11078 17768 11084
rect 17808 11136 17860 11142
rect 17808 11078 17860 11084
rect 16244 10592 16296 10598
rect 16244 10534 16296 10540
rect 17624 10592 17676 10598
rect 17624 10534 17676 10540
rect 16060 10320 16112 10326
rect 16060 10262 16112 10268
rect 16072 10122 16100 10262
rect 16256 10122 16284 10534
rect 17728 10530 17756 11078
rect 17820 11006 17848 11078
rect 17808 11000 17860 11006
rect 17808 10942 17860 10948
rect 16336 10524 16388 10530
rect 16336 10466 16388 10472
rect 17716 10524 17768 10530
rect 17716 10466 17768 10472
rect 16060 10116 16112 10122
rect 16060 10058 16112 10064
rect 16244 10116 16296 10122
rect 16244 10058 16296 10064
rect 16348 10054 16376 10466
rect 16612 10320 16664 10326
rect 16612 10262 16664 10268
rect 17440 10320 17492 10326
rect 17440 10262 17492 10268
rect 16624 10122 16652 10262
rect 17452 10122 17480 10262
rect 16612 10116 16664 10122
rect 16612 10058 16664 10064
rect 17440 10116 17492 10122
rect 17912 10074 17940 14070
rect 18188 12638 18216 14186
rect 18280 13930 18308 15158
rect 18360 14944 18412 14950
rect 18360 14886 18412 14892
rect 18268 13924 18320 13930
rect 18268 13866 18320 13872
rect 18176 12632 18228 12638
rect 18176 12574 18228 12580
rect 18372 11550 18400 14886
rect 18464 14134 18492 15226
rect 18556 14950 18584 15362
rect 18648 15018 18676 15380
rect 18924 15358 18952 15702
rect 19016 15426 19044 15702
rect 19004 15420 19056 15426
rect 19004 15362 19056 15368
rect 18912 15352 18964 15358
rect 18740 15312 18912 15340
rect 18636 15012 18688 15018
rect 18636 14954 18688 14960
rect 18544 14944 18596 14950
rect 18544 14886 18596 14892
rect 18740 14474 18768 15312
rect 18912 15294 18964 15300
rect 18864 15116 19184 15136
rect 18864 15114 18876 15116
rect 18932 15114 18956 15116
rect 19012 15114 19036 15116
rect 19092 15114 19116 15116
rect 19172 15114 19184 15116
rect 18864 15062 18870 15114
rect 18932 15062 18934 15114
rect 19114 15062 19116 15114
rect 19178 15062 19184 15114
rect 18864 15060 18876 15062
rect 18932 15060 18956 15062
rect 19012 15060 19036 15062
rect 19092 15060 19116 15062
rect 19172 15060 19184 15062
rect 18864 15040 19184 15060
rect 19188 14672 19240 14678
rect 19188 14614 19240 14620
rect 18728 14468 18780 14474
rect 18728 14410 18780 14416
rect 19200 14338 19228 14614
rect 18544 14332 18596 14338
rect 18544 14274 18596 14280
rect 19188 14332 19240 14338
rect 19188 14274 19240 14280
rect 18452 14128 18504 14134
rect 18452 14070 18504 14076
rect 18452 13584 18504 13590
rect 18452 13526 18504 13532
rect 18464 13386 18492 13526
rect 18452 13380 18504 13386
rect 18452 13322 18504 13328
rect 18556 12774 18584 14274
rect 18864 14028 19184 14048
rect 18864 14026 18876 14028
rect 18932 14026 18956 14028
rect 19012 14026 19036 14028
rect 19092 14026 19116 14028
rect 19172 14026 19184 14028
rect 18864 13974 18870 14026
rect 18932 13974 18934 14026
rect 19114 13974 19116 14026
rect 19178 13974 19184 14026
rect 18864 13972 18876 13974
rect 18932 13972 18956 13974
rect 19012 13972 19036 13974
rect 19092 13972 19116 13974
rect 19172 13972 19184 13974
rect 18864 13952 19184 13972
rect 19384 13862 19412 16382
rect 19464 16372 19516 16378
rect 19464 16314 19516 16320
rect 19476 15970 19504 16314
rect 19464 15964 19516 15970
rect 19464 15906 19516 15912
rect 19464 14264 19516 14270
rect 19568 14252 19596 17062
rect 19844 16446 19872 17878
rect 19936 17670 19964 19782
rect 20292 19704 20344 19710
rect 20292 19646 20344 19652
rect 20200 19568 20252 19574
rect 20200 19510 20252 19516
rect 20212 17738 20240 19510
rect 20304 19370 20332 19646
rect 20292 19364 20344 19370
rect 20292 19306 20344 19312
rect 20672 19234 20700 22230
rect 21500 21886 21528 23318
rect 21592 22974 21620 23522
rect 21672 23376 21724 23382
rect 21672 23318 21724 23324
rect 21684 23178 21712 23318
rect 21672 23172 21724 23178
rect 21672 23114 21724 23120
rect 21580 22968 21632 22974
rect 21580 22910 21632 22916
rect 21776 22616 21804 31662
rect 23052 30108 23104 30114
rect 23052 30050 23104 30056
rect 23064 29706 23092 30050
rect 23248 29706 23276 31664
rect 24444 31662 24564 31690
rect 24678 31664 24790 32088
rect 23604 30040 23656 30046
rect 23604 29982 23656 29988
rect 23420 29972 23472 29978
rect 23420 29914 23472 29920
rect 23052 29700 23104 29706
rect 23052 29642 23104 29648
rect 23236 29700 23288 29706
rect 23236 29642 23288 29648
rect 23064 28482 23092 29642
rect 23432 29094 23460 29914
rect 23616 29706 23644 29982
rect 23788 29904 23840 29910
rect 23788 29846 23840 29852
rect 23604 29700 23656 29706
rect 23604 29642 23656 29648
rect 23800 29394 23828 29846
rect 24156 29700 24208 29706
rect 24156 29642 24208 29648
rect 24168 29502 24196 29642
rect 24156 29496 24208 29502
rect 24156 29438 24208 29444
rect 23880 29428 23932 29434
rect 23800 29376 23880 29394
rect 23800 29370 23932 29376
rect 23800 29366 23920 29370
rect 23696 29360 23748 29366
rect 23696 29302 23748 29308
rect 23420 29088 23472 29094
rect 23420 29030 23472 29036
rect 23512 29020 23564 29026
rect 23512 28962 23564 28968
rect 23524 28618 23552 28962
rect 23512 28612 23564 28618
rect 23512 28554 23564 28560
rect 21856 28476 21908 28482
rect 21856 28418 21908 28424
rect 23052 28476 23104 28482
rect 23052 28418 23104 28424
rect 21868 26850 21896 28418
rect 23708 28414 23736 29302
rect 24168 29162 24196 29438
rect 24156 29156 24208 29162
rect 24156 29098 24208 29104
rect 23696 28408 23748 28414
rect 23696 28350 23748 28356
rect 22500 28340 22552 28346
rect 22500 28282 22552 28288
rect 23052 28340 23104 28346
rect 23052 28282 23104 28288
rect 22512 27938 22540 28282
rect 23064 28074 23092 28282
rect 23052 28068 23104 28074
rect 23052 28010 23104 28016
rect 22408 27932 22460 27938
rect 22408 27874 22460 27880
rect 22500 27932 22552 27938
rect 22500 27874 22552 27880
rect 22224 27864 22276 27870
rect 22224 27806 22276 27812
rect 22236 27190 22264 27806
rect 22420 27258 22448 27874
rect 22960 27388 23012 27394
rect 23064 27376 23092 28010
rect 24340 27932 24392 27938
rect 24340 27874 24392 27880
rect 23512 27796 23564 27802
rect 23512 27738 23564 27744
rect 23012 27348 23092 27376
rect 22960 27330 23012 27336
rect 22408 27252 22460 27258
rect 22408 27194 22460 27200
rect 23328 27252 23380 27258
rect 23328 27194 23380 27200
rect 22224 27184 22276 27190
rect 22224 27126 22276 27132
rect 22236 26986 22264 27126
rect 22224 26980 22276 26986
rect 22224 26922 22276 26928
rect 21856 26844 21908 26850
rect 21856 26786 21908 26792
rect 21868 26442 21896 26786
rect 21856 26436 21908 26442
rect 21856 26378 21908 26384
rect 22500 25824 22552 25830
rect 22500 25766 22552 25772
rect 21856 25688 21908 25694
rect 21856 25630 21908 25636
rect 22224 25688 22276 25694
rect 22224 25630 22276 25636
rect 21868 25082 21896 25630
rect 22236 25354 22264 25630
rect 22512 25354 22540 25766
rect 23236 25688 23288 25694
rect 23236 25630 23288 25636
rect 22224 25348 22276 25354
rect 22224 25290 22276 25296
rect 22500 25348 22552 25354
rect 22500 25290 22552 25296
rect 21856 25076 21908 25082
rect 21856 25018 21908 25024
rect 21684 22588 21804 22616
rect 21488 21880 21540 21886
rect 21488 21822 21540 21828
rect 21396 20384 21448 20390
rect 21396 20326 21448 20332
rect 21028 20316 21080 20322
rect 21028 20258 21080 20264
rect 20752 20112 20804 20118
rect 20752 20054 20804 20060
rect 20764 19778 20792 20054
rect 20752 19772 20804 19778
rect 20752 19714 20804 19720
rect 20764 19370 20792 19714
rect 20752 19364 20804 19370
rect 20752 19306 20804 19312
rect 20660 19228 20712 19234
rect 20660 19170 20712 19176
rect 21040 19030 21068 20258
rect 21212 19840 21264 19846
rect 21212 19782 21264 19788
rect 21224 19710 21252 19782
rect 21212 19704 21264 19710
rect 21212 19646 21264 19652
rect 21408 19370 21436 20326
rect 21684 20322 21712 22588
rect 21868 22566 21896 25018
rect 22592 25008 22644 25014
rect 22592 24950 22644 24956
rect 21948 23988 22000 23994
rect 21948 23930 22000 23936
rect 21856 22560 21908 22566
rect 21856 22502 21908 22508
rect 21764 22492 21816 22498
rect 21764 22434 21816 22440
rect 21776 22090 21804 22434
rect 21868 22090 21896 22502
rect 21764 22084 21816 22090
rect 21764 22026 21816 22032
rect 21856 22084 21908 22090
rect 21856 22026 21908 22032
rect 21776 20390 21804 22026
rect 21960 21478 21988 23930
rect 21948 21472 22000 21478
rect 21948 21414 22000 21420
rect 21960 21002 21988 21414
rect 22604 21410 22632 24950
rect 22960 24600 23012 24606
rect 22960 24542 23012 24548
rect 22972 24198 23000 24542
rect 22960 24192 23012 24198
rect 22960 24134 23012 24140
rect 22972 23874 23000 24134
rect 22880 23846 23000 23874
rect 22880 23518 22908 23846
rect 22960 23580 23012 23586
rect 22960 23522 23012 23528
rect 22868 23512 22920 23518
rect 22868 23454 22920 23460
rect 22684 22968 22736 22974
rect 22684 22910 22736 22916
rect 22696 22498 22724 22910
rect 22880 22838 22908 23454
rect 22972 23042 23000 23522
rect 23144 23376 23196 23382
rect 23144 23318 23196 23324
rect 22960 23036 23012 23042
rect 22960 22978 23012 22984
rect 23156 22974 23184 23318
rect 23144 22968 23196 22974
rect 23144 22910 23196 22916
rect 22868 22832 22920 22838
rect 22868 22774 22920 22780
rect 22684 22492 22736 22498
rect 22684 22434 22736 22440
rect 22696 22022 22724 22434
rect 22684 22016 22736 22022
rect 22684 21958 22736 21964
rect 22776 21948 22828 21954
rect 22776 21890 22828 21896
rect 22132 21404 22184 21410
rect 22132 21346 22184 21352
rect 22316 21404 22368 21410
rect 22316 21346 22368 21352
rect 22592 21404 22644 21410
rect 22592 21346 22644 21352
rect 22144 21002 22172 21346
rect 21948 20996 22000 21002
rect 21948 20938 22000 20944
rect 22132 20996 22184 21002
rect 22132 20938 22184 20944
rect 22328 20730 22356 21346
rect 22604 20934 22632 21346
rect 22788 21206 22816 21890
rect 22880 21342 22908 22774
rect 23248 22566 23276 25630
rect 23340 25354 23368 27194
rect 23328 25348 23380 25354
rect 23328 25290 23380 25296
rect 23420 24464 23472 24470
rect 23420 24406 23472 24412
rect 23236 22560 23288 22566
rect 23156 22520 23236 22548
rect 22960 22492 23012 22498
rect 22960 22434 23012 22440
rect 22972 21886 23000 22434
rect 23156 21954 23184 22520
rect 23236 22502 23288 22508
rect 23236 22424 23288 22430
rect 23236 22366 23288 22372
rect 23144 21948 23196 21954
rect 23144 21890 23196 21896
rect 22960 21880 23012 21886
rect 22960 21822 23012 21828
rect 23248 21750 23276 22366
rect 23236 21744 23288 21750
rect 23236 21686 23288 21692
rect 23248 21410 23276 21686
rect 23432 21546 23460 24406
rect 23420 21540 23472 21546
rect 23420 21482 23472 21488
rect 23236 21404 23288 21410
rect 23236 21346 23288 21352
rect 22868 21336 22920 21342
rect 22868 21278 22920 21284
rect 22776 21200 22828 21206
rect 22776 21142 22828 21148
rect 22788 20934 22816 21142
rect 22592 20928 22644 20934
rect 22592 20870 22644 20876
rect 22776 20928 22828 20934
rect 22776 20870 22828 20876
rect 22880 20798 22908 21278
rect 23248 20866 23276 21346
rect 23432 21002 23460 21482
rect 23420 20996 23472 21002
rect 23420 20938 23472 20944
rect 23236 20860 23288 20866
rect 23236 20802 23288 20808
rect 22868 20792 22920 20798
rect 22868 20734 22920 20740
rect 22316 20724 22368 20730
rect 22316 20666 22368 20672
rect 22132 20656 22184 20662
rect 22132 20598 22184 20604
rect 21764 20384 21816 20390
rect 21764 20326 21816 20332
rect 21856 20384 21908 20390
rect 21856 20326 21908 20332
rect 21672 20316 21724 20322
rect 21672 20258 21724 20264
rect 21684 19846 21712 20258
rect 21868 19914 21896 20326
rect 22040 20248 22092 20254
rect 22040 20190 22092 20196
rect 21856 19908 21908 19914
rect 21856 19850 21908 19856
rect 21672 19840 21724 19846
rect 21672 19782 21724 19788
rect 21396 19364 21448 19370
rect 21396 19306 21448 19312
rect 21028 19024 21080 19030
rect 21028 18966 21080 18972
rect 20752 18072 20804 18078
rect 20752 18014 20804 18020
rect 20764 17738 20792 18014
rect 20936 17936 20988 17942
rect 20936 17878 20988 17884
rect 20200 17732 20252 17738
rect 20200 17674 20252 17680
rect 20752 17732 20804 17738
rect 20752 17674 20804 17680
rect 20844 17732 20896 17738
rect 20844 17674 20896 17680
rect 19924 17664 19976 17670
rect 19924 17606 19976 17612
rect 19936 16990 19964 17606
rect 20108 17460 20160 17466
rect 20108 17402 20160 17408
rect 20120 17058 20148 17402
rect 20200 17392 20252 17398
rect 20200 17334 20252 17340
rect 20108 17052 20160 17058
rect 20108 16994 20160 17000
rect 19924 16984 19976 16990
rect 19924 16926 19976 16932
rect 19832 16440 19884 16446
rect 19832 16382 19884 16388
rect 19844 15902 19872 16382
rect 19832 15896 19884 15902
rect 19832 15838 19884 15844
rect 20212 15204 20240 17334
rect 20764 17194 20792 17674
rect 20856 17534 20884 17674
rect 20948 17534 20976 17878
rect 20844 17528 20896 17534
rect 20844 17470 20896 17476
rect 20936 17528 20988 17534
rect 20936 17470 20988 17476
rect 20752 17188 20804 17194
rect 20752 17130 20804 17136
rect 20476 16984 20528 16990
rect 20476 16926 20528 16932
rect 20292 16916 20344 16922
rect 20292 16858 20344 16864
rect 20304 16650 20332 16858
rect 20292 16644 20344 16650
rect 20292 16586 20344 16592
rect 20488 16310 20516 16926
rect 20764 16650 20792 17130
rect 20936 17052 20988 17058
rect 20936 16994 20988 17000
rect 20752 16644 20804 16650
rect 20752 16586 20804 16592
rect 20948 16582 20976 16994
rect 20936 16576 20988 16582
rect 20936 16518 20988 16524
rect 20476 16304 20528 16310
rect 20476 16246 20528 16252
rect 20292 15216 20344 15222
rect 20212 15176 20292 15204
rect 20292 15158 20344 15164
rect 20108 15012 20160 15018
rect 20108 14954 20160 14960
rect 20016 14332 20068 14338
rect 20016 14274 20068 14280
rect 19516 14224 19596 14252
rect 19464 14206 19516 14212
rect 19372 13856 19424 13862
rect 19372 13798 19424 13804
rect 18636 13788 18688 13794
rect 18636 13730 18688 13736
rect 18728 13788 18780 13794
rect 18728 13730 18780 13736
rect 18648 13386 18676 13730
rect 18636 13380 18688 13386
rect 18636 13322 18688 13328
rect 18544 12768 18596 12774
rect 18544 12710 18596 12716
rect 18452 12496 18504 12502
rect 18452 12438 18504 12444
rect 18464 12298 18492 12438
rect 18452 12292 18504 12298
rect 18452 12234 18504 12240
rect 18556 12230 18584 12710
rect 18648 12280 18676 13322
rect 18740 13318 18768 13730
rect 19384 13386 19412 13798
rect 19568 13590 19596 14224
rect 20028 13794 20056 14274
rect 20120 14270 20148 14954
rect 20108 14264 20160 14270
rect 20108 14206 20160 14212
rect 20108 13924 20160 13930
rect 20108 13866 20160 13872
rect 20016 13788 20068 13794
rect 20016 13730 20068 13736
rect 19556 13584 19608 13590
rect 19556 13526 19608 13532
rect 19740 13584 19792 13590
rect 19740 13526 19792 13532
rect 19372 13380 19424 13386
rect 19372 13322 19424 13328
rect 18728 13312 18780 13318
rect 18728 13254 18780 13260
rect 19372 13244 19424 13250
rect 19372 13186 19424 13192
rect 18864 12940 19184 12960
rect 18864 12938 18876 12940
rect 18932 12938 18956 12940
rect 19012 12938 19036 12940
rect 19092 12938 19116 12940
rect 19172 12938 19184 12940
rect 18864 12886 18870 12938
rect 18932 12886 18934 12938
rect 19114 12886 19116 12938
rect 19178 12886 19184 12938
rect 18864 12884 18876 12886
rect 18932 12884 18956 12886
rect 19012 12884 19036 12886
rect 19092 12884 19116 12886
rect 19172 12884 19184 12886
rect 18864 12864 19184 12884
rect 18820 12700 18872 12706
rect 18820 12642 18872 12648
rect 18728 12292 18780 12298
rect 18648 12252 18728 12280
rect 18728 12234 18780 12240
rect 18544 12224 18596 12230
rect 18544 12166 18596 12172
rect 18740 11754 18768 12234
rect 18832 12094 18860 12642
rect 18820 12088 18872 12094
rect 18820 12030 18872 12036
rect 18864 11852 19184 11872
rect 18864 11850 18876 11852
rect 18932 11850 18956 11852
rect 19012 11850 19036 11852
rect 19092 11850 19116 11852
rect 19172 11850 19184 11852
rect 18864 11798 18870 11850
rect 18932 11798 18934 11850
rect 19114 11798 19116 11850
rect 19178 11798 19184 11850
rect 18864 11796 18876 11798
rect 18932 11796 18956 11798
rect 19012 11796 19036 11798
rect 19092 11796 19116 11798
rect 19172 11796 19184 11798
rect 18864 11776 19184 11796
rect 18728 11748 18780 11754
rect 18728 11690 18780 11696
rect 19280 11680 19332 11686
rect 19280 11622 19332 11628
rect 18360 11544 18412 11550
rect 18360 11486 18412 11492
rect 18728 10932 18780 10938
rect 18728 10874 18780 10880
rect 18452 10660 18504 10666
rect 18452 10602 18504 10608
rect 18464 10462 18492 10602
rect 18636 10524 18688 10530
rect 18636 10466 18688 10472
rect 18740 10512 18768 10874
rect 18864 10764 19184 10784
rect 18864 10762 18876 10764
rect 18932 10762 18956 10764
rect 19012 10762 19036 10764
rect 19092 10762 19116 10764
rect 19172 10762 19184 10764
rect 18864 10710 18870 10762
rect 18932 10710 18934 10762
rect 19114 10710 19116 10762
rect 19178 10710 19184 10762
rect 18864 10708 18876 10710
rect 18932 10708 18956 10710
rect 19012 10708 19036 10710
rect 19092 10708 19116 10710
rect 19172 10708 19184 10710
rect 18864 10688 19184 10708
rect 19292 10666 19320 11622
rect 19280 10660 19332 10666
rect 19108 10620 19280 10648
rect 18820 10524 18872 10530
rect 18740 10484 18820 10512
rect 18452 10456 18504 10462
rect 18452 10398 18504 10404
rect 18360 10320 18412 10326
rect 18360 10262 18412 10268
rect 18372 10122 18400 10262
rect 17440 10058 17492 10064
rect 16336 10048 16388 10054
rect 16336 9990 16388 9996
rect 15876 9912 15928 9918
rect 15876 9854 15928 9860
rect 15968 9912 16020 9918
rect 15968 9854 16020 9860
rect 15980 9442 16008 9854
rect 17348 9504 17400 9510
rect 17348 9446 17400 9452
rect 15968 9436 16020 9442
rect 15968 9378 16020 9384
rect 15980 9034 16008 9378
rect 16152 9232 16204 9238
rect 16152 9174 16204 9180
rect 16164 9034 16192 9174
rect 15692 9028 15744 9034
rect 15692 8970 15744 8976
rect 15968 9028 16020 9034
rect 15968 8970 16020 8976
rect 16152 9028 16204 9034
rect 16152 8970 16204 8976
rect 15784 7804 15836 7810
rect 15784 7746 15836 7752
rect 15416 6580 15468 6586
rect 15336 6540 15416 6568
rect 15232 6308 15284 6314
rect 15232 6250 15284 6256
rect 15140 5424 15192 5430
rect 15140 5366 15192 5372
rect 15152 4886 15180 5366
rect 15336 5072 15364 6540
rect 15416 6522 15468 6528
rect 15796 5770 15824 7746
rect 16164 6178 16192 8970
rect 17360 8762 17388 9446
rect 17452 8830 17480 10058
rect 17532 10048 17584 10054
rect 17532 9990 17584 9996
rect 17728 10046 17940 10074
rect 18360 10116 18412 10122
rect 18360 10058 18412 10064
rect 17544 9238 17572 9990
rect 17532 9232 17584 9238
rect 17532 9174 17584 9180
rect 17440 8824 17492 8830
rect 17440 8766 17492 8772
rect 17348 8756 17400 8762
rect 17348 8698 17400 8704
rect 17452 7946 17480 8766
rect 17544 8422 17572 9174
rect 17532 8416 17584 8422
rect 17532 8358 17584 8364
rect 17440 7940 17492 7946
rect 17440 7882 17492 7888
rect 16796 7600 16848 7606
rect 16796 7542 16848 7548
rect 16336 6512 16388 6518
rect 16336 6454 16388 6460
rect 15968 6172 16020 6178
rect 15968 6114 16020 6120
rect 16152 6172 16204 6178
rect 16152 6114 16204 6120
rect 15980 5770 16008 6114
rect 16244 6104 16296 6110
rect 16244 6046 16296 6052
rect 15784 5764 15836 5770
rect 15784 5706 15836 5712
rect 15968 5764 16020 5770
rect 15968 5706 16020 5712
rect 15796 5566 15824 5706
rect 15784 5560 15836 5566
rect 15784 5502 15836 5508
rect 16256 5430 16284 6046
rect 16348 5673 16376 6454
rect 16334 5664 16390 5673
rect 16334 5599 16390 5608
rect 15416 5424 15468 5430
rect 15416 5366 15468 5372
rect 16244 5424 16296 5430
rect 16244 5366 16296 5372
rect 15428 5090 15456 5366
rect 15244 5044 15364 5072
rect 15416 5084 15468 5090
rect 15140 4880 15192 4886
rect 15140 4822 15192 4828
rect 15244 4614 15272 5044
rect 15416 5026 15468 5032
rect 15876 5084 15928 5090
rect 15876 5026 15928 5032
rect 15324 4948 15376 4954
rect 15324 4890 15376 4896
rect 15336 4682 15364 4890
rect 15324 4676 15376 4682
rect 15324 4618 15376 4624
rect 15232 4608 15284 4614
rect 15232 4550 15284 4556
rect 15048 4336 15100 4342
rect 15048 4278 15100 4284
rect 14956 3996 15008 4002
rect 14956 3938 15008 3944
rect 14496 3860 14548 3866
rect 14496 3802 14548 3808
rect 14968 3594 14996 3938
rect 14956 3588 15008 3594
rect 14956 3530 15008 3536
rect 14404 3384 14456 3390
rect 14404 3326 14456 3332
rect 14772 3384 14824 3390
rect 14772 3326 14824 3332
rect 14784 3050 14812 3326
rect 15060 3322 15088 4278
rect 15428 4138 15456 5026
rect 15888 4682 15916 5026
rect 15876 4676 15928 4682
rect 15876 4618 15928 4624
rect 15692 4472 15744 4478
rect 15692 4414 15744 4420
rect 16060 4472 16112 4478
rect 16060 4414 16112 4420
rect 15416 4132 15468 4138
rect 15416 4074 15468 4080
rect 15428 3526 15456 4074
rect 15704 3934 15732 4414
rect 15692 3928 15744 3934
rect 15692 3870 15744 3876
rect 16072 3866 16100 4414
rect 16060 3860 16112 3866
rect 16060 3802 16112 3808
rect 16072 3594 16100 3802
rect 15508 3588 15560 3594
rect 15508 3530 15560 3536
rect 16060 3588 16112 3594
rect 16060 3530 16112 3536
rect 15416 3520 15468 3526
rect 15416 3462 15468 3468
rect 15048 3316 15100 3322
rect 15048 3258 15100 3264
rect 14772 3044 14824 3050
rect 14772 2986 14824 2992
rect 15520 2982 15548 3530
rect 15692 3384 15744 3390
rect 15692 3326 15744 3332
rect 15508 2976 15560 2982
rect 15508 2918 15560 2924
rect 15520 2506 15548 2918
rect 15704 2914 15732 3326
rect 16256 2914 16284 5366
rect 16348 5090 16376 5599
rect 16336 5084 16388 5090
rect 16336 5026 16388 5032
rect 16348 4342 16376 5026
rect 16336 4336 16388 4342
rect 16336 4278 16388 4284
rect 16808 4070 16836 7542
rect 16888 5152 16940 5158
rect 16888 5094 16940 5100
rect 17624 5152 17676 5158
rect 17624 5094 17676 5100
rect 16900 4682 16928 5094
rect 17072 5016 17124 5022
rect 17072 4958 17124 4964
rect 16888 4676 16940 4682
rect 16888 4618 16940 4624
rect 16796 4064 16848 4070
rect 16796 4006 16848 4012
rect 16808 3594 16836 4006
rect 16796 3588 16848 3594
rect 16796 3530 16848 3536
rect 16980 3384 17032 3390
rect 16980 3326 17032 3332
rect 15692 2908 15744 2914
rect 15692 2850 15744 2856
rect 16244 2908 16296 2914
rect 16244 2850 16296 2856
rect 16888 2908 16940 2914
rect 16888 2850 16940 2856
rect 15508 2500 15560 2506
rect 15508 2442 15560 2448
rect 15704 2234 15732 2850
rect 16060 2840 16112 2846
rect 16060 2782 16112 2788
rect 16072 2506 16100 2782
rect 16060 2500 16112 2506
rect 16060 2442 16112 2448
rect 16900 2370 16928 2850
rect 16888 2364 16940 2370
rect 16888 2306 16940 2312
rect 15692 2228 15744 2234
rect 15692 2170 15744 2176
rect 16992 1962 17020 3326
rect 17084 2982 17112 4958
rect 17636 4614 17664 5094
rect 17624 4608 17676 4614
rect 17624 4550 17676 4556
rect 17348 4064 17400 4070
rect 17348 4006 17400 4012
rect 17360 3254 17388 4006
rect 17532 3860 17584 3866
rect 17532 3802 17584 3808
rect 17544 3254 17572 3802
rect 17348 3248 17400 3254
rect 17348 3190 17400 3196
rect 17532 3248 17584 3254
rect 17532 3190 17584 3196
rect 17072 2976 17124 2982
rect 17072 2918 17124 2924
rect 17084 2438 17112 2918
rect 17164 2908 17216 2914
rect 17164 2850 17216 2856
rect 17176 2506 17204 2850
rect 17164 2500 17216 2506
rect 17164 2442 17216 2448
rect 17072 2432 17124 2438
rect 17072 2374 17124 2380
rect 16980 1956 17032 1962
rect 16980 1898 17032 1904
rect 17360 1758 17388 3190
rect 17544 2166 17572 3190
rect 17532 2160 17584 2166
rect 17532 2102 17584 2108
rect 17348 1752 17400 1758
rect 17348 1694 17400 1700
rect 15140 1616 15192 1622
rect 15140 1558 15192 1564
rect 16612 1616 16664 1622
rect 16612 1558 16664 1564
rect 15152 1078 15180 1558
rect 16624 1078 16652 1558
rect 15140 1072 15192 1078
rect 15140 1014 15192 1020
rect 15508 1072 15560 1078
rect 15508 1014 15560 1020
rect 16612 1072 16664 1078
rect 16612 1014 16664 1020
rect 15520 424 15548 1014
rect 16624 426 16652 1014
rect 17728 777 17756 10046
rect 18360 9776 18412 9782
rect 18464 9764 18492 10398
rect 18412 9736 18492 9764
rect 18360 9718 18412 9724
rect 18266 9472 18322 9481
rect 17992 9436 18044 9442
rect 18266 9407 18322 9416
rect 17992 9378 18044 9384
rect 18004 8898 18032 9378
rect 18084 9368 18136 9374
rect 18084 9310 18136 9316
rect 17992 8892 18044 8898
rect 17992 8834 18044 8840
rect 17808 8756 17860 8762
rect 17808 8698 17860 8704
rect 17820 8257 17848 8698
rect 18004 8490 18032 8834
rect 18096 8762 18124 9310
rect 18280 8966 18308 9407
rect 18268 8960 18320 8966
rect 18268 8902 18320 8908
rect 18084 8756 18136 8762
rect 18084 8698 18136 8704
rect 17992 8484 18044 8490
rect 17992 8426 18044 8432
rect 17806 8248 17862 8257
rect 17806 8183 17862 8192
rect 17820 7266 17848 8183
rect 18004 7946 18032 8426
rect 17992 7940 18044 7946
rect 17992 7882 18044 7888
rect 17808 7260 17860 7266
rect 17808 7202 17860 7208
rect 18176 7260 18228 7266
rect 18176 7202 18228 7208
rect 17820 6790 17848 7202
rect 18188 6858 18216 7202
rect 18176 6852 18228 6858
rect 18176 6794 18228 6800
rect 17808 6784 17860 6790
rect 17808 6726 17860 6732
rect 18268 6648 18320 6654
rect 18268 6590 18320 6596
rect 18280 6178 18308 6590
rect 18268 6172 18320 6178
rect 18268 6114 18320 6120
rect 18280 5770 18308 6114
rect 18268 5764 18320 5770
rect 18268 5706 18320 5712
rect 18372 5650 18400 9718
rect 18648 9578 18676 10466
rect 18740 9578 18768 10484
rect 18820 10466 18872 10472
rect 18912 10456 18964 10462
rect 18912 10398 18964 10404
rect 18924 9850 18952 10398
rect 19108 9918 19136 10620
rect 19280 10602 19332 10608
rect 19280 9980 19332 9986
rect 19280 9922 19332 9928
rect 19096 9912 19148 9918
rect 19096 9854 19148 9860
rect 18912 9844 18964 9850
rect 18912 9786 18964 9792
rect 18864 9676 19184 9696
rect 18864 9674 18876 9676
rect 18932 9674 18956 9676
rect 19012 9674 19036 9676
rect 19092 9674 19116 9676
rect 19172 9674 19184 9676
rect 18864 9622 18870 9674
rect 18932 9622 18934 9674
rect 19114 9622 19116 9674
rect 19178 9622 19184 9674
rect 18864 9620 18876 9622
rect 18932 9620 18956 9622
rect 19012 9620 19036 9622
rect 19092 9620 19116 9622
rect 19172 9620 19184 9622
rect 18864 9600 19184 9620
rect 19292 9578 19320 9922
rect 18636 9572 18688 9578
rect 18636 9514 18688 9520
rect 18728 9572 18780 9578
rect 18728 9514 18780 9520
rect 19280 9572 19332 9578
rect 19280 9514 19332 9520
rect 18450 9472 18506 9481
rect 19384 9442 19412 13186
rect 19752 13182 19780 13526
rect 19740 13176 19792 13182
rect 19740 13118 19792 13124
rect 19752 13046 19780 13118
rect 19464 13040 19516 13046
rect 19464 12982 19516 12988
rect 19740 13040 19792 13046
rect 19740 12982 19792 12988
rect 19476 12502 19504 12982
rect 19556 12632 19608 12638
rect 19556 12574 19608 12580
rect 19464 12496 19516 12502
rect 19464 12438 19516 12444
rect 19464 11952 19516 11958
rect 19464 11894 19516 11900
rect 19476 10462 19504 11894
rect 19464 10456 19516 10462
rect 19464 10398 19516 10404
rect 19464 9912 19516 9918
rect 19464 9854 19516 9860
rect 18450 9407 18506 9416
rect 19372 9436 19424 9442
rect 18464 9374 18492 9407
rect 19372 9378 19424 9384
rect 18452 9368 18504 9374
rect 18452 9310 18504 9316
rect 18464 9034 18492 9310
rect 19384 9034 19412 9378
rect 18452 9028 18504 9034
rect 18452 8970 18504 8976
rect 19372 9028 19424 9034
rect 19372 8970 19424 8976
rect 18728 8824 18780 8830
rect 18728 8766 18780 8772
rect 18740 7334 18768 8766
rect 18864 8588 19184 8608
rect 18864 8586 18876 8588
rect 18932 8586 18956 8588
rect 19012 8586 19036 8588
rect 19092 8586 19116 8588
rect 19172 8586 19184 8588
rect 18864 8534 18870 8586
rect 18932 8534 18934 8586
rect 19114 8534 19116 8586
rect 19178 8534 19184 8586
rect 18864 8532 18876 8534
rect 18932 8532 18956 8534
rect 19012 8532 19036 8534
rect 19092 8532 19116 8534
rect 19172 8532 19184 8534
rect 18864 8512 19184 8532
rect 18864 7500 19184 7520
rect 18864 7498 18876 7500
rect 18932 7498 18956 7500
rect 19012 7498 19036 7500
rect 19092 7498 19116 7500
rect 19172 7498 19184 7500
rect 18864 7446 18870 7498
rect 18932 7446 18934 7498
rect 19114 7446 19116 7498
rect 19178 7446 19184 7498
rect 18864 7444 18876 7446
rect 18932 7444 18956 7446
rect 19012 7444 19036 7446
rect 19092 7444 19116 7446
rect 19172 7444 19184 7446
rect 18864 7424 19184 7444
rect 18728 7328 18780 7334
rect 18728 7270 18780 7276
rect 18452 7260 18504 7266
rect 18452 7202 18504 7208
rect 18464 6518 18492 7202
rect 18740 6858 18768 7270
rect 18728 6852 18780 6858
rect 18728 6794 18780 6800
rect 18452 6512 18504 6518
rect 18452 6454 18504 6460
rect 18280 5622 18400 5650
rect 18280 4886 18308 5622
rect 18360 5084 18412 5090
rect 18360 5026 18412 5032
rect 18268 4880 18320 4886
rect 18268 4822 18320 4828
rect 18176 4608 18228 4614
rect 18176 4550 18228 4556
rect 18188 4138 18216 4550
rect 18372 4478 18400 5026
rect 18360 4472 18412 4478
rect 18360 4414 18412 4420
rect 18176 4132 18228 4138
rect 18176 4074 18228 4080
rect 17900 3996 17952 4002
rect 17900 3938 17952 3944
rect 17808 3928 17860 3934
rect 17808 3870 17860 3876
rect 17820 3526 17848 3870
rect 17808 3520 17860 3526
rect 17808 3462 17860 3468
rect 17820 3050 17848 3462
rect 17912 3390 17940 3938
rect 17900 3384 17952 3390
rect 17900 3326 17952 3332
rect 17808 3044 17860 3050
rect 17808 2986 17860 2992
rect 17912 2982 17940 3326
rect 18188 3050 18216 4074
rect 18372 4070 18400 4414
rect 18360 4064 18412 4070
rect 18360 4006 18412 4012
rect 18464 3594 18492 6454
rect 18864 6412 19184 6432
rect 18864 6410 18876 6412
rect 18932 6410 18956 6412
rect 19012 6410 19036 6412
rect 19092 6410 19116 6412
rect 19172 6410 19184 6412
rect 18864 6358 18870 6410
rect 18932 6358 18934 6410
rect 19114 6358 19116 6410
rect 19178 6358 19184 6410
rect 18864 6356 18876 6358
rect 18932 6356 18956 6358
rect 19012 6356 19036 6358
rect 19092 6356 19116 6358
rect 19172 6356 19184 6358
rect 18864 6336 19184 6356
rect 19476 6178 19504 9854
rect 19464 6172 19516 6178
rect 19464 6114 19516 6120
rect 18636 5968 18688 5974
rect 18636 5910 18688 5916
rect 18648 5430 18676 5910
rect 19372 5628 19424 5634
rect 19372 5570 19424 5576
rect 19464 5628 19516 5634
rect 19464 5570 19516 5576
rect 18636 5424 18688 5430
rect 18636 5366 18688 5372
rect 19280 5424 19332 5430
rect 19384 5401 19412 5570
rect 19280 5366 19332 5372
rect 19370 5392 19426 5401
rect 18648 5022 18676 5366
rect 18864 5324 19184 5344
rect 18864 5322 18876 5324
rect 18932 5322 18956 5324
rect 19012 5322 19036 5324
rect 19092 5322 19116 5324
rect 19172 5322 19184 5324
rect 18864 5270 18870 5322
rect 18932 5270 18934 5322
rect 19114 5270 19116 5322
rect 19178 5270 19184 5322
rect 18864 5268 18876 5270
rect 18932 5268 18956 5270
rect 19012 5268 19036 5270
rect 19092 5268 19116 5270
rect 19172 5268 19184 5270
rect 18864 5248 19184 5268
rect 18544 5016 18596 5022
rect 18544 4958 18596 4964
rect 18636 5016 18688 5022
rect 18636 4958 18688 4964
rect 18556 4614 18584 4958
rect 18648 4682 18676 4958
rect 18636 4676 18688 4682
rect 18636 4618 18688 4624
rect 18728 4676 18780 4682
rect 18728 4618 18780 4624
rect 18544 4608 18596 4614
rect 18544 4550 18596 4556
rect 18634 4576 18690 4585
rect 18634 4511 18690 4520
rect 18648 4478 18676 4511
rect 18636 4472 18688 4478
rect 18636 4414 18688 4420
rect 18452 3588 18504 3594
rect 18452 3530 18504 3536
rect 18636 3452 18688 3458
rect 18740 3440 18768 4618
rect 19292 4585 19320 5366
rect 19370 5327 19426 5336
rect 19278 4576 19334 4585
rect 19476 4554 19504 5570
rect 19278 4511 19334 4520
rect 19384 4526 19504 4554
rect 18864 4236 19184 4256
rect 18864 4234 18876 4236
rect 18932 4234 18956 4236
rect 19012 4234 19036 4236
rect 19092 4234 19116 4236
rect 19172 4234 19184 4236
rect 18864 4182 18870 4234
rect 18932 4182 18934 4234
rect 19114 4182 19116 4234
rect 19178 4182 19184 4234
rect 18864 4180 18876 4182
rect 18932 4180 18956 4182
rect 19012 4180 19036 4182
rect 19092 4180 19116 4182
rect 19172 4180 19184 4182
rect 18864 4160 19184 4180
rect 19188 3860 19240 3866
rect 19188 3802 19240 3808
rect 18912 3792 18964 3798
rect 18912 3734 18964 3740
rect 18924 3594 18952 3734
rect 18912 3588 18964 3594
rect 18912 3530 18964 3536
rect 19200 3458 19228 3802
rect 18688 3412 18768 3440
rect 19188 3452 19240 3458
rect 18636 3394 18688 3400
rect 19188 3394 19240 3400
rect 19280 3384 19332 3390
rect 19280 3326 19332 3332
rect 18636 3316 18688 3322
rect 18636 3258 18688 3264
rect 18176 3044 18228 3050
rect 18176 2986 18228 2992
rect 17900 2976 17952 2982
rect 17900 2918 17952 2924
rect 18648 2710 18676 3258
rect 18864 3148 19184 3168
rect 18864 3146 18876 3148
rect 18932 3146 18956 3148
rect 19012 3146 19036 3148
rect 19092 3146 19116 3148
rect 19172 3146 19184 3148
rect 18864 3094 18870 3146
rect 18932 3094 18934 3146
rect 19114 3094 19116 3146
rect 19178 3094 19184 3146
rect 18864 3092 18876 3094
rect 18932 3092 18956 3094
rect 19012 3092 19036 3094
rect 19092 3092 19116 3094
rect 19172 3092 19184 3094
rect 18864 3072 19184 3092
rect 18452 2704 18504 2710
rect 18452 2646 18504 2652
rect 18636 2704 18688 2710
rect 18636 2646 18688 2652
rect 19096 2704 19148 2710
rect 19096 2646 19148 2652
rect 18360 2364 18412 2370
rect 18360 2306 18412 2312
rect 18176 2228 18228 2234
rect 18228 2188 18308 2216
rect 18176 2170 18228 2176
rect 18176 1752 18228 1758
rect 18176 1694 18228 1700
rect 18188 1418 18216 1694
rect 18176 1412 18228 1418
rect 18176 1354 18228 1360
rect 17714 768 17770 777
rect 17714 703 17770 712
rect 16624 424 17020 426
rect 18280 424 18308 2188
rect 18372 1962 18400 2306
rect 18464 2302 18492 2646
rect 18452 2296 18504 2302
rect 18452 2238 18504 2244
rect 18544 2296 18596 2302
rect 18544 2238 18596 2244
rect 18464 1962 18492 2238
rect 18360 1956 18412 1962
rect 18360 1898 18412 1904
rect 18452 1956 18504 1962
rect 18452 1898 18504 1904
rect 18372 1350 18400 1898
rect 18452 1820 18504 1826
rect 18452 1762 18504 1768
rect 18464 1418 18492 1762
rect 18556 1690 18584 2238
rect 18648 1894 18676 2646
rect 19108 2302 19136 2646
rect 19096 2296 19148 2302
rect 19096 2238 19148 2244
rect 18864 2060 19184 2080
rect 18864 2058 18876 2060
rect 18932 2058 18956 2060
rect 19012 2058 19036 2060
rect 19092 2058 19116 2060
rect 19172 2058 19184 2060
rect 18864 2006 18870 2058
rect 18932 2006 18934 2058
rect 19114 2006 19116 2058
rect 19178 2006 19184 2058
rect 18864 2004 18876 2006
rect 18932 2004 18956 2006
rect 19012 2004 19036 2006
rect 19092 2004 19116 2006
rect 19172 2004 19184 2006
rect 18864 1984 19184 2004
rect 18636 1888 18688 1894
rect 18636 1830 18688 1836
rect 18728 1820 18780 1826
rect 18728 1762 18780 1768
rect 19096 1820 19148 1826
rect 19096 1762 19148 1768
rect 18544 1684 18596 1690
rect 18544 1626 18596 1632
rect 18740 1418 18768 1762
rect 18452 1412 18504 1418
rect 18452 1354 18504 1360
rect 18728 1412 18780 1418
rect 18728 1354 18780 1360
rect 18360 1344 18412 1350
rect 18360 1286 18412 1292
rect 19108 1282 19136 1762
rect 19096 1276 19148 1282
rect 19096 1218 19148 1224
rect 19292 1146 19320 3326
rect 19384 2506 19412 4526
rect 19372 2500 19424 2506
rect 19372 2442 19424 2448
rect 19384 2234 19412 2442
rect 19372 2228 19424 2234
rect 19372 2170 19424 2176
rect 19464 2160 19516 2166
rect 19464 2102 19516 2108
rect 19476 1758 19504 2102
rect 19464 1752 19516 1758
rect 19464 1694 19516 1700
rect 19280 1140 19332 1146
rect 19280 1082 19332 1088
rect 18864 972 19184 992
rect 18864 970 18876 972
rect 18932 970 18956 972
rect 19012 970 19036 972
rect 19092 970 19116 972
rect 19172 970 19184 972
rect 18864 918 18870 970
rect 18932 918 18934 970
rect 19114 918 19116 970
rect 19178 918 19184 970
rect 18864 916 18876 918
rect 18932 916 18956 918
rect 19012 916 19036 918
rect 19092 916 19116 918
rect 19172 916 19184 918
rect 18864 896 19184 916
rect 19568 777 19596 12574
rect 19924 10864 19976 10870
rect 19924 10806 19976 10812
rect 19936 10122 19964 10806
rect 19924 10116 19976 10122
rect 19924 10058 19976 10064
rect 19936 9850 19964 10058
rect 19924 9844 19976 9850
rect 19924 9786 19976 9792
rect 20028 7044 20056 13730
rect 20120 13386 20148 13866
rect 20108 13380 20160 13386
rect 20108 13322 20160 13328
rect 20108 11952 20160 11958
rect 20108 11894 20160 11900
rect 20120 11754 20148 11894
rect 20108 11748 20160 11754
rect 20108 11690 20160 11696
rect 20120 10394 20148 11690
rect 20304 10870 20332 15158
rect 20292 10864 20344 10870
rect 20292 10806 20344 10812
rect 20108 10388 20160 10394
rect 20108 10330 20160 10336
rect 20384 9980 20436 9986
rect 20384 9922 20436 9928
rect 20396 9889 20424 9922
rect 20382 9880 20438 9889
rect 20382 9815 20438 9824
rect 20200 7056 20252 7062
rect 20028 7016 20200 7044
rect 20200 6998 20252 7004
rect 20212 6722 20240 6998
rect 20200 6716 20252 6722
rect 20200 6658 20252 6664
rect 19832 6172 19884 6178
rect 19832 6114 19884 6120
rect 19844 5770 19872 6114
rect 20212 6042 20240 6658
rect 20384 6512 20436 6518
rect 20384 6454 20436 6460
rect 20396 6110 20424 6454
rect 20384 6104 20436 6110
rect 20384 6046 20436 6052
rect 20200 6036 20252 6042
rect 20200 5978 20252 5984
rect 19832 5764 19884 5770
rect 19832 5706 19884 5712
rect 19844 5090 19872 5706
rect 20396 5702 20424 6046
rect 20384 5696 20436 5702
rect 20384 5638 20436 5644
rect 19832 5084 19884 5090
rect 19832 5026 19884 5032
rect 20488 3934 20516 16246
rect 20568 15420 20620 15426
rect 20568 15362 20620 15368
rect 20580 14270 20608 15362
rect 20568 14264 20620 14270
rect 20568 14206 20620 14212
rect 21040 13930 21068 18966
rect 21120 18208 21172 18214
rect 21120 18150 21172 18156
rect 21132 17398 21160 18150
rect 21684 18078 21712 19782
rect 22052 19642 22080 20190
rect 22040 19636 22092 19642
rect 22040 19578 22092 19584
rect 22040 19228 22092 19234
rect 22040 19170 22092 19176
rect 22052 18622 22080 19170
rect 22144 19166 22172 20598
rect 22132 19160 22184 19166
rect 22132 19102 22184 19108
rect 22040 18616 22092 18622
rect 22040 18558 22092 18564
rect 21672 18072 21724 18078
rect 21672 18014 21724 18020
rect 21684 17670 21712 18014
rect 21672 17664 21724 17670
rect 21672 17606 21724 17612
rect 21396 17460 21448 17466
rect 21396 17402 21448 17408
rect 21120 17392 21172 17398
rect 21120 17334 21172 17340
rect 21408 17058 21436 17402
rect 21396 17052 21448 17058
rect 21396 16994 21448 17000
rect 21408 16650 21436 16994
rect 21684 16990 21712 17606
rect 21856 17392 21908 17398
rect 21856 17334 21908 17340
rect 21672 16984 21724 16990
rect 21672 16926 21724 16932
rect 21396 16644 21448 16650
rect 21396 16586 21448 16592
rect 21580 16372 21632 16378
rect 21580 16314 21632 16320
rect 21028 13924 21080 13930
rect 21028 13866 21080 13872
rect 20752 13176 20804 13182
rect 20752 13118 20804 13124
rect 20568 12496 20620 12502
rect 20568 12438 20620 12444
rect 20580 12065 20608 12438
rect 20764 12094 20792 13118
rect 21028 12224 21080 12230
rect 21028 12166 21080 12172
rect 20752 12088 20804 12094
rect 20566 12056 20622 12065
rect 20752 12030 20804 12036
rect 20566 11991 20622 12000
rect 20660 12020 20712 12026
rect 20580 11958 20608 11991
rect 20660 11962 20712 11968
rect 20568 11952 20620 11958
rect 20568 11894 20620 11900
rect 20672 11618 20700 11962
rect 20660 11612 20712 11618
rect 20660 11554 20712 11560
rect 20660 11476 20712 11482
rect 20764 11464 20792 12030
rect 20712 11436 20792 11464
rect 20660 11418 20712 11424
rect 20672 11385 20700 11418
rect 20658 11376 20714 11385
rect 20658 11311 20714 11320
rect 20658 9880 20714 9889
rect 20658 9815 20714 9824
rect 20672 9209 20700 9815
rect 20658 9200 20714 9209
rect 20658 9135 20714 9144
rect 20936 8348 20988 8354
rect 20936 8290 20988 8296
rect 20568 8212 20620 8218
rect 20568 8154 20620 8160
rect 20580 7606 20608 8154
rect 20948 7878 20976 8290
rect 20936 7872 20988 7878
rect 20764 7832 20936 7860
rect 20568 7600 20620 7606
rect 20568 7542 20620 7548
rect 20580 7305 20608 7542
rect 20566 7296 20622 7305
rect 20566 7231 20622 7240
rect 20568 6580 20620 6586
rect 20568 6522 20620 6528
rect 20580 6178 20608 6522
rect 20568 6172 20620 6178
rect 20568 6114 20620 6120
rect 20580 5770 20608 6114
rect 20568 5764 20620 5770
rect 20568 5706 20620 5712
rect 20660 5628 20712 5634
rect 20660 5570 20712 5576
rect 20672 5430 20700 5570
rect 20660 5424 20712 5430
rect 20660 5366 20712 5372
rect 20672 5158 20700 5366
rect 20764 5226 20792 7832
rect 20936 7814 20988 7820
rect 20936 7056 20988 7062
rect 20936 6998 20988 7004
rect 20948 6654 20976 6998
rect 20936 6648 20988 6654
rect 20936 6590 20988 6596
rect 20936 5424 20988 5430
rect 20936 5366 20988 5372
rect 20948 5226 20976 5366
rect 20752 5220 20804 5226
rect 20752 5162 20804 5168
rect 20936 5220 20988 5226
rect 20936 5162 20988 5168
rect 20660 5152 20712 5158
rect 20660 5094 20712 5100
rect 20672 4614 20700 5094
rect 20660 4608 20712 4614
rect 20660 4550 20712 4556
rect 21040 4554 21068 12166
rect 21304 12088 21356 12094
rect 21304 12030 21356 12036
rect 21316 11754 21344 12030
rect 21304 11748 21356 11754
rect 21304 11690 21356 11696
rect 21304 11612 21356 11618
rect 21304 11554 21356 11560
rect 21316 11210 21344 11554
rect 21488 11544 21540 11550
rect 21488 11486 21540 11492
rect 21500 11210 21528 11486
rect 21304 11204 21356 11210
rect 21304 11146 21356 11152
rect 21488 11204 21540 11210
rect 21488 11146 21540 11152
rect 21488 9776 21540 9782
rect 21488 9718 21540 9724
rect 21212 8824 21264 8830
rect 21212 8766 21264 8772
rect 21224 8354 21252 8766
rect 21212 8348 21264 8354
rect 21212 8290 21264 8296
rect 21224 7946 21252 8290
rect 21212 7940 21264 7946
rect 21212 7882 21264 7888
rect 21120 6648 21172 6654
rect 21120 6590 21172 6596
rect 21132 5770 21160 6590
rect 21120 5764 21172 5770
rect 21120 5706 21172 5712
rect 21132 5158 21160 5706
rect 21212 5560 21264 5566
rect 21212 5502 21264 5508
rect 21120 5152 21172 5158
rect 21120 5094 21172 5100
rect 21224 4886 21252 5502
rect 21396 5084 21448 5090
rect 21396 5026 21448 5032
rect 21212 4880 21264 4886
rect 21212 4822 21264 4828
rect 21212 4676 21264 4682
rect 21212 4618 21264 4624
rect 20948 4526 21068 4554
rect 21120 4540 21172 4546
rect 20568 4404 20620 4410
rect 20568 4346 20620 4352
rect 20476 3928 20528 3934
rect 20476 3870 20528 3876
rect 20488 3769 20516 3870
rect 19646 3760 19702 3769
rect 19646 3695 19702 3704
rect 20474 3760 20530 3769
rect 20474 3695 20530 3704
rect 19660 1282 19688 3695
rect 20200 3588 20252 3594
rect 20200 3530 20252 3536
rect 19740 2704 19792 2710
rect 19740 2646 19792 2652
rect 19648 1276 19700 1282
rect 19648 1218 19700 1224
rect 19660 806 19688 1218
rect 19648 800 19700 806
rect 19554 768 19610 777
rect 19648 742 19700 748
rect 19554 703 19610 712
rect 19752 424 19780 2646
rect 20212 1826 20240 3530
rect 20200 1820 20252 1826
rect 20200 1762 20252 1768
rect 20212 1214 20240 1762
rect 20200 1208 20252 1214
rect 20200 1150 20252 1156
rect 20212 874 20240 1150
rect 20200 868 20252 874
rect 20200 810 20252 816
rect 20580 505 20608 4346
rect 20752 2160 20804 2166
rect 20752 2102 20804 2108
rect 20660 1752 20712 1758
rect 20660 1694 20712 1700
rect 20672 1418 20700 1694
rect 20660 1412 20712 1418
rect 20660 1354 20712 1360
rect 20764 505 20792 2102
rect 20948 641 20976 4526
rect 21120 4482 21172 4488
rect 21028 4336 21080 4342
rect 21028 4278 21080 4284
rect 21040 3866 21068 4278
rect 21028 3860 21080 3866
rect 21028 3802 21080 3808
rect 21040 3594 21068 3802
rect 21028 3588 21080 3594
rect 21028 3530 21080 3536
rect 21040 2370 21068 3530
rect 21132 2914 21160 4482
rect 21224 3526 21252 4618
rect 21408 4546 21436 5026
rect 21500 4585 21528 9718
rect 21592 8218 21620 16314
rect 21868 15902 21896 17334
rect 21856 15896 21908 15902
rect 21856 15838 21908 15844
rect 21868 15766 21896 15838
rect 21856 15760 21908 15766
rect 21856 15702 21908 15708
rect 21672 13924 21724 13930
rect 21672 13866 21724 13872
rect 21684 13386 21712 13866
rect 21856 13720 21908 13726
rect 21856 13662 21908 13668
rect 21672 13380 21724 13386
rect 21672 13322 21724 13328
rect 21868 13182 21896 13662
rect 21856 13176 21908 13182
rect 21856 13118 21908 13124
rect 21672 13040 21724 13046
rect 21672 12982 21724 12988
rect 21684 12094 21712 12982
rect 21948 12700 22000 12706
rect 21948 12642 22000 12648
rect 21764 12496 21816 12502
rect 21764 12438 21816 12444
rect 21672 12088 21724 12094
rect 21672 12030 21724 12036
rect 21776 12026 21804 12438
rect 21960 12298 21988 12642
rect 21948 12292 22000 12298
rect 21948 12234 22000 12240
rect 21856 12088 21908 12094
rect 21856 12030 21908 12036
rect 21764 12020 21816 12026
rect 21764 11962 21816 11968
rect 21672 11680 21724 11686
rect 21672 11622 21724 11628
rect 21684 10870 21712 11622
rect 21672 10864 21724 10870
rect 21672 10806 21724 10812
rect 21776 8762 21804 11962
rect 21868 11142 21896 12030
rect 21856 11136 21908 11142
rect 21856 11078 21908 11084
rect 21960 10938 21988 12234
rect 21948 10932 22000 10938
rect 21948 10874 22000 10880
rect 21764 8756 21816 8762
rect 21764 8698 21816 8704
rect 21764 8348 21816 8354
rect 21764 8290 21816 8296
rect 21580 8212 21632 8218
rect 21580 8154 21632 8160
rect 21592 7946 21620 8154
rect 21580 7940 21632 7946
rect 21580 7882 21632 7888
rect 21776 7742 21804 8290
rect 22052 8286 22080 18558
rect 22144 18486 22172 19102
rect 22132 18480 22184 18486
rect 22132 18422 22184 18428
rect 22144 17738 22172 18422
rect 22132 17732 22184 17738
rect 22132 17674 22184 17680
rect 22132 16100 22184 16106
rect 22132 16042 22184 16048
rect 22144 15562 22172 16042
rect 22328 15970 22356 20666
rect 23248 20322 23276 20802
rect 23420 20792 23472 20798
rect 23420 20734 23472 20740
rect 23432 20458 23460 20734
rect 23420 20452 23472 20458
rect 23420 20394 23472 20400
rect 23236 20316 23288 20322
rect 23236 20258 23288 20264
rect 23432 19370 23460 20394
rect 23420 19364 23472 19370
rect 23420 19306 23472 19312
rect 23236 19228 23288 19234
rect 23236 19170 23288 19176
rect 23248 18826 23276 19170
rect 23236 18820 23288 18826
rect 23236 18762 23288 18768
rect 22500 17528 22552 17534
rect 22500 17470 22552 17476
rect 22512 16990 22540 17470
rect 22592 17460 22644 17466
rect 22592 17402 22644 17408
rect 22500 16984 22552 16990
rect 22500 16926 22552 16932
rect 22512 16650 22540 16926
rect 22500 16644 22552 16650
rect 22500 16586 22552 16592
rect 22604 16038 22632 17402
rect 22960 17052 23012 17058
rect 22960 16994 23012 17000
rect 22972 16378 23000 16994
rect 23144 16984 23196 16990
rect 23144 16926 23196 16932
rect 23156 16446 23184 16926
rect 23248 16922 23276 18762
rect 23432 18758 23460 19306
rect 23524 18826 23552 27738
rect 24352 27530 24380 27874
rect 24340 27524 24392 27530
rect 24340 27466 24392 27472
rect 24444 27410 24472 31662
rect 24536 31626 24564 31662
rect 24720 31626 24748 31664
rect 24536 31598 24748 31626
rect 25640 31662 25852 31690
rect 25966 31664 26078 32088
rect 27438 31664 27550 32088
rect 28726 31664 28838 32088
rect 30198 31690 30310 32088
rect 29504 31664 30310 31690
rect 31486 31664 31598 32088
rect 24524 30108 24576 30114
rect 24524 30050 24576 30056
rect 24616 30108 24668 30114
rect 24616 30050 24668 30056
rect 24536 29570 24564 30050
rect 24524 29564 24576 29570
rect 24524 29506 24576 29512
rect 24524 29428 24576 29434
rect 24524 29370 24576 29376
rect 24536 28618 24564 29370
rect 24628 28958 24656 30050
rect 25350 29464 25406 29473
rect 24892 29428 24944 29434
rect 25350 29399 25406 29408
rect 24892 29370 24944 29376
rect 24904 29162 24932 29370
rect 24892 29156 24944 29162
rect 24892 29098 24944 29104
rect 24616 28952 24668 28958
rect 24616 28894 24668 28900
rect 24524 28612 24576 28618
rect 24524 28554 24576 28560
rect 24628 28550 24656 28894
rect 24616 28544 24668 28550
rect 24616 28486 24668 28492
rect 24984 28408 25036 28414
rect 24984 28350 25036 28356
rect 24996 28074 25024 28350
rect 24984 28068 25036 28074
rect 24984 28010 25036 28016
rect 24616 28000 24668 28006
rect 24616 27942 24668 27948
rect 24352 27382 24472 27410
rect 23696 27252 23748 27258
rect 23696 27194 23748 27200
rect 23708 26986 23736 27194
rect 23696 26980 23748 26986
rect 23696 26922 23748 26928
rect 24248 26164 24300 26170
rect 24248 26106 24300 26112
rect 24260 23722 24288 26106
rect 24248 23716 24300 23722
rect 24248 23658 24300 23664
rect 24260 23178 24288 23658
rect 24248 23172 24300 23178
rect 24248 23114 24300 23120
rect 24156 23104 24208 23110
rect 24156 23046 24208 23052
rect 23972 22900 24024 22906
rect 23972 22842 24024 22848
rect 23984 22634 24012 22842
rect 23972 22628 24024 22634
rect 23972 22570 24024 22576
rect 24168 21410 24196 23046
rect 24156 21404 24208 21410
rect 24156 21346 24208 21352
rect 23788 21200 23840 21206
rect 23788 21142 23840 21148
rect 23800 20866 23828 21142
rect 24168 21002 24196 21346
rect 24156 20996 24208 21002
rect 24156 20938 24208 20944
rect 23788 20860 23840 20866
rect 23788 20802 23840 20808
rect 23604 20792 23656 20798
rect 23604 20734 23656 20740
rect 23616 20390 23644 20734
rect 23604 20384 23656 20390
rect 23604 20326 23656 20332
rect 24168 19914 24196 20938
rect 24156 19908 24208 19914
rect 24156 19850 24208 19856
rect 24156 19024 24208 19030
rect 24156 18966 24208 18972
rect 23512 18820 23564 18826
rect 23512 18762 23564 18768
rect 23420 18752 23472 18758
rect 23420 18694 23472 18700
rect 23420 17936 23472 17942
rect 23420 17878 23472 17884
rect 23432 17398 23460 17878
rect 23420 17392 23472 17398
rect 23420 17334 23472 17340
rect 23328 17052 23380 17058
rect 23328 16994 23380 17000
rect 23236 16916 23288 16922
rect 23236 16858 23288 16864
rect 23248 16650 23276 16858
rect 23236 16644 23288 16650
rect 23236 16586 23288 16592
rect 23340 16514 23368 16994
rect 23524 16582 23552 18762
rect 24168 18690 24196 18966
rect 24156 18684 24208 18690
rect 24156 18626 24208 18632
rect 23788 18616 23840 18622
rect 23788 18558 23840 18564
rect 23696 18480 23748 18486
rect 23696 18422 23748 18428
rect 23708 17466 23736 18422
rect 23800 17942 23828 18558
rect 23788 17936 23840 17942
rect 23788 17878 23840 17884
rect 23972 17936 24024 17942
rect 23972 17878 24024 17884
rect 23880 17732 23932 17738
rect 23880 17674 23932 17680
rect 23696 17460 23748 17466
rect 23696 17402 23748 17408
rect 23604 17392 23656 17398
rect 23604 17334 23656 17340
rect 23512 16576 23564 16582
rect 23512 16518 23564 16524
rect 23328 16508 23380 16514
rect 23328 16450 23380 16456
rect 23144 16440 23196 16446
rect 23144 16382 23196 16388
rect 22960 16372 23012 16378
rect 22960 16314 23012 16320
rect 22592 16032 22644 16038
rect 22592 15974 22644 15980
rect 22316 15964 22368 15970
rect 22316 15906 22368 15912
rect 22224 15896 22276 15902
rect 22224 15838 22276 15844
rect 22132 15556 22184 15562
rect 22132 15498 22184 15504
rect 22236 15222 22264 15838
rect 22408 15760 22460 15766
rect 22408 15702 22460 15708
rect 22420 15562 22448 15702
rect 22316 15556 22368 15562
rect 22316 15498 22368 15504
rect 22408 15556 22460 15562
rect 22408 15498 22460 15504
rect 22224 15216 22276 15222
rect 22224 15158 22276 15164
rect 22236 13930 22264 15158
rect 22224 13924 22276 13930
rect 22224 13866 22276 13872
rect 22132 13788 22184 13794
rect 22132 13730 22184 13736
rect 22144 13386 22172 13730
rect 22328 13726 22356 15498
rect 22604 15290 22632 15974
rect 23616 15494 23644 17334
rect 23892 15970 23920 17674
rect 23984 17602 24012 17878
rect 23972 17596 24024 17602
rect 23972 17538 24024 17544
rect 24064 16848 24116 16854
rect 24064 16790 24116 16796
rect 24076 16582 24104 16790
rect 24168 16650 24196 18626
rect 24248 17936 24300 17942
rect 24248 17878 24300 17884
rect 24260 17602 24288 17878
rect 24248 17596 24300 17602
rect 24248 17538 24300 17544
rect 24156 16644 24208 16650
rect 24156 16586 24208 16592
rect 24064 16576 24116 16582
rect 24064 16518 24116 16524
rect 24076 16106 24104 16518
rect 24156 16440 24208 16446
rect 24156 16382 24208 16388
rect 24064 16100 24116 16106
rect 24064 16042 24116 16048
rect 23880 15964 23932 15970
rect 23880 15906 23932 15912
rect 24064 15760 24116 15766
rect 24064 15702 24116 15708
rect 23604 15488 23656 15494
rect 23604 15430 23656 15436
rect 22592 15284 22644 15290
rect 22592 15226 22644 15232
rect 23420 14876 23472 14882
rect 23420 14818 23472 14824
rect 22408 14196 22460 14202
rect 22408 14138 22460 14144
rect 22420 13794 22448 14138
rect 23432 14134 23460 14818
rect 23420 14128 23472 14134
rect 23420 14070 23472 14076
rect 23432 13794 23460 14070
rect 22408 13788 22460 13794
rect 22408 13730 22460 13736
rect 23420 13788 23472 13794
rect 23420 13730 23472 13736
rect 22316 13720 22368 13726
rect 22316 13662 22368 13668
rect 22132 13380 22184 13386
rect 22132 13322 22184 13328
rect 22328 13318 22356 13662
rect 22316 13312 22368 13318
rect 22316 13254 22368 13260
rect 22420 13114 22448 13730
rect 23432 13386 23460 13730
rect 23420 13380 23472 13386
rect 23420 13322 23472 13328
rect 22408 13108 22460 13114
rect 22408 13050 22460 13056
rect 23050 12736 23106 12745
rect 23432 12706 23460 13322
rect 23972 13040 24024 13046
rect 23972 12982 24024 12988
rect 23050 12671 23106 12680
rect 23420 12700 23472 12706
rect 23064 12094 23092 12671
rect 23420 12642 23472 12648
rect 23144 12564 23196 12570
rect 23144 12506 23196 12512
rect 23156 12230 23184 12506
rect 23880 12496 23932 12502
rect 23880 12438 23932 12444
rect 23144 12224 23196 12230
rect 23144 12166 23196 12172
rect 23052 12088 23104 12094
rect 23052 12030 23104 12036
rect 23064 11754 23092 12030
rect 23156 11754 23184 12166
rect 23236 12156 23288 12162
rect 23236 12098 23288 12104
rect 23248 11958 23276 12098
rect 23892 12094 23920 12438
rect 23512 12088 23564 12094
rect 23512 12030 23564 12036
rect 23880 12088 23932 12094
rect 23880 12030 23932 12036
rect 23236 11952 23288 11958
rect 23236 11894 23288 11900
rect 23052 11748 23104 11754
rect 23052 11690 23104 11696
rect 23144 11748 23196 11754
rect 23144 11690 23196 11696
rect 22500 11544 22552 11550
rect 22500 11486 22552 11492
rect 22512 9442 22540 11486
rect 23248 10870 23276 11894
rect 23524 11550 23552 12030
rect 23892 11754 23920 12030
rect 23880 11748 23932 11754
rect 23880 11690 23932 11696
rect 23512 11544 23564 11550
rect 23512 11486 23564 11492
rect 23984 10977 24012 12982
rect 24076 11686 24104 15702
rect 24168 15358 24196 16382
rect 24260 15562 24288 17538
rect 24248 15556 24300 15562
rect 24248 15498 24300 15504
rect 24156 15352 24208 15358
rect 24156 15294 24208 15300
rect 24168 14678 24196 15294
rect 24248 14808 24300 14814
rect 24248 14750 24300 14756
rect 24156 14672 24208 14678
rect 24156 14614 24208 14620
rect 24168 13726 24196 14614
rect 24260 14134 24288 14750
rect 24352 14214 24380 27382
rect 24524 27184 24576 27190
rect 24524 27126 24576 27132
rect 24536 25762 24564 27126
rect 24628 26986 24656 27942
rect 24616 26980 24668 26986
rect 24616 26922 24668 26928
rect 24996 26442 25024 28010
rect 24984 26436 25036 26442
rect 24984 26378 25036 26384
rect 24892 25892 24944 25898
rect 24892 25834 24944 25840
rect 24524 25756 24576 25762
rect 24524 25698 24576 25704
rect 24432 25552 24484 25558
rect 24432 25494 24484 25500
rect 24444 25082 24472 25494
rect 24536 25354 24564 25698
rect 24524 25348 24576 25354
rect 24524 25290 24576 25296
rect 24904 25286 24932 25834
rect 24892 25280 24944 25286
rect 24892 25222 24944 25228
rect 24524 25144 24576 25150
rect 24524 25086 24576 25092
rect 24708 25144 24760 25150
rect 24708 25086 24760 25092
rect 24432 25076 24484 25082
rect 24432 25018 24484 25024
rect 24444 23042 24472 25018
rect 24536 23178 24564 25086
rect 24720 24810 24748 25086
rect 24708 24804 24760 24810
rect 24708 24746 24760 24752
rect 24800 23376 24852 23382
rect 24800 23318 24852 23324
rect 24524 23172 24576 23178
rect 24524 23114 24576 23120
rect 24432 23036 24484 23042
rect 24432 22978 24484 22984
rect 24444 22634 24472 22978
rect 24812 22974 24840 23318
rect 24616 22968 24668 22974
rect 24616 22910 24668 22916
rect 24800 22968 24852 22974
rect 24800 22910 24852 22916
rect 24432 22628 24484 22634
rect 24432 22570 24484 22576
rect 24524 21812 24576 21818
rect 24524 21754 24576 21760
rect 24536 21342 24564 21754
rect 24524 21336 24576 21342
rect 24524 21278 24576 21284
rect 24536 21002 24564 21278
rect 24524 20996 24576 21002
rect 24524 20938 24576 20944
rect 24628 20798 24656 22910
rect 24616 20792 24668 20798
rect 24616 20734 24668 20740
rect 24708 19024 24760 19030
rect 24708 18966 24760 18972
rect 24720 18554 24748 18966
rect 24708 18548 24760 18554
rect 24708 18490 24760 18496
rect 24720 17466 24748 18490
rect 24708 17460 24760 17466
rect 24708 17402 24760 17408
rect 24616 16440 24668 16446
rect 24616 16382 24668 16388
rect 24628 15834 24656 16382
rect 24616 15828 24668 15834
rect 24616 15770 24668 15776
rect 24708 15216 24760 15222
rect 24708 15158 24760 15164
rect 24352 14186 24472 14214
rect 24720 14202 24748 15158
rect 24248 14128 24300 14134
rect 24248 14070 24300 14076
rect 24156 13720 24208 13726
rect 24156 13662 24208 13668
rect 24168 13182 24196 13662
rect 24260 13386 24288 14070
rect 24248 13380 24300 13386
rect 24248 13322 24300 13328
rect 24156 13176 24208 13182
rect 24156 13118 24208 13124
rect 24168 12638 24196 13118
rect 24340 12700 24392 12706
rect 24340 12642 24392 12648
rect 24156 12632 24208 12638
rect 24156 12574 24208 12580
rect 24168 11754 24196 12574
rect 24248 12156 24300 12162
rect 24248 12098 24300 12104
rect 24260 12026 24288 12098
rect 24248 12020 24300 12026
rect 24248 11962 24300 11968
rect 24156 11748 24208 11754
rect 24156 11690 24208 11696
rect 24064 11680 24116 11686
rect 24064 11622 24116 11628
rect 23970 10968 24026 10977
rect 23970 10903 24026 10912
rect 23236 10864 23288 10870
rect 23236 10806 23288 10812
rect 22958 10560 23014 10569
rect 22958 10495 23014 10504
rect 22972 10462 23000 10495
rect 22960 10456 23012 10462
rect 22960 10398 23012 10404
rect 22972 9900 23000 10398
rect 23144 10320 23196 10326
rect 23144 10262 23196 10268
rect 23052 9912 23104 9918
rect 22972 9872 23052 9900
rect 23052 9854 23104 9860
rect 23156 9850 23184 10262
rect 22868 9844 22920 9850
rect 22868 9786 22920 9792
rect 23144 9844 23196 9850
rect 23144 9786 23196 9792
rect 22880 9442 22908 9786
rect 22500 9436 22552 9442
rect 22500 9378 22552 9384
rect 22868 9436 22920 9442
rect 22868 9378 22920 9384
rect 22512 8966 22540 9378
rect 22776 9368 22828 9374
rect 22776 9310 22828 9316
rect 22788 9034 22816 9310
rect 22880 9034 22908 9378
rect 23156 9345 23184 9786
rect 23248 9510 23276 10806
rect 23788 10456 23840 10462
rect 23788 10398 23840 10404
rect 23420 9912 23472 9918
rect 23420 9854 23472 9860
rect 23236 9504 23288 9510
rect 23288 9464 23368 9492
rect 23236 9446 23288 9452
rect 23142 9336 23198 9345
rect 23198 9294 23276 9322
rect 23142 9271 23198 9280
rect 22776 9028 22828 9034
rect 22776 8970 22828 8976
rect 22868 9028 22920 9034
rect 22868 8970 22920 8976
rect 22500 8960 22552 8966
rect 22500 8902 22552 8908
rect 22868 8348 22920 8354
rect 22868 8290 22920 8296
rect 22040 8280 22092 8286
rect 22040 8222 22092 8228
rect 22880 7878 22908 8290
rect 23052 8144 23104 8150
rect 23052 8086 23104 8092
rect 23064 7946 23092 8086
rect 23052 7940 23104 7946
rect 23052 7882 23104 7888
rect 22868 7872 22920 7878
rect 22868 7814 22920 7820
rect 21764 7736 21816 7742
rect 21764 7678 21816 7684
rect 23064 7266 23092 7882
rect 23248 7810 23276 9294
rect 23340 8898 23368 9464
rect 23328 8892 23380 8898
rect 23328 8834 23380 8840
rect 23236 7804 23288 7810
rect 23236 7746 23288 7752
rect 23248 7402 23276 7746
rect 23236 7396 23288 7402
rect 23236 7338 23288 7344
rect 23052 7260 23104 7266
rect 23052 7202 23104 7208
rect 23064 6858 23092 7202
rect 23052 6852 23104 6858
rect 23052 6794 23104 6800
rect 21948 6648 22000 6654
rect 21948 6590 22000 6596
rect 21672 6580 21724 6586
rect 21672 6522 21724 6528
rect 21580 6512 21632 6518
rect 21580 6454 21632 6460
rect 21592 6246 21620 6454
rect 21580 6240 21632 6246
rect 21580 6182 21632 6188
rect 21592 5702 21620 6182
rect 21684 5702 21712 6522
rect 21960 6110 21988 6590
rect 23340 6586 23368 8834
rect 23432 6654 23460 9854
rect 23696 9776 23748 9782
rect 23696 9718 23748 9724
rect 23512 8280 23564 8286
rect 23512 8222 23564 8228
rect 23524 7878 23552 8222
rect 23512 7872 23564 7878
rect 23512 7814 23564 7820
rect 23604 7668 23656 7674
rect 23604 7610 23656 7616
rect 23420 6648 23472 6654
rect 23420 6590 23472 6596
rect 23328 6580 23380 6586
rect 23328 6522 23380 6528
rect 23616 6518 23644 7610
rect 23708 7334 23736 9718
rect 23800 9220 23828 10398
rect 24076 9889 24104 11622
rect 24352 11414 24380 12642
rect 24340 11408 24392 11414
rect 24340 11350 24392 11356
rect 24352 10462 24380 11350
rect 24340 10456 24392 10462
rect 24340 10398 24392 10404
rect 24248 10388 24300 10394
rect 24248 10330 24300 10336
rect 24062 9880 24118 9889
rect 24062 9815 24118 9824
rect 23800 9192 23920 9220
rect 23786 8112 23842 8121
rect 23786 8047 23842 8056
rect 23800 7878 23828 8047
rect 23892 7985 23920 9192
rect 23878 7976 23934 7985
rect 23878 7911 23934 7920
rect 23972 7940 24024 7946
rect 23972 7882 24024 7888
rect 23788 7872 23840 7878
rect 23880 7872 23932 7878
rect 23840 7832 23880 7860
rect 23788 7814 23840 7820
rect 23880 7814 23932 7820
rect 23984 7674 24012 7882
rect 23972 7668 24024 7674
rect 23972 7610 24024 7616
rect 23696 7328 23748 7334
rect 23696 7270 23748 7276
rect 23708 6790 23736 7270
rect 23696 6784 23748 6790
rect 23696 6726 23748 6732
rect 24260 6654 24288 10330
rect 24338 9472 24394 9481
rect 24338 9407 24394 9416
rect 24352 8694 24380 9407
rect 24340 8688 24392 8694
rect 24340 8630 24392 8636
rect 24352 8354 24380 8630
rect 24340 8348 24392 8354
rect 24340 8290 24392 8296
rect 24340 7668 24392 7674
rect 24340 7610 24392 7616
rect 24352 7402 24380 7610
rect 24340 7396 24392 7402
rect 24340 7338 24392 7344
rect 24352 6654 24380 7338
rect 23696 6648 23748 6654
rect 23696 6590 23748 6596
rect 24248 6648 24300 6654
rect 24248 6590 24300 6596
rect 24340 6648 24392 6654
rect 24340 6590 24392 6596
rect 22132 6512 22184 6518
rect 22132 6454 22184 6460
rect 23604 6512 23656 6518
rect 23604 6454 23656 6460
rect 21948 6104 22000 6110
rect 21948 6046 22000 6052
rect 21856 5764 21908 5770
rect 21856 5706 21908 5712
rect 21580 5696 21632 5702
rect 21580 5638 21632 5644
rect 21672 5696 21724 5702
rect 21672 5638 21724 5644
rect 21684 5566 21712 5638
rect 21868 5566 21896 5706
rect 21672 5560 21724 5566
rect 21672 5502 21724 5508
rect 21856 5560 21908 5566
rect 21856 5502 21908 5508
rect 21486 4576 21542 4585
rect 21396 4540 21448 4546
rect 21486 4511 21542 4520
rect 21396 4482 21448 4488
rect 21580 4336 21632 4342
rect 21580 4278 21632 4284
rect 21488 3928 21540 3934
rect 21488 3870 21540 3876
rect 21304 3792 21356 3798
rect 21304 3734 21356 3740
rect 21316 3594 21344 3734
rect 21304 3588 21356 3594
rect 21304 3530 21356 3536
rect 21212 3520 21264 3526
rect 21212 3462 21264 3468
rect 21212 3044 21264 3050
rect 21212 2986 21264 2992
rect 21120 2908 21172 2914
rect 21120 2850 21172 2856
rect 21132 2438 21160 2850
rect 21224 2506 21252 2986
rect 21316 2982 21344 3530
rect 21500 3458 21528 3870
rect 21488 3452 21540 3458
rect 21488 3394 21540 3400
rect 21592 3050 21620 4278
rect 21684 4002 21712 5502
rect 21764 5152 21816 5158
rect 21764 5094 21816 5100
rect 21776 4682 21804 5094
rect 21764 4676 21816 4682
rect 21764 4618 21816 4624
rect 21868 4002 21896 5502
rect 22144 5158 22172 6454
rect 23420 5628 23472 5634
rect 23420 5570 23472 5576
rect 22222 5256 22278 5265
rect 22222 5191 22278 5200
rect 22132 5152 22184 5158
rect 22132 5094 22184 5100
rect 21672 3996 21724 4002
rect 21672 3938 21724 3944
rect 21856 3996 21908 4002
rect 21856 3938 21908 3944
rect 21684 3322 21712 3938
rect 21868 3594 21896 3938
rect 22236 3934 22264 5191
rect 23432 5158 23460 5570
rect 23420 5152 23472 5158
rect 23420 5094 23472 5100
rect 22224 3928 22276 3934
rect 22224 3870 22276 3876
rect 21856 3588 21908 3594
rect 21856 3530 21908 3536
rect 21868 3458 21896 3530
rect 21856 3452 21908 3458
rect 21856 3394 21908 3400
rect 21672 3316 21724 3322
rect 21672 3258 21724 3264
rect 22236 3050 22264 3870
rect 23144 3860 23196 3866
rect 23144 3802 23196 3808
rect 23156 3254 23184 3802
rect 23328 3792 23380 3798
rect 23328 3734 23380 3740
rect 23340 3594 23368 3734
rect 23328 3588 23380 3594
rect 23328 3530 23380 3536
rect 23144 3248 23196 3254
rect 23144 3190 23196 3196
rect 21580 3044 21632 3050
rect 21580 2986 21632 2992
rect 22224 3044 22276 3050
rect 22224 2986 22276 2992
rect 21304 2976 21356 2982
rect 21304 2918 21356 2924
rect 21316 2506 21344 2918
rect 21212 2500 21264 2506
rect 21212 2442 21264 2448
rect 21304 2500 21356 2506
rect 21304 2442 21356 2448
rect 21120 2432 21172 2438
rect 21120 2374 21172 2380
rect 21028 2364 21080 2370
rect 21028 2306 21080 2312
rect 21224 1894 21252 2442
rect 23156 2234 23184 3190
rect 23340 3050 23368 3530
rect 23418 3352 23474 3361
rect 23418 3287 23474 3296
rect 23432 3254 23460 3287
rect 23420 3248 23472 3254
rect 23420 3190 23472 3196
rect 23328 3044 23380 3050
rect 23328 2986 23380 2992
rect 23236 2500 23288 2506
rect 23236 2442 23288 2448
rect 23248 2250 23276 2442
rect 23340 2370 23368 2986
rect 23616 2710 23644 6454
rect 23708 2846 23736 6590
rect 24260 6314 24288 6590
rect 24248 6308 24300 6314
rect 24248 6250 24300 6256
rect 24248 5764 24300 5770
rect 24248 5706 24300 5712
rect 24260 5090 24288 5706
rect 24444 5158 24472 14186
rect 24708 14196 24760 14202
rect 24708 14138 24760 14144
rect 24720 13658 24748 14138
rect 24812 13930 24840 22910
rect 25168 21200 25220 21206
rect 25168 21142 25220 21148
rect 25180 19030 25208 21142
rect 25168 19024 25220 19030
rect 25168 18966 25220 18972
rect 25260 16440 25312 16446
rect 25260 16382 25312 16388
rect 25272 15358 25300 16382
rect 24892 15352 24944 15358
rect 24892 15294 24944 15300
rect 25260 15352 25312 15358
rect 25260 15294 25312 15300
rect 24800 13924 24852 13930
rect 24800 13866 24852 13872
rect 24708 13652 24760 13658
rect 24708 13594 24760 13600
rect 24720 12706 24748 13594
rect 24812 13386 24840 13866
rect 24800 13380 24852 13386
rect 24800 13322 24852 13328
rect 24708 12700 24760 12706
rect 24708 12642 24760 12648
rect 24720 12298 24748 12642
rect 24708 12292 24760 12298
rect 24708 12234 24760 12240
rect 24904 11006 24932 15294
rect 25260 14332 25312 14338
rect 25260 14274 25312 14280
rect 25272 12706 25300 14274
rect 25260 12700 25312 12706
rect 25260 12642 25312 12648
rect 25272 12162 25300 12642
rect 25260 12156 25312 12162
rect 25260 12098 25312 12104
rect 25364 11142 25392 29399
rect 25536 22288 25588 22294
rect 25536 22230 25588 22236
rect 25548 22022 25576 22230
rect 25536 22016 25588 22022
rect 25536 21958 25588 21964
rect 25640 19734 25668 31662
rect 25824 31626 25852 31662
rect 26008 31626 26036 31664
rect 25824 31598 26036 31626
rect 27480 30794 27508 31664
rect 27468 30788 27520 30794
rect 27468 30730 27520 30736
rect 26916 30584 26968 30590
rect 26916 30526 26968 30532
rect 25996 30040 26048 30046
rect 25996 29982 26048 29988
rect 26008 29366 26036 29982
rect 26928 29706 26956 30526
rect 27836 30108 27888 30114
rect 27836 30050 27888 30056
rect 27652 30040 27704 30046
rect 27652 29982 27704 29988
rect 26916 29700 26968 29706
rect 26916 29642 26968 29648
rect 26456 29564 26508 29570
rect 26456 29506 26508 29512
rect 26088 29428 26140 29434
rect 26088 29370 26140 29376
rect 25996 29360 26048 29366
rect 25996 29302 26048 29308
rect 26100 28346 26128 29370
rect 26180 28816 26232 28822
rect 26180 28758 26232 28764
rect 26192 28482 26220 28758
rect 26180 28476 26232 28482
rect 26180 28418 26232 28424
rect 26088 28340 26140 28346
rect 26088 28282 26140 28288
rect 25904 26844 25956 26850
rect 25904 26786 25956 26792
rect 25916 26102 25944 26786
rect 25904 26096 25956 26102
rect 25904 26038 25956 26044
rect 25916 25082 25944 26038
rect 25904 25076 25956 25082
rect 25904 25018 25956 25024
rect 25904 24668 25956 24674
rect 25904 24610 25956 24616
rect 25916 24266 25944 24610
rect 25904 24260 25956 24266
rect 25956 24220 26036 24248
rect 25904 24202 25956 24208
rect 25904 23988 25956 23994
rect 25904 23930 25956 23936
rect 25916 22362 25944 23930
rect 26008 22974 26036 24220
rect 26100 23874 26128 28282
rect 26192 26918 26220 28418
rect 26180 26912 26232 26918
rect 26180 26854 26232 26860
rect 26192 26442 26220 26854
rect 26180 26436 26232 26442
rect 26180 26378 26232 26384
rect 26192 25286 26220 26378
rect 26180 25280 26232 25286
rect 26232 25240 26312 25268
rect 26180 25222 26232 25228
rect 26180 25144 26232 25150
rect 26180 25086 26232 25092
rect 26192 24742 26220 25086
rect 26180 24736 26232 24742
rect 26180 24678 26232 24684
rect 26192 24266 26220 24678
rect 26284 24674 26312 25240
rect 26272 24668 26324 24674
rect 26272 24610 26324 24616
rect 26180 24260 26232 24266
rect 26180 24202 26232 24208
rect 26100 23846 26220 23874
rect 25996 22968 26048 22974
rect 25996 22910 26048 22916
rect 26192 22498 26220 23846
rect 26180 22492 26232 22498
rect 26180 22434 26232 22440
rect 25996 22424 26048 22430
rect 25996 22366 26048 22372
rect 25812 22356 25864 22362
rect 25812 22298 25864 22304
rect 25904 22356 25956 22362
rect 25904 22298 25956 22304
rect 25824 21342 25852 22298
rect 25916 22090 25944 22298
rect 25904 22084 25956 22090
rect 25904 22026 25956 22032
rect 26008 21750 26036 22366
rect 26192 22022 26220 22434
rect 26272 22288 26324 22294
rect 26272 22230 26324 22236
rect 26180 22016 26232 22022
rect 26180 21958 26232 21964
rect 25996 21744 26048 21750
rect 25996 21686 26048 21692
rect 25812 21336 25864 21342
rect 25812 21278 25864 21284
rect 26008 20730 26036 21686
rect 25996 20724 26048 20730
rect 25996 20666 26048 20672
rect 25548 19706 25668 19734
rect 25548 17602 25576 19706
rect 25904 18820 25956 18826
rect 25904 18762 25956 18768
rect 25536 17596 25588 17602
rect 25536 17538 25588 17544
rect 25444 16440 25496 16446
rect 25444 16382 25496 16388
rect 25456 16038 25484 16382
rect 25444 16032 25496 16038
rect 25444 15974 25496 15980
rect 25548 15426 25576 17538
rect 25916 17534 25944 18762
rect 25904 17528 25956 17534
rect 25904 17470 25956 17476
rect 26180 16508 26232 16514
rect 26180 16450 26232 16456
rect 26192 16378 26220 16450
rect 26180 16372 26232 16378
rect 26180 16314 26232 16320
rect 25812 15964 25864 15970
rect 25812 15906 25864 15912
rect 25536 15420 25588 15426
rect 25536 15362 25588 15368
rect 25548 15329 25576 15362
rect 25534 15320 25590 15329
rect 25534 15255 25590 15264
rect 25824 13794 25852 15906
rect 26088 15488 26140 15494
rect 26088 15430 26140 15436
rect 25996 14944 26048 14950
rect 25996 14886 26048 14892
rect 26008 14134 26036 14886
rect 26100 14474 26128 15430
rect 26192 15222 26220 16314
rect 26180 15216 26232 15222
rect 26180 15158 26232 15164
rect 26192 14814 26220 15158
rect 26284 14882 26312 22230
rect 26364 22016 26416 22022
rect 26364 21958 26416 21964
rect 26376 21886 26404 21958
rect 26468 21886 26496 29506
rect 27664 29434 27692 29982
rect 27848 29706 27876 30050
rect 27836 29700 27888 29706
rect 27756 29660 27836 29688
rect 26916 29428 26968 29434
rect 26916 29370 26968 29376
rect 27652 29428 27704 29434
rect 27652 29370 27704 29376
rect 26928 29026 26956 29370
rect 27664 29094 27692 29370
rect 27756 29366 27784 29660
rect 27836 29642 27888 29648
rect 27836 29496 27888 29502
rect 27836 29438 27888 29444
rect 27744 29360 27796 29366
rect 27744 29302 27796 29308
rect 27652 29088 27704 29094
rect 27652 29030 27704 29036
rect 26916 29020 26968 29026
rect 26916 28962 26968 28968
rect 26928 28550 26956 28962
rect 27192 28952 27244 28958
rect 27192 28894 27244 28900
rect 27284 28952 27336 28958
rect 27284 28894 27336 28900
rect 27204 28618 27232 28894
rect 27192 28612 27244 28618
rect 27192 28554 27244 28560
rect 26916 28544 26968 28550
rect 26916 28486 26968 28492
rect 27204 28006 27232 28554
rect 27296 28278 27324 28894
rect 27664 28618 27692 29030
rect 27652 28612 27704 28618
rect 27652 28554 27704 28560
rect 27284 28272 27336 28278
rect 27284 28214 27336 28220
rect 27192 28000 27244 28006
rect 27192 27942 27244 27948
rect 27204 27530 27232 27942
rect 27296 27938 27324 28214
rect 27848 28074 27876 29438
rect 28204 29428 28256 29434
rect 28204 29370 28256 29376
rect 28768 29394 28796 31664
rect 29504 31662 30268 31664
rect 28848 30516 28900 30522
rect 28848 30458 28900 30464
rect 28860 30250 28888 30458
rect 28848 30244 28900 30250
rect 28848 30186 28900 30192
rect 28860 29570 28888 30186
rect 29400 30040 29452 30046
rect 29400 29982 29452 29988
rect 28848 29564 28900 29570
rect 28848 29506 28900 29512
rect 29412 29434 29440 29982
rect 29400 29428 29452 29434
rect 28216 28618 28244 29370
rect 28768 29366 28980 29394
rect 29400 29370 29452 29376
rect 28480 29360 28532 29366
rect 28480 29302 28532 29308
rect 28204 28612 28256 28618
rect 28204 28554 28256 28560
rect 28112 28476 28164 28482
rect 28112 28418 28164 28424
rect 28020 28408 28072 28414
rect 28020 28350 28072 28356
rect 27836 28068 27888 28074
rect 27836 28010 27888 28016
rect 27284 27932 27336 27938
rect 27284 27874 27336 27880
rect 27192 27524 27244 27530
rect 27192 27466 27244 27472
rect 27296 27190 27324 27874
rect 27560 27864 27612 27870
rect 27560 27806 27612 27812
rect 27572 27530 27600 27806
rect 27560 27524 27612 27530
rect 27560 27466 27612 27472
rect 27284 27184 27336 27190
rect 27284 27126 27336 27132
rect 27100 26232 27152 26238
rect 27100 26174 27152 26180
rect 27112 25762 27140 26174
rect 27192 26096 27244 26102
rect 27192 26038 27244 26044
rect 26732 25756 26784 25762
rect 26732 25698 26784 25704
rect 27100 25756 27152 25762
rect 27100 25698 27152 25704
rect 26744 25150 26772 25698
rect 27112 25354 27140 25698
rect 27100 25348 27152 25354
rect 27100 25290 27152 25296
rect 26732 25144 26784 25150
rect 26732 25086 26784 25092
rect 26548 25008 26600 25014
rect 26548 24950 26600 24956
rect 26364 21880 26416 21886
rect 26364 21822 26416 21828
rect 26456 21880 26508 21886
rect 26456 21822 26508 21828
rect 26560 20322 26588 24950
rect 26744 21342 26772 25086
rect 26916 23580 26968 23586
rect 26916 23522 26968 23528
rect 26928 23178 26956 23522
rect 27204 23450 27232 26038
rect 27296 23586 27324 27126
rect 27572 25830 27600 27466
rect 27560 25824 27612 25830
rect 27560 25766 27612 25772
rect 27572 25354 27600 25766
rect 27848 25762 27876 28010
rect 28032 26306 28060 28350
rect 28124 27938 28152 28418
rect 28492 28278 28520 29302
rect 28480 28272 28532 28278
rect 28480 28214 28532 28220
rect 28112 27932 28164 27938
rect 28112 27874 28164 27880
rect 28124 27462 28152 27874
rect 28112 27456 28164 27462
rect 28112 27398 28164 27404
rect 28296 27184 28348 27190
rect 28296 27126 28348 27132
rect 28020 26300 28072 26306
rect 28020 26242 28072 26248
rect 27836 25756 27888 25762
rect 27836 25698 27888 25704
rect 27560 25348 27612 25354
rect 27560 25290 27612 25296
rect 27848 25014 27876 25698
rect 27836 25008 27888 25014
rect 27836 24950 27888 24956
rect 27376 24668 27428 24674
rect 27376 24610 27428 24616
rect 27560 24668 27612 24674
rect 27560 24610 27612 24616
rect 27388 24266 27416 24610
rect 27376 24260 27428 24266
rect 27376 24202 27428 24208
rect 27376 24056 27428 24062
rect 27376 23998 27428 24004
rect 27284 23580 27336 23586
rect 27284 23522 27336 23528
rect 27008 23444 27060 23450
rect 27008 23386 27060 23392
rect 27192 23444 27244 23450
rect 27192 23386 27244 23392
rect 26916 23172 26968 23178
rect 26916 23114 26968 23120
rect 27020 22838 27048 23386
rect 27204 23178 27232 23386
rect 27192 23172 27244 23178
rect 27192 23114 27244 23120
rect 27192 22968 27244 22974
rect 27192 22910 27244 22916
rect 27284 22968 27336 22974
rect 27284 22910 27336 22916
rect 27008 22832 27060 22838
rect 27008 22774 27060 22780
rect 27020 22548 27048 22774
rect 27100 22560 27152 22566
rect 27020 22520 27100 22548
rect 26916 22492 26968 22498
rect 26916 22434 26968 22440
rect 26928 21954 26956 22434
rect 26916 21948 26968 21954
rect 26916 21890 26968 21896
rect 27020 21410 27048 22520
rect 27100 22502 27152 22508
rect 27100 21744 27152 21750
rect 27100 21686 27152 21692
rect 27112 21449 27140 21686
rect 27098 21440 27154 21449
rect 27008 21404 27060 21410
rect 27098 21375 27154 21384
rect 27008 21346 27060 21352
rect 26732 21336 26784 21342
rect 26732 21278 26784 21284
rect 26744 21002 26772 21278
rect 26732 20996 26784 21002
rect 26732 20938 26784 20944
rect 27020 20866 27048 21346
rect 27008 20860 27060 20866
rect 27008 20802 27060 20808
rect 27204 20458 27232 22910
rect 27192 20452 27244 20458
rect 27192 20394 27244 20400
rect 26548 20316 26600 20322
rect 26548 20258 26600 20264
rect 27204 19914 27232 20394
rect 27192 19908 27244 19914
rect 27192 19850 27244 19856
rect 26732 19636 26784 19642
rect 26732 19578 26784 19584
rect 26456 19568 26508 19574
rect 26456 19510 26508 19516
rect 26468 18146 26496 19510
rect 26744 19166 26772 19578
rect 26916 19228 26968 19234
rect 26916 19170 26968 19176
rect 26732 19160 26784 19166
rect 26732 19102 26784 19108
rect 26744 18826 26772 19102
rect 26928 18826 26956 19170
rect 26732 18820 26784 18826
rect 26732 18762 26784 18768
rect 26916 18820 26968 18826
rect 26916 18762 26968 18768
rect 26640 18548 26692 18554
rect 26640 18490 26692 18496
rect 26652 18214 26680 18490
rect 26640 18208 26692 18214
rect 26640 18150 26692 18156
rect 26456 18140 26508 18146
rect 26456 18082 26508 18088
rect 26468 17670 26496 18082
rect 26456 17664 26508 17670
rect 26456 17606 26508 17612
rect 26652 17602 26680 18150
rect 26916 17936 26968 17942
rect 26916 17878 26968 17884
rect 26928 17738 26956 17878
rect 26916 17732 26968 17738
rect 26968 17692 27140 17720
rect 26916 17674 26968 17680
rect 26640 17596 26692 17602
rect 26640 17538 26692 17544
rect 26914 17360 26970 17369
rect 26914 17295 26970 17304
rect 26928 16650 26956 17295
rect 26916 16644 26968 16650
rect 26916 16586 26968 16592
rect 26732 16100 26784 16106
rect 26732 16042 26784 16048
rect 26548 15760 26600 15766
rect 26548 15702 26600 15708
rect 26560 15426 26588 15702
rect 26744 15562 26772 16042
rect 27112 15816 27140 17692
rect 27192 17392 27244 17398
rect 27192 17334 27244 17340
rect 27204 17194 27232 17334
rect 27192 17188 27244 17194
rect 27192 17130 27244 17136
rect 27296 16106 27324 22910
rect 27388 21392 27416 23998
rect 27572 23994 27600 24610
rect 27560 23988 27612 23994
rect 27560 23930 27612 23936
rect 27560 23580 27612 23586
rect 27560 23522 27612 23528
rect 27468 23512 27520 23518
rect 27468 23454 27520 23460
rect 27480 23110 27508 23454
rect 27468 23104 27520 23110
rect 27468 23046 27520 23052
rect 27572 23042 27600 23522
rect 27560 23036 27612 23042
rect 27560 22978 27612 22984
rect 27572 21546 27600 22978
rect 27848 22786 27876 24950
rect 28204 24668 28256 24674
rect 28204 24610 28256 24616
rect 28216 24266 28244 24610
rect 27928 24260 27980 24266
rect 27928 24202 27980 24208
rect 28204 24260 28256 24266
rect 28204 24202 28256 24208
rect 27940 22906 27968 24202
rect 27928 22900 27980 22906
rect 27928 22842 27980 22848
rect 27848 22758 27968 22786
rect 27560 21540 27612 21546
rect 27560 21482 27612 21488
rect 27468 21404 27520 21410
rect 27388 21364 27468 21392
rect 27468 21346 27520 21352
rect 27744 21404 27796 21410
rect 27744 21346 27796 21352
rect 27480 21002 27508 21346
rect 27652 21336 27704 21342
rect 27652 21278 27704 21284
rect 27664 21002 27692 21278
rect 27468 20996 27520 21002
rect 27468 20938 27520 20944
rect 27652 20996 27704 21002
rect 27652 20938 27704 20944
rect 27560 20928 27612 20934
rect 27560 20870 27612 20876
rect 27376 20316 27428 20322
rect 27376 20258 27428 20264
rect 27388 19846 27416 20258
rect 27468 20248 27520 20254
rect 27468 20190 27520 20196
rect 27376 19840 27428 19846
rect 27376 19782 27428 19788
rect 27376 19568 27428 19574
rect 27480 19556 27508 20190
rect 27428 19528 27508 19556
rect 27376 19510 27428 19516
rect 27284 16100 27336 16106
rect 27284 16042 27336 16048
rect 27112 15788 27232 15816
rect 27204 15562 27232 15788
rect 26732 15556 26784 15562
rect 26732 15498 26784 15504
rect 27192 15556 27244 15562
rect 27192 15498 27244 15504
rect 26916 15488 26968 15494
rect 26916 15430 26968 15436
rect 26548 15420 26600 15426
rect 26548 15362 26600 15368
rect 26272 14876 26324 14882
rect 26272 14818 26324 14824
rect 26456 14876 26508 14882
rect 26456 14818 26508 14824
rect 26180 14808 26232 14814
rect 26180 14750 26232 14756
rect 26272 14740 26324 14746
rect 26272 14682 26324 14688
rect 26088 14468 26140 14474
rect 26088 14410 26140 14416
rect 26284 14134 26312 14682
rect 26468 14214 26496 14818
rect 26928 14474 26956 15430
rect 27204 15358 27232 15498
rect 27100 15352 27152 15358
rect 27100 15294 27152 15300
rect 27192 15352 27244 15358
rect 27192 15294 27244 15300
rect 27112 15018 27140 15294
rect 27100 15012 27152 15018
rect 27100 14954 27152 14960
rect 27204 14882 27232 15294
rect 27008 14876 27060 14882
rect 27008 14818 27060 14824
rect 27192 14876 27244 14882
rect 27192 14818 27244 14824
rect 26916 14468 26968 14474
rect 26916 14410 26968 14416
rect 26824 14400 26876 14406
rect 26824 14342 26876 14348
rect 26836 14270 26864 14342
rect 26376 14186 26496 14214
rect 26824 14264 26876 14270
rect 26824 14206 26876 14212
rect 25996 14128 26048 14134
rect 25916 14088 25996 14116
rect 25916 13794 25944 14088
rect 25996 14070 26048 14076
rect 26272 14128 26324 14134
rect 26272 14070 26324 14076
rect 25812 13788 25864 13794
rect 25812 13730 25864 13736
rect 25904 13788 25956 13794
rect 25904 13730 25956 13736
rect 25536 13584 25588 13590
rect 25536 13526 25588 13532
rect 25548 13182 25576 13526
rect 25824 13386 25852 13730
rect 25812 13380 25864 13386
rect 25812 13322 25864 13328
rect 25536 13176 25588 13182
rect 25536 13118 25588 13124
rect 25812 13176 25864 13182
rect 25812 13118 25864 13124
rect 25352 11136 25404 11142
rect 25352 11078 25404 11084
rect 24892 11000 24944 11006
rect 24812 10960 24892 10988
rect 24616 10116 24668 10122
rect 24616 10058 24668 10064
rect 24628 9918 24656 10058
rect 24616 9912 24668 9918
rect 24616 9854 24668 9860
rect 24628 9578 24656 9854
rect 24616 9572 24668 9578
rect 24616 9514 24668 9520
rect 24708 9572 24760 9578
rect 24708 9514 24760 9520
rect 24628 9374 24656 9514
rect 24616 9368 24668 9374
rect 24616 9310 24668 9316
rect 24720 9034 24748 9514
rect 24708 9028 24760 9034
rect 24708 8970 24760 8976
rect 24616 8960 24668 8966
rect 24616 8902 24668 8908
rect 24628 8422 24656 8902
rect 24616 8416 24668 8422
rect 24668 8376 24748 8404
rect 24616 8358 24668 8364
rect 24524 8348 24576 8354
rect 24524 8290 24576 8296
rect 24536 7402 24564 8290
rect 24616 7668 24668 7674
rect 24616 7610 24668 7616
rect 24524 7396 24576 7402
rect 24524 7338 24576 7344
rect 24628 6858 24656 7610
rect 24720 7402 24748 8376
rect 24812 7878 24840 10960
rect 24892 10942 24944 10948
rect 25352 10048 25404 10054
rect 25352 9990 25404 9996
rect 25364 9782 25392 9990
rect 25352 9776 25404 9782
rect 25352 9718 25404 9724
rect 25364 8830 25392 9718
rect 25548 9578 25576 13118
rect 25628 10388 25680 10394
rect 25628 10330 25680 10336
rect 25536 9572 25588 9578
rect 25536 9514 25588 9520
rect 25536 9028 25588 9034
rect 25536 8970 25588 8976
rect 25352 8824 25404 8830
rect 25352 8766 25404 8772
rect 25168 8756 25220 8762
rect 25168 8698 25220 8704
rect 25076 8144 25128 8150
rect 25076 8086 25128 8092
rect 24800 7872 24852 7878
rect 24800 7814 24852 7820
rect 24892 7804 24944 7810
rect 24892 7746 24944 7752
rect 24904 7402 24932 7746
rect 25088 7674 25116 8086
rect 25076 7668 25128 7674
rect 25076 7610 25128 7616
rect 24708 7396 24760 7402
rect 24708 7338 24760 7344
rect 24892 7396 24944 7402
rect 24892 7338 24944 7344
rect 24904 6858 24932 7338
rect 24616 6852 24668 6858
rect 24616 6794 24668 6800
rect 24892 6852 24944 6858
rect 24892 6794 24944 6800
rect 24892 5560 24944 5566
rect 24892 5502 24944 5508
rect 24800 5424 24852 5430
rect 24800 5366 24852 5372
rect 24432 5152 24484 5158
rect 24432 5094 24484 5100
rect 24248 5084 24300 5090
rect 24248 5026 24300 5032
rect 24260 4682 24288 5026
rect 24432 5016 24484 5022
rect 24432 4958 24484 4964
rect 24248 4676 24300 4682
rect 24248 4618 24300 4624
rect 24444 4342 24472 4958
rect 24064 4336 24116 4342
rect 24064 4278 24116 4284
rect 24432 4336 24484 4342
rect 24432 4278 24484 4284
rect 24076 4002 24104 4278
rect 24812 4138 24840 5366
rect 24800 4132 24852 4138
rect 24800 4074 24852 4080
rect 23880 3996 23932 4002
rect 23880 3938 23932 3944
rect 24064 3996 24116 4002
rect 24064 3938 24116 3944
rect 23788 3928 23840 3934
rect 23788 3870 23840 3876
rect 23800 3458 23828 3870
rect 23788 3452 23840 3458
rect 23788 3394 23840 3400
rect 23800 3361 23828 3394
rect 23786 3352 23842 3361
rect 23786 3287 23842 3296
rect 23892 3254 23920 3938
rect 24076 3390 24104 3938
rect 24904 3526 24932 5502
rect 25180 4138 25208 8698
rect 25364 8354 25392 8766
rect 25352 8348 25404 8354
rect 25352 8290 25404 8296
rect 25548 7946 25576 8970
rect 25640 8966 25668 10330
rect 25718 10152 25774 10161
rect 25718 10087 25774 10096
rect 25732 9918 25760 10087
rect 25720 9912 25772 9918
rect 25720 9854 25772 9860
rect 25720 9300 25772 9306
rect 25720 9242 25772 9248
rect 25628 8960 25680 8966
rect 25628 8902 25680 8908
rect 25640 8830 25668 8902
rect 25628 8824 25680 8830
rect 25628 8766 25680 8772
rect 25732 8694 25760 9242
rect 25720 8688 25772 8694
rect 25720 8630 25772 8636
rect 25536 7940 25588 7946
rect 25536 7882 25588 7888
rect 25548 7742 25576 7882
rect 25536 7736 25588 7742
rect 25536 7678 25588 7684
rect 25548 6790 25576 7678
rect 25536 6784 25588 6790
rect 25536 6726 25588 6732
rect 25444 6648 25496 6654
rect 25444 6590 25496 6596
rect 25456 5770 25484 6590
rect 25444 5764 25496 5770
rect 25444 5706 25496 5712
rect 25824 5226 25852 13118
rect 25916 13114 25944 13730
rect 26284 13697 26312 14070
rect 26376 13930 26404 14186
rect 26364 13924 26416 13930
rect 26364 13866 26416 13872
rect 26270 13688 26326 13697
rect 26270 13623 26326 13632
rect 26180 13584 26232 13590
rect 26180 13526 26232 13532
rect 26192 13386 26220 13526
rect 26180 13380 26232 13386
rect 26180 13322 26232 13328
rect 26548 13312 26600 13318
rect 26548 13254 26600 13260
rect 25904 13108 25956 13114
rect 25904 13050 25956 13056
rect 26364 12632 26416 12638
rect 26364 12574 26416 12580
rect 26376 11550 26404 12574
rect 26364 11544 26416 11550
rect 26364 11486 26416 11492
rect 26088 10524 26140 10530
rect 26088 10466 26140 10472
rect 25904 10320 25956 10326
rect 25904 10262 25956 10268
rect 25916 9578 25944 10262
rect 26100 10122 26128 10466
rect 26376 10462 26404 11486
rect 26364 10456 26416 10462
rect 26364 10398 26416 10404
rect 26088 10116 26140 10122
rect 26088 10058 26140 10064
rect 26180 10048 26232 10054
rect 26180 9990 26232 9996
rect 26192 9918 26220 9990
rect 26180 9912 26232 9918
rect 26180 9854 26232 9860
rect 25904 9572 25956 9578
rect 25904 9514 25956 9520
rect 25916 8898 25944 9514
rect 26364 9504 26416 9510
rect 26364 9446 26416 9452
rect 25996 9368 26048 9374
rect 25996 9310 26048 9316
rect 25904 8892 25956 8898
rect 25904 8834 25956 8840
rect 25904 8688 25956 8694
rect 26008 8676 26036 9310
rect 25956 8648 26036 8676
rect 25904 8630 25956 8636
rect 25916 8286 25944 8630
rect 26376 8490 26404 9446
rect 26456 8756 26508 8762
rect 26456 8698 26508 8704
rect 26364 8484 26416 8490
rect 26364 8426 26416 8432
rect 26468 8422 26496 8698
rect 26456 8416 26508 8422
rect 26456 8358 26508 8364
rect 25904 8280 25956 8286
rect 25902 8248 25904 8257
rect 25956 8248 25958 8257
rect 25902 8183 25958 8192
rect 25916 8157 25944 8183
rect 26560 7198 26588 13254
rect 26732 13040 26784 13046
rect 26732 12982 26784 12988
rect 26744 12026 26772 12982
rect 26836 12162 26864 14206
rect 26928 13930 26956 14410
rect 27020 14202 27048 14818
rect 27008 14196 27060 14202
rect 27008 14138 27060 14144
rect 26916 13924 26968 13930
rect 26916 13866 26968 13872
rect 27020 12842 27048 14138
rect 27388 13182 27416 19510
rect 27572 16038 27600 20870
rect 27756 20798 27784 21346
rect 27744 20792 27796 20798
rect 27744 20734 27796 20740
rect 27652 20724 27704 20730
rect 27652 20666 27704 20672
rect 27664 19166 27692 20666
rect 27836 20316 27888 20322
rect 27836 20258 27888 20264
rect 27848 19642 27876 20258
rect 27940 19710 27968 22758
rect 28308 21206 28336 27126
rect 28492 25098 28520 28214
rect 28572 26844 28624 26850
rect 28572 26786 28624 26792
rect 28584 26442 28612 26786
rect 28754 26744 28810 26753
rect 28754 26679 28810 26688
rect 28768 26646 28796 26679
rect 28756 26640 28808 26646
rect 28756 26582 28808 26588
rect 28768 26442 28796 26582
rect 28572 26436 28624 26442
rect 28572 26378 28624 26384
rect 28756 26436 28808 26442
rect 28756 26378 28808 26384
rect 28572 25688 28624 25694
rect 28572 25630 28624 25636
rect 28584 25218 28612 25630
rect 28572 25212 28624 25218
rect 28572 25154 28624 25160
rect 28388 25076 28440 25082
rect 28492 25070 28612 25098
rect 28388 25018 28440 25024
rect 28400 24538 28428 25018
rect 28480 25008 28532 25014
rect 28480 24950 28532 24956
rect 28388 24532 28440 24538
rect 28388 24474 28440 24480
rect 28400 24198 28428 24474
rect 28388 24192 28440 24198
rect 28388 24134 28440 24140
rect 28492 24062 28520 24950
rect 28480 24056 28532 24062
rect 28480 23998 28532 24004
rect 28480 23580 28532 23586
rect 28480 23522 28532 23528
rect 28492 23110 28520 23522
rect 28480 23104 28532 23110
rect 28480 23046 28532 23052
rect 28584 22498 28612 25070
rect 28572 22492 28624 22498
rect 28572 22434 28624 22440
rect 28756 22492 28808 22498
rect 28756 22434 28808 22440
rect 28584 22090 28612 22434
rect 28768 22090 28796 22434
rect 28848 22288 28900 22294
rect 28848 22230 28900 22236
rect 28860 22090 28888 22230
rect 28572 22084 28624 22090
rect 28572 22026 28624 22032
rect 28756 22084 28808 22090
rect 28756 22026 28808 22032
rect 28848 22084 28900 22090
rect 28848 22026 28900 22032
rect 28664 22016 28716 22022
rect 28664 21958 28716 21964
rect 28572 21404 28624 21410
rect 28492 21364 28572 21392
rect 28296 21200 28348 21206
rect 28296 21142 28348 21148
rect 28492 20934 28520 21364
rect 28572 21346 28624 21352
rect 28572 21200 28624 21206
rect 28572 21142 28624 21148
rect 28480 20928 28532 20934
rect 28480 20870 28532 20876
rect 28584 20866 28612 21142
rect 28572 20860 28624 20866
rect 28572 20802 28624 20808
rect 28112 20656 28164 20662
rect 28112 20598 28164 20604
rect 28296 20656 28348 20662
rect 28296 20598 28348 20604
rect 28020 20384 28072 20390
rect 28020 20326 28072 20332
rect 28032 19846 28060 20326
rect 28124 20236 28152 20598
rect 28204 20248 28256 20254
rect 28124 20208 28204 20236
rect 28124 19914 28152 20208
rect 28204 20190 28256 20196
rect 28308 20186 28336 20598
rect 28388 20452 28440 20458
rect 28388 20394 28440 20400
rect 28400 20322 28428 20394
rect 28388 20316 28440 20322
rect 28388 20258 28440 20264
rect 28296 20180 28348 20186
rect 28296 20122 28348 20128
rect 28112 19908 28164 19914
rect 28112 19850 28164 19856
rect 28020 19840 28072 19846
rect 28020 19782 28072 19788
rect 27928 19704 27980 19710
rect 27980 19664 28060 19692
rect 27928 19646 27980 19652
rect 27836 19636 27888 19642
rect 27836 19578 27888 19584
rect 27928 19228 27980 19234
rect 27928 19170 27980 19176
rect 27652 19160 27704 19166
rect 27652 19102 27704 19108
rect 27664 18758 27692 19102
rect 27652 18752 27704 18758
rect 27652 18694 27704 18700
rect 27744 18616 27796 18622
rect 27744 18558 27796 18564
rect 27756 17058 27784 18558
rect 27836 17120 27888 17126
rect 27836 17062 27888 17068
rect 27744 17052 27796 17058
rect 27744 16994 27796 17000
rect 27756 16582 27784 16994
rect 27848 16650 27876 17062
rect 27940 16854 27968 19170
rect 28032 18146 28060 19664
rect 28204 19296 28256 19302
rect 28204 19238 28256 19244
rect 28112 19160 28164 19166
rect 28112 19102 28164 19108
rect 28124 18826 28152 19102
rect 28112 18820 28164 18826
rect 28112 18762 28164 18768
rect 28216 18758 28244 19238
rect 28204 18752 28256 18758
rect 28204 18694 28256 18700
rect 28216 18622 28244 18694
rect 28204 18616 28256 18622
rect 28204 18558 28256 18564
rect 28112 18480 28164 18486
rect 28112 18422 28164 18428
rect 28020 18140 28072 18146
rect 28020 18082 28072 18088
rect 28032 17670 28060 18082
rect 28020 17664 28072 17670
rect 28020 17606 28072 17612
rect 28020 17052 28072 17058
rect 28020 16994 28072 17000
rect 27928 16848 27980 16854
rect 27928 16790 27980 16796
rect 27940 16650 27968 16790
rect 27836 16644 27888 16650
rect 27836 16586 27888 16592
rect 27928 16644 27980 16650
rect 27928 16586 27980 16592
rect 27744 16576 27796 16582
rect 27744 16518 27796 16524
rect 28032 16310 28060 16994
rect 28020 16304 28072 16310
rect 28020 16246 28072 16252
rect 27560 16032 27612 16038
rect 27612 15992 27784 16020
rect 27560 15974 27612 15980
rect 27560 15420 27612 15426
rect 27560 15362 27612 15368
rect 27376 13176 27428 13182
rect 27376 13118 27428 13124
rect 27008 12836 27060 12842
rect 27008 12778 27060 12784
rect 27020 12298 27048 12778
rect 27376 12700 27428 12706
rect 27376 12642 27428 12648
rect 27008 12292 27060 12298
rect 27008 12234 27060 12240
rect 26824 12156 26876 12162
rect 26824 12098 26876 12104
rect 27284 12088 27336 12094
rect 27284 12030 27336 12036
rect 26732 12020 26784 12026
rect 26732 11962 26784 11968
rect 27192 12020 27244 12026
rect 27192 11962 27244 11968
rect 27204 11686 27232 11962
rect 27192 11680 27244 11686
rect 27192 11622 27244 11628
rect 26732 11544 26784 11550
rect 26732 11486 26784 11492
rect 26744 11210 26772 11486
rect 26732 11204 26784 11210
rect 26732 11146 26784 11152
rect 26640 11000 26692 11006
rect 26640 10942 26692 10948
rect 26652 10598 26680 10942
rect 26744 10666 26772 11146
rect 27008 11068 27060 11074
rect 27008 11010 27060 11016
rect 26916 10864 26968 10870
rect 26916 10806 26968 10812
rect 26732 10660 26784 10666
rect 26732 10602 26784 10608
rect 26640 10592 26692 10598
rect 26640 10534 26692 10540
rect 26640 9436 26692 9442
rect 26640 9378 26692 9384
rect 26652 8898 26680 9378
rect 26640 8892 26692 8898
rect 26640 8834 26692 8840
rect 26652 8218 26680 8834
rect 26640 8212 26692 8218
rect 26640 8154 26692 8160
rect 26652 7334 26680 8154
rect 26640 7328 26692 7334
rect 26640 7270 26692 7276
rect 26548 7192 26600 7198
rect 26548 7134 26600 7140
rect 26560 6654 26588 7134
rect 26652 6790 26680 7270
rect 26928 7062 26956 10806
rect 27020 9442 27048 11010
rect 27100 11000 27152 11006
rect 27100 10942 27152 10948
rect 27112 10666 27140 10942
rect 27204 10938 27232 11622
rect 27192 10932 27244 10938
rect 27192 10874 27244 10880
rect 27100 10660 27152 10666
rect 27100 10602 27152 10608
rect 27296 9782 27324 12030
rect 27388 11958 27416 12642
rect 27376 11952 27428 11958
rect 27376 11894 27428 11900
rect 27100 9776 27152 9782
rect 27100 9718 27152 9724
rect 27284 9776 27336 9782
rect 27284 9718 27336 9724
rect 27008 9436 27060 9442
rect 27008 9378 27060 9384
rect 27020 8966 27048 9378
rect 27008 8960 27060 8966
rect 27008 8902 27060 8908
rect 27112 8830 27140 9718
rect 27192 9368 27244 9374
rect 27192 9310 27244 9316
rect 27204 9034 27232 9310
rect 27192 9028 27244 9034
rect 27192 8970 27244 8976
rect 27296 8830 27324 9718
rect 27100 8824 27152 8830
rect 27100 8766 27152 8772
rect 27284 8824 27336 8830
rect 27284 8766 27336 8772
rect 27112 8490 27140 8766
rect 27100 8484 27152 8490
rect 27100 8426 27152 8432
rect 27296 8150 27324 8766
rect 27388 8422 27416 11894
rect 27468 11476 27520 11482
rect 27468 11418 27520 11424
rect 27480 11006 27508 11418
rect 27468 11000 27520 11006
rect 27468 10942 27520 10948
rect 27480 10870 27508 10942
rect 27468 10864 27520 10870
rect 27468 10806 27520 10812
rect 27572 9510 27600 15362
rect 27652 15284 27704 15290
rect 27652 15226 27704 15232
rect 27664 9510 27692 15226
rect 27756 14950 27784 15992
rect 27836 15420 27888 15426
rect 27836 15362 27888 15368
rect 27848 15329 27876 15362
rect 27834 15320 27890 15329
rect 27834 15255 27890 15264
rect 27744 14944 27796 14950
rect 27744 14886 27796 14892
rect 28032 10666 28060 16246
rect 28124 15902 28152 18422
rect 28400 18214 28428 20258
rect 28584 19778 28612 20802
rect 28572 19772 28624 19778
rect 28572 19714 28624 19720
rect 28676 19302 28704 21958
rect 28860 20390 28888 22026
rect 28848 20384 28900 20390
rect 28848 20326 28900 20332
rect 28664 19296 28716 19302
rect 28664 19238 28716 19244
rect 28388 18208 28440 18214
rect 28388 18150 28440 18156
rect 28756 18208 28808 18214
rect 28756 18150 28808 18156
rect 28400 17602 28428 18150
rect 28388 17596 28440 17602
rect 28388 17538 28440 17544
rect 28480 17460 28532 17466
rect 28480 17402 28532 17408
rect 28492 15970 28520 17402
rect 28572 17392 28624 17398
rect 28768 17380 28796 18150
rect 28624 17352 28796 17380
rect 28572 17334 28624 17340
rect 28204 15964 28256 15970
rect 28204 15906 28256 15912
rect 28480 15964 28532 15970
rect 28480 15906 28532 15912
rect 28112 15896 28164 15902
rect 28112 15838 28164 15844
rect 28124 15562 28152 15838
rect 28112 15556 28164 15562
rect 28112 15498 28164 15504
rect 28216 15494 28244 15906
rect 28388 15896 28440 15902
rect 28388 15838 28440 15844
rect 28204 15488 28256 15494
rect 28204 15430 28256 15436
rect 28400 15290 28428 15838
rect 28492 15358 28520 15906
rect 28480 15352 28532 15358
rect 28480 15294 28532 15300
rect 28388 15284 28440 15290
rect 28388 15226 28440 15232
rect 28584 14241 28612 17334
rect 28848 15556 28900 15562
rect 28848 15498 28900 15504
rect 28664 15352 28716 15358
rect 28664 15294 28716 15300
rect 28676 14474 28704 15294
rect 28860 15018 28888 15498
rect 28848 15012 28900 15018
rect 28848 14954 28900 14960
rect 28664 14468 28716 14474
rect 28664 14410 28716 14416
rect 28570 14232 28626 14241
rect 28952 14214 28980 29366
rect 29412 29162 29440 29370
rect 29400 29156 29452 29162
rect 29400 29098 29452 29104
rect 29032 28272 29084 28278
rect 29032 28214 29084 28220
rect 29044 18758 29072 28214
rect 29308 26164 29360 26170
rect 29308 26106 29360 26112
rect 29320 25082 29348 26106
rect 29308 25076 29360 25082
rect 29308 25018 29360 25024
rect 29320 24810 29348 25018
rect 29308 24804 29360 24810
rect 29308 24746 29360 24752
rect 29216 24600 29268 24606
rect 29216 24542 29268 24548
rect 29228 24062 29256 24542
rect 29308 24260 29360 24266
rect 29308 24202 29360 24208
rect 29216 24056 29268 24062
rect 29216 23998 29268 24004
rect 29320 21002 29348 24202
rect 29308 20996 29360 21002
rect 29308 20938 29360 20944
rect 29320 20730 29348 20938
rect 29308 20724 29360 20730
rect 29308 20666 29360 20672
rect 29504 20254 29532 31662
rect 29860 30108 29912 30114
rect 29860 30050 29912 30056
rect 29768 29020 29820 29026
rect 29768 28962 29820 28968
rect 29584 28408 29636 28414
rect 29584 28350 29636 28356
rect 29596 28074 29624 28350
rect 29780 28278 29808 28962
rect 29872 28822 29900 30050
rect 29950 29600 30006 29609
rect 29950 29535 30006 29544
rect 29964 29162 29992 29535
rect 29952 29156 30004 29162
rect 29952 29098 30004 29104
rect 29860 28816 29912 28822
rect 29860 28758 29912 28764
rect 29768 28272 29820 28278
rect 29768 28214 29820 28220
rect 29584 28068 29636 28074
rect 29584 28010 29636 28016
rect 29676 27932 29728 27938
rect 29676 27874 29728 27880
rect 29688 27190 29716 27874
rect 29676 27184 29728 27190
rect 29676 27126 29728 27132
rect 29872 26238 29900 28758
rect 29964 28618 29992 29098
rect 29952 28612 30004 28618
rect 29952 28554 30004 28560
rect 30044 27864 30096 27870
rect 30044 27806 30096 27812
rect 30056 27705 30084 27806
rect 30042 27696 30098 27705
rect 30042 27631 30098 27640
rect 30056 27530 30084 27631
rect 30044 27524 30096 27530
rect 30044 27466 30096 27472
rect 30044 26368 30096 26374
rect 30044 26310 30096 26316
rect 29860 26232 29912 26238
rect 29860 26174 29912 26180
rect 29872 26102 29900 26174
rect 29860 26096 29912 26102
rect 29860 26038 29912 26044
rect 29872 24674 29900 26038
rect 30056 25529 30084 26310
rect 30042 25520 30098 25529
rect 30042 25455 30098 25464
rect 29860 24668 29912 24674
rect 29860 24610 29912 24616
rect 29768 24600 29820 24606
rect 29768 24542 29820 24548
rect 29780 24266 29808 24542
rect 29872 24266 29900 24610
rect 29768 24260 29820 24266
rect 29768 24202 29820 24208
rect 29860 24260 29912 24266
rect 29860 24202 29912 24208
rect 29768 24124 29820 24130
rect 29768 24066 29820 24072
rect 29584 21336 29636 21342
rect 29584 21278 29636 21284
rect 29492 20248 29544 20254
rect 29492 20190 29544 20196
rect 29400 19296 29452 19302
rect 29400 19238 29452 19244
rect 29124 19228 29176 19234
rect 29124 19170 29176 19176
rect 29136 18826 29164 19170
rect 29124 18820 29176 18826
rect 29124 18762 29176 18768
rect 29032 18752 29084 18758
rect 29032 18694 29084 18700
rect 29412 18690 29440 19238
rect 29596 19166 29624 21278
rect 29584 19160 29636 19166
rect 29584 19102 29636 19108
rect 29596 18826 29624 19102
rect 29492 18820 29544 18826
rect 29492 18762 29544 18768
rect 29584 18820 29636 18826
rect 29584 18762 29636 18768
rect 29400 18684 29452 18690
rect 29400 18626 29452 18632
rect 29504 18570 29532 18762
rect 29412 18542 29532 18570
rect 29412 18486 29440 18542
rect 29400 18480 29452 18486
rect 29400 18422 29452 18428
rect 28952 14186 29072 14214
rect 28570 14167 28626 14176
rect 28848 14128 28900 14134
rect 28848 14070 28900 14076
rect 28388 13720 28440 13726
rect 28388 13662 28440 13668
rect 28756 13720 28808 13726
rect 28756 13662 28808 13668
rect 28400 13114 28428 13662
rect 28768 13386 28796 13662
rect 28756 13380 28808 13386
rect 28756 13322 28808 13328
rect 28388 13108 28440 13114
rect 28388 13050 28440 13056
rect 28400 12638 28428 13050
rect 28572 13040 28624 13046
rect 28572 12982 28624 12988
rect 28584 12824 28612 12982
rect 28664 12836 28716 12842
rect 28584 12796 28664 12824
rect 28388 12632 28440 12638
rect 28388 12574 28440 12580
rect 28400 12230 28428 12574
rect 28388 12224 28440 12230
rect 28388 12166 28440 12172
rect 28584 12026 28612 12796
rect 28664 12778 28716 12784
rect 28756 12632 28808 12638
rect 28756 12574 28808 12580
rect 28768 12298 28796 12574
rect 28756 12292 28808 12298
rect 28756 12234 28808 12240
rect 28572 12020 28624 12026
rect 28572 11962 28624 11968
rect 28768 11754 28796 12234
rect 28756 11748 28808 11754
rect 28756 11690 28808 11696
rect 28112 11544 28164 11550
rect 28112 11486 28164 11492
rect 28204 11544 28256 11550
rect 28860 11521 28888 14070
rect 29044 13726 29072 14186
rect 29412 14134 29440 18422
rect 29400 14128 29452 14134
rect 29400 14070 29452 14076
rect 29124 13856 29176 13862
rect 29124 13798 29176 13804
rect 29032 13720 29084 13726
rect 29032 13662 29084 13668
rect 29044 13046 29072 13662
rect 29032 13040 29084 13046
rect 29032 12982 29084 12988
rect 28940 12156 28992 12162
rect 28940 12098 28992 12104
rect 28204 11486 28256 11492
rect 28846 11512 28902 11521
rect 28124 11074 28152 11486
rect 28112 11068 28164 11074
rect 28112 11010 28164 11016
rect 28020 10660 28072 10666
rect 28020 10602 28072 10608
rect 28216 10598 28244 11486
rect 28846 11447 28902 11456
rect 28664 11408 28716 11414
rect 28716 11368 28796 11396
rect 28664 11350 28716 11356
rect 28768 11006 28796 11368
rect 28756 11000 28808 11006
rect 28756 10942 28808 10948
rect 28664 10660 28716 10666
rect 28664 10602 28716 10608
rect 28204 10592 28256 10598
rect 28204 10534 28256 10540
rect 27560 9504 27612 9510
rect 27560 9446 27612 9452
rect 27652 9504 27704 9510
rect 27652 9446 27704 9452
rect 27468 9436 27520 9442
rect 27468 9378 27520 9384
rect 27480 9034 27508 9378
rect 27468 9028 27520 9034
rect 27468 8970 27520 8976
rect 27468 8824 27520 8830
rect 27468 8766 27520 8772
rect 27652 8824 27704 8830
rect 27652 8766 27704 8772
rect 27376 8416 27428 8422
rect 27376 8358 27428 8364
rect 27480 8354 27508 8766
rect 27468 8348 27520 8354
rect 27468 8290 27520 8296
rect 27284 8144 27336 8150
rect 27284 8086 27336 8092
rect 27480 7946 27508 8290
rect 27664 8218 27692 8766
rect 27652 8212 27704 8218
rect 27652 8154 27704 8160
rect 27468 7940 27520 7946
rect 27468 7882 27520 7888
rect 26916 7056 26968 7062
rect 26916 6998 26968 7004
rect 26928 6790 26956 6998
rect 26640 6784 26692 6790
rect 26640 6726 26692 6732
rect 26916 6784 26968 6790
rect 26916 6726 26968 6732
rect 26548 6648 26600 6654
rect 26548 6590 26600 6596
rect 26652 6178 26680 6726
rect 26640 6172 26692 6178
rect 26640 6114 26692 6120
rect 26652 5770 26680 6114
rect 26640 5764 26692 5770
rect 26640 5706 26692 5712
rect 26180 5696 26232 5702
rect 26180 5638 26232 5644
rect 26546 5664 26602 5673
rect 25260 5220 25312 5226
rect 25260 5162 25312 5168
rect 25812 5220 25864 5226
rect 25812 5162 25864 5168
rect 25168 4132 25220 4138
rect 25168 4074 25220 4080
rect 25180 3526 25208 4074
rect 24892 3520 24944 3526
rect 24892 3462 24944 3468
rect 25168 3520 25220 3526
rect 25168 3462 25220 3468
rect 24064 3384 24116 3390
rect 24064 3326 24116 3332
rect 23880 3248 23932 3254
rect 23880 3190 23932 3196
rect 23696 2840 23748 2846
rect 23696 2782 23748 2788
rect 23604 2704 23656 2710
rect 23604 2646 23656 2652
rect 23328 2364 23380 2370
rect 23328 2306 23380 2312
rect 23420 2296 23472 2302
rect 22500 2228 22552 2234
rect 22500 2170 22552 2176
rect 23144 2228 23196 2234
rect 23248 2222 23368 2250
rect 23420 2238 23472 2244
rect 23144 2170 23196 2176
rect 21212 1888 21264 1894
rect 21212 1830 21264 1836
rect 21764 1888 21816 1894
rect 21764 1830 21816 1836
rect 21224 1282 21252 1830
rect 21776 1418 21804 1830
rect 22040 1752 22092 1758
rect 22040 1694 22092 1700
rect 21764 1412 21816 1418
rect 21764 1354 21816 1360
rect 21212 1276 21264 1282
rect 21212 1218 21264 1224
rect 22052 1214 22080 1694
rect 22040 1208 22092 1214
rect 22040 1150 22092 1156
rect 20934 632 20990 641
rect 20934 567 20990 576
rect 21028 528 21080 534
rect 20566 496 20622 505
rect 20566 431 20622 440
rect 20750 496 20806 505
rect 21028 470 21080 476
rect 20750 431 20806 440
rect 21040 424 21068 470
rect 22512 424 22540 2170
rect 23340 2166 23368 2222
rect 23328 2160 23380 2166
rect 23328 2102 23380 2108
rect 23052 1820 23104 1826
rect 23052 1762 23104 1768
rect 22592 1752 22644 1758
rect 22592 1694 22644 1700
rect 22604 1350 22632 1694
rect 22592 1344 22644 1350
rect 22592 1286 22644 1292
rect 23064 1078 23092 1762
rect 23340 1350 23368 2102
rect 23328 1344 23380 1350
rect 23328 1286 23380 1292
rect 23432 1214 23460 2238
rect 23708 1758 23736 2782
rect 23892 1826 23920 3190
rect 24076 1826 24104 3326
rect 24800 3248 24852 3254
rect 24800 3190 24852 3196
rect 24432 2500 24484 2506
rect 24432 2442 24484 2448
rect 24444 2234 24472 2442
rect 24432 2228 24484 2234
rect 24432 2170 24484 2176
rect 23880 1820 23932 1826
rect 23880 1762 23932 1768
rect 24064 1820 24116 1826
rect 24064 1762 24116 1768
rect 23696 1752 23748 1758
rect 23696 1694 23748 1700
rect 23696 1616 23748 1622
rect 23696 1558 23748 1564
rect 23708 1282 23736 1558
rect 23696 1276 23748 1282
rect 23696 1218 23748 1224
rect 23420 1208 23472 1214
rect 23420 1150 23472 1156
rect 23052 1072 23104 1078
rect 23052 1014 23104 1020
rect 23064 534 23092 1014
rect 23432 806 23460 1150
rect 23708 874 23736 1218
rect 23788 1072 23840 1078
rect 23788 1014 23840 1020
rect 23696 868 23748 874
rect 23696 810 23748 816
rect 23420 800 23472 806
rect 23420 742 23472 748
rect 23052 528 23104 534
rect 23052 470 23104 476
rect 23800 424 23828 1014
rect 23892 874 23920 1762
rect 24076 1418 24104 1762
rect 24444 1418 24472 2170
rect 24812 1826 24840 3190
rect 24800 1820 24852 1826
rect 24800 1762 24852 1768
rect 24064 1412 24116 1418
rect 24064 1354 24116 1360
rect 24432 1412 24484 1418
rect 24432 1354 24484 1360
rect 24444 1146 24472 1354
rect 24812 1350 24840 1762
rect 24800 1344 24852 1350
rect 24800 1286 24852 1292
rect 24432 1140 24484 1146
rect 24432 1082 24484 1088
rect 23880 868 23932 874
rect 23880 810 23932 816
rect 25272 424 25300 5162
rect 26192 4070 26220 5638
rect 26652 5634 26680 5706
rect 26546 5599 26602 5608
rect 26640 5628 26692 5634
rect 26560 5566 26588 5599
rect 26640 5570 26692 5576
rect 26548 5560 26600 5566
rect 26548 5502 26600 5508
rect 26180 4064 26232 4070
rect 26180 4006 26232 4012
rect 26088 3996 26140 4002
rect 26088 3938 26140 3944
rect 25442 3488 25498 3497
rect 25442 3423 25498 3432
rect 25456 2506 25484 3423
rect 26100 3390 26128 3938
rect 25536 3384 25588 3390
rect 26088 3384 26140 3390
rect 25588 3344 25668 3372
rect 25536 3326 25588 3332
rect 25444 2500 25496 2506
rect 25444 2442 25496 2448
rect 25640 2234 25668 3344
rect 26088 3326 26140 3332
rect 26100 2982 26128 3326
rect 26192 3050 26220 4006
rect 26560 3390 26588 5502
rect 26928 5430 26956 6726
rect 27664 6042 27692 8154
rect 28112 7600 28164 7606
rect 28112 7542 28164 7548
rect 28124 7266 28152 7542
rect 28112 7260 28164 7266
rect 28112 7202 28164 7208
rect 27836 7192 27888 7198
rect 27836 7134 27888 7140
rect 27848 6790 27876 7134
rect 28020 7124 28072 7130
rect 28020 7066 28072 7072
rect 27836 6784 27888 6790
rect 27836 6726 27888 6732
rect 28032 6722 28060 7066
rect 28124 6858 28152 7202
rect 28112 6852 28164 6858
rect 28112 6794 28164 6800
rect 28020 6716 28072 6722
rect 28020 6658 28072 6664
rect 28020 6308 28072 6314
rect 28020 6250 28072 6256
rect 27744 6172 27796 6178
rect 27744 6114 27796 6120
rect 27652 6036 27704 6042
rect 27652 5978 27704 5984
rect 27100 5492 27152 5498
rect 27100 5434 27152 5440
rect 26916 5424 26968 5430
rect 26916 5366 26968 5372
rect 27112 5090 27140 5434
rect 27664 5226 27692 5978
rect 27756 5702 27784 6114
rect 27744 5696 27796 5702
rect 27744 5638 27796 5644
rect 27652 5220 27704 5226
rect 27652 5162 27704 5168
rect 28032 5090 28060 6250
rect 28216 6178 28244 10534
rect 28676 10122 28704 10602
rect 28664 10116 28716 10122
rect 28664 10058 28716 10064
rect 28296 9980 28348 9986
rect 28296 9922 28348 9928
rect 28308 6858 28336 9922
rect 28388 9504 28440 9510
rect 28388 9446 28440 9452
rect 28572 9504 28624 9510
rect 28572 9446 28624 9452
rect 28400 8490 28428 9446
rect 28480 9300 28532 9306
rect 28480 9242 28532 9248
rect 28492 9034 28520 9242
rect 28480 9028 28532 9034
rect 28480 8970 28532 8976
rect 28388 8484 28440 8490
rect 28388 8426 28440 8432
rect 28584 8286 28612 9446
rect 28664 9368 28716 9374
rect 28664 9310 28716 9316
rect 28676 8694 28704 9310
rect 28664 8688 28716 8694
rect 28664 8630 28716 8636
rect 28572 8280 28624 8286
rect 28572 8222 28624 8228
rect 28584 7742 28612 8222
rect 28572 7736 28624 7742
rect 28572 7678 28624 7684
rect 28676 7334 28704 8630
rect 28664 7328 28716 7334
rect 28664 7270 28716 7276
rect 28480 7056 28532 7062
rect 28480 6998 28532 7004
rect 28296 6852 28348 6858
rect 28348 6812 28428 6840
rect 28296 6794 28348 6800
rect 28204 6172 28256 6178
rect 28204 6114 28256 6120
rect 28216 5702 28244 6114
rect 28296 6104 28348 6110
rect 28296 6046 28348 6052
rect 28308 5770 28336 6046
rect 28296 5764 28348 5770
rect 28296 5706 28348 5712
rect 28204 5696 28256 5702
rect 28204 5638 28256 5644
rect 28216 5498 28244 5638
rect 28204 5492 28256 5498
rect 28204 5434 28256 5440
rect 27100 5084 27152 5090
rect 27100 5026 27152 5032
rect 28020 5084 28072 5090
rect 28020 5026 28072 5032
rect 27112 4682 27140 5026
rect 27284 5016 27336 5022
rect 27284 4958 27336 4964
rect 27100 4676 27152 4682
rect 27100 4618 27152 4624
rect 27296 4342 27324 4958
rect 28032 4478 28060 5026
rect 28020 4472 28072 4478
rect 28020 4414 28072 4420
rect 27284 4336 27336 4342
rect 27284 4278 27336 4284
rect 27296 3526 27324 4278
rect 28032 4138 28060 4414
rect 28020 4132 28072 4138
rect 28020 4074 28072 4080
rect 27284 3520 27336 3526
rect 27284 3462 27336 3468
rect 26548 3384 26600 3390
rect 26548 3326 26600 3332
rect 26180 3044 26232 3050
rect 26180 2986 26232 2992
rect 26088 2976 26140 2982
rect 26088 2918 26140 2924
rect 26560 2914 26588 3326
rect 26548 2908 26600 2914
rect 26548 2850 26600 2856
rect 26824 2840 26876 2846
rect 26824 2782 26876 2788
rect 25812 2704 25864 2710
rect 25812 2646 25864 2652
rect 25824 2370 25852 2646
rect 26836 2370 26864 2782
rect 27296 2506 27324 3462
rect 28032 2914 28060 4074
rect 28308 3390 28336 5706
rect 28296 3384 28348 3390
rect 28296 3326 28348 3332
rect 28296 3248 28348 3254
rect 28216 3208 28296 3236
rect 28020 2908 28072 2914
rect 28020 2850 28072 2856
rect 27284 2500 27336 2506
rect 27284 2442 27336 2448
rect 27468 2432 27520 2438
rect 27468 2374 27520 2380
rect 25812 2364 25864 2370
rect 25812 2306 25864 2312
rect 26824 2364 26876 2370
rect 26824 2306 26876 2312
rect 27376 2296 27428 2302
rect 27376 2238 27428 2244
rect 25628 2228 25680 2234
rect 25628 2170 25680 2176
rect 27388 1962 27416 2238
rect 27376 1956 27428 1962
rect 27376 1898 27428 1904
rect 26548 1684 26600 1690
rect 26548 1626 26600 1632
rect 25996 1616 26048 1622
rect 25996 1558 26048 1564
rect 26008 1078 26036 1558
rect 25996 1072 26048 1078
rect 25996 1014 26048 1020
rect 26560 424 26588 1626
rect 27480 1418 27508 2374
rect 28032 2302 28060 2850
rect 28216 2438 28244 3208
rect 28296 3190 28348 3196
rect 28204 2432 28256 2438
rect 28204 2374 28256 2380
rect 27744 2296 27796 2302
rect 27744 2238 27796 2244
rect 28020 2296 28072 2302
rect 28020 2238 28072 2244
rect 27756 2166 27784 2238
rect 27836 2228 27888 2234
rect 27836 2170 27888 2176
rect 27744 2160 27796 2166
rect 27744 2102 27796 2108
rect 27756 1622 27784 2102
rect 27848 1826 27876 2170
rect 27836 1820 27888 1826
rect 27836 1762 27888 1768
rect 27744 1616 27796 1622
rect 27744 1558 27796 1564
rect 27468 1412 27520 1418
rect 27468 1354 27520 1360
rect 27756 1350 27784 1558
rect 27848 1418 27876 1762
rect 28032 1758 28060 2238
rect 28216 1894 28244 2374
rect 28400 2234 28428 6812
rect 28492 6586 28520 6998
rect 28480 6580 28532 6586
rect 28480 6522 28532 6528
rect 28676 6518 28704 7270
rect 28768 7198 28796 10942
rect 28952 10682 28980 12098
rect 29044 10852 29072 12982
rect 29136 12774 29164 13798
rect 29308 13380 29360 13386
rect 29308 13322 29360 13328
rect 29124 12768 29176 12774
rect 29124 12710 29176 12716
rect 29216 12088 29268 12094
rect 29216 12030 29268 12036
rect 29124 12020 29176 12026
rect 29124 11962 29176 11968
rect 29136 11686 29164 11962
rect 29124 11680 29176 11686
rect 29124 11622 29176 11628
rect 29136 11074 29164 11622
rect 29228 11550 29256 12030
rect 29320 11686 29348 13322
rect 29584 12088 29636 12094
rect 29584 12030 29636 12036
rect 29308 11680 29360 11686
rect 29308 11622 29360 11628
rect 29216 11544 29268 11550
rect 29216 11486 29268 11492
rect 29320 11210 29348 11622
rect 29596 11482 29624 12030
rect 29676 11544 29728 11550
rect 29676 11486 29728 11492
rect 29584 11476 29636 11482
rect 29584 11418 29636 11424
rect 29308 11204 29360 11210
rect 29308 11146 29360 11152
rect 29124 11068 29176 11074
rect 29124 11010 29176 11016
rect 29308 11068 29360 11074
rect 29308 11010 29360 11016
rect 29124 10864 29176 10870
rect 29044 10824 29124 10852
rect 29124 10806 29176 10812
rect 28952 10654 29072 10682
rect 28848 9436 28900 9442
rect 28848 9378 28900 9384
rect 28860 8830 28888 9378
rect 29044 8966 29072 10654
rect 29136 9442 29164 10806
rect 29216 9912 29268 9918
rect 29216 9854 29268 9860
rect 29124 9436 29176 9442
rect 29124 9378 29176 9384
rect 29136 9034 29164 9378
rect 29228 9034 29256 9854
rect 29124 9028 29176 9034
rect 29124 8970 29176 8976
rect 29216 9028 29268 9034
rect 29216 8970 29268 8976
rect 29032 8960 29084 8966
rect 29032 8902 29084 8908
rect 28848 8824 28900 8830
rect 28848 8766 28900 8772
rect 29216 8756 29268 8762
rect 29216 8698 29268 8704
rect 29228 8354 29256 8698
rect 29216 8348 29268 8354
rect 29216 8290 29268 8296
rect 29228 7946 29256 8290
rect 29216 7940 29268 7946
rect 29216 7882 29268 7888
rect 28756 7192 28808 7198
rect 28756 7134 28808 7140
rect 29320 6722 29348 11010
rect 29688 11006 29716 11486
rect 29676 11000 29728 11006
rect 29676 10942 29728 10948
rect 29780 10530 29808 24066
rect 30056 23586 30084 25455
rect 30596 25076 30648 25082
rect 30596 25018 30648 25024
rect 30608 24198 30636 25018
rect 30596 24192 30648 24198
rect 30596 24134 30648 24140
rect 31528 24130 31556 31664
rect 31516 24124 31568 24130
rect 31516 24066 31568 24072
rect 30228 23648 30280 23654
rect 30134 23616 30190 23625
rect 30044 23580 30096 23586
rect 30228 23590 30280 23596
rect 30134 23551 30190 23560
rect 30044 23522 30096 23528
rect 30056 23110 30084 23522
rect 30148 23110 30176 23551
rect 30044 23104 30096 23110
rect 30044 23046 30096 23052
rect 30136 23104 30188 23110
rect 30136 23046 30188 23052
rect 30240 22838 30268 23590
rect 30412 23512 30464 23518
rect 30412 23454 30464 23460
rect 30424 23178 30452 23454
rect 30412 23172 30464 23178
rect 30412 23114 30464 23120
rect 30228 22832 30280 22838
rect 30228 22774 30280 22780
rect 30240 22022 30268 22774
rect 30228 22016 30280 22022
rect 30228 21958 30280 21964
rect 30136 20248 30188 20254
rect 30136 20190 30188 20196
rect 30044 18072 30096 18078
rect 30044 18014 30096 18020
rect 30056 17738 30084 18014
rect 30044 17732 30096 17738
rect 30044 17674 30096 17680
rect 30056 16446 30084 17674
rect 30044 16440 30096 16446
rect 30044 16382 30096 16388
rect 29952 16304 30004 16310
rect 29952 16246 30004 16252
rect 29860 11612 29912 11618
rect 29860 11554 29912 11560
rect 29872 11210 29900 11554
rect 29860 11204 29912 11210
rect 29860 11146 29912 11152
rect 29768 10524 29820 10530
rect 29768 10466 29820 10472
rect 29676 10320 29728 10326
rect 29676 10262 29728 10268
rect 29688 10074 29716 10262
rect 29584 10048 29636 10054
rect 29688 10046 29808 10074
rect 29584 9990 29636 9996
rect 29596 9918 29624 9990
rect 29780 9918 29808 10046
rect 29584 9912 29636 9918
rect 29584 9854 29636 9860
rect 29768 9912 29820 9918
rect 29768 9854 29820 9860
rect 29964 9209 29992 16246
rect 30148 12638 30176 20190
rect 30502 19536 30558 19545
rect 30502 19471 30558 19480
rect 30516 19234 30544 19471
rect 30504 19228 30556 19234
rect 30504 19170 30556 19176
rect 30516 18826 30544 19170
rect 30504 18820 30556 18826
rect 30504 18762 30556 18768
rect 30502 15456 30558 15465
rect 30502 15391 30558 15400
rect 30516 13833 30544 15391
rect 30502 13824 30558 13833
rect 30502 13759 30558 13768
rect 30136 12632 30188 12638
rect 30136 12574 30188 12580
rect 30148 12094 30176 12574
rect 30136 12088 30188 12094
rect 30136 12030 30188 12036
rect 30228 11544 30280 11550
rect 30228 11486 30280 11492
rect 30044 11476 30096 11482
rect 30044 11418 30096 11424
rect 30056 11210 30084 11418
rect 30044 11204 30096 11210
rect 30044 11146 30096 11152
rect 30240 10938 30268 11486
rect 30228 10932 30280 10938
rect 30228 10874 30280 10880
rect 30044 9300 30096 9306
rect 30044 9242 30096 9248
rect 29950 9200 30006 9209
rect 29950 9135 30006 9144
rect 29400 8824 29452 8830
rect 29400 8766 29452 8772
rect 29412 8490 29440 8766
rect 30056 8490 30084 9242
rect 29400 8484 29452 8490
rect 29400 8426 29452 8432
rect 30044 8484 30096 8490
rect 30044 8426 30096 8432
rect 30056 7946 30084 8426
rect 30044 7940 30096 7946
rect 30044 7882 30096 7888
rect 30502 7296 30558 7305
rect 30502 7231 30558 7240
rect 29584 7124 29636 7130
rect 29584 7066 29636 7072
rect 29308 6716 29360 6722
rect 29308 6658 29360 6664
rect 29216 6648 29268 6654
rect 29216 6590 29268 6596
rect 28940 6580 28992 6586
rect 28940 6522 28992 6528
rect 28664 6512 28716 6518
rect 28664 6454 28716 6460
rect 28848 6512 28900 6518
rect 28848 6454 28900 6460
rect 28676 5208 28704 6454
rect 28860 5974 28888 6454
rect 28848 5968 28900 5974
rect 28848 5910 28900 5916
rect 28756 5492 28808 5498
rect 28756 5434 28808 5440
rect 28768 5401 28796 5434
rect 28754 5392 28810 5401
rect 28754 5327 28810 5336
rect 28756 5220 28808 5226
rect 28676 5180 28756 5208
rect 28756 5162 28808 5168
rect 28768 4410 28796 5162
rect 28756 4404 28808 4410
rect 28756 4346 28808 4352
rect 28664 4336 28716 4342
rect 28664 4278 28716 4284
rect 28676 4138 28704 4278
rect 28664 4132 28716 4138
rect 28664 4074 28716 4080
rect 28676 3236 28704 4074
rect 28756 3928 28808 3934
rect 28756 3870 28808 3876
rect 28768 3594 28796 3870
rect 28756 3588 28808 3594
rect 28756 3530 28808 3536
rect 28756 3248 28808 3254
rect 28676 3208 28756 3236
rect 28756 3190 28808 3196
rect 28768 2982 28796 3190
rect 28756 2976 28808 2982
rect 28756 2918 28808 2924
rect 28860 2846 28888 5910
rect 28952 5022 28980 6522
rect 29228 6314 29256 6590
rect 29216 6308 29268 6314
rect 29216 6250 29268 6256
rect 29320 6246 29348 6658
rect 29596 6654 29624 7066
rect 29584 6648 29636 6654
rect 29584 6590 29636 6596
rect 29308 6240 29360 6246
rect 29308 6182 29360 6188
rect 29308 5492 29360 5498
rect 29308 5434 29360 5440
rect 29124 5152 29176 5158
rect 29124 5094 29176 5100
rect 28940 5016 28992 5022
rect 28940 4958 28992 4964
rect 28952 4682 28980 4958
rect 28940 4676 28992 4682
rect 28940 4618 28992 4624
rect 29136 4070 29164 5094
rect 29124 4064 29176 4070
rect 29124 4006 29176 4012
rect 29216 3520 29268 3526
rect 29216 3462 29268 3468
rect 29228 3390 29256 3462
rect 29320 3390 29348 5434
rect 30516 5265 30544 7231
rect 30502 5256 30558 5265
rect 30502 5191 30558 5200
rect 30504 3792 30556 3798
rect 30504 3734 30556 3740
rect 30516 3390 30544 3734
rect 29216 3384 29268 3390
rect 29216 3326 29268 3332
rect 29308 3384 29360 3390
rect 29308 3326 29360 3332
rect 29584 3384 29636 3390
rect 29584 3326 29636 3332
rect 30504 3384 30556 3390
rect 30504 3326 30556 3332
rect 29596 3254 29624 3326
rect 29584 3248 29636 3254
rect 30516 3225 30544 3326
rect 29584 3190 29636 3196
rect 30502 3216 30558 3225
rect 28848 2840 28900 2846
rect 28848 2782 28900 2788
rect 29308 2840 29360 2846
rect 29308 2782 29360 2788
rect 28860 2506 28888 2782
rect 28848 2500 28900 2506
rect 28848 2442 28900 2448
rect 29320 2234 29348 2782
rect 29596 2370 29624 3190
rect 30502 3151 30558 3160
rect 29584 2364 29636 2370
rect 29584 2306 29636 2312
rect 28388 2228 28440 2234
rect 28388 2170 28440 2176
rect 29308 2228 29360 2234
rect 29308 2170 29360 2176
rect 28204 1888 28256 1894
rect 28204 1830 28256 1836
rect 28020 1752 28072 1758
rect 28020 1694 28072 1700
rect 28032 1418 28060 1694
rect 27836 1412 27888 1418
rect 27836 1354 27888 1360
rect 28020 1412 28072 1418
rect 28020 1354 28072 1360
rect 27744 1344 27796 1350
rect 27744 1286 27796 1292
rect 28018 768 28074 777
rect 28018 703 28074 712
rect 28032 424 28060 703
rect 29320 424 29348 2170
rect 30780 1616 30832 1622
rect 30780 1558 30832 1564
rect 30792 424 30820 1558
rect 12802 384 12830 424
rect 12718 0 12830 384
rect 14190 0 14302 424
rect 15478 0 15590 424
rect 16624 398 17062 424
rect 16950 0 17062 398
rect 18238 0 18350 424
rect 19710 0 19822 424
rect 20998 0 21110 424
rect 22470 0 22582 424
rect 23758 0 23870 424
rect 25230 0 25342 424
rect 26518 0 26630 424
rect 27990 0 28102 424
rect 29278 0 29390 424
rect 30750 0 30862 424
<< via2 >>
rect 418 30904 474 30960
rect 3516 30890 3572 30892
rect 3596 30890 3652 30892
rect 3676 30890 3732 30892
rect 3756 30890 3812 30892
rect 3516 30838 3562 30890
rect 3562 30838 3572 30890
rect 3596 30838 3626 30890
rect 3626 30838 3638 30890
rect 3638 30838 3652 30890
rect 3676 30838 3690 30890
rect 3690 30838 3702 30890
rect 3702 30838 3732 30890
rect 3756 30838 3766 30890
rect 3766 30838 3812 30890
rect 3516 30836 3572 30838
rect 3596 30836 3652 30838
rect 3676 30836 3732 30838
rect 3756 30836 3812 30838
rect 3516 29802 3572 29804
rect 3596 29802 3652 29804
rect 3676 29802 3732 29804
rect 3756 29802 3812 29804
rect 3516 29750 3562 29802
rect 3562 29750 3572 29802
rect 3596 29750 3626 29802
rect 3626 29750 3638 29802
rect 3638 29750 3652 29802
rect 3676 29750 3690 29802
rect 3690 29750 3702 29802
rect 3702 29750 3732 29802
rect 3756 29750 3766 29802
rect 3766 29750 3812 29802
rect 3516 29748 3572 29750
rect 3596 29748 3652 29750
rect 3676 29748 3732 29750
rect 3756 29748 3812 29750
rect 1614 28728 1670 28784
rect 1154 20568 1210 20624
rect 3516 28714 3572 28716
rect 3596 28714 3652 28716
rect 3676 28714 3732 28716
rect 3756 28714 3812 28716
rect 3516 28662 3562 28714
rect 3562 28662 3572 28714
rect 3596 28662 3626 28714
rect 3626 28662 3638 28714
rect 3638 28662 3652 28714
rect 3676 28662 3690 28714
rect 3690 28662 3702 28714
rect 3702 28662 3732 28714
rect 3756 28662 3766 28714
rect 3766 28662 3812 28714
rect 3516 28660 3572 28662
rect 3596 28660 3652 28662
rect 3676 28660 3732 28662
rect 3756 28660 3812 28662
rect 3516 27626 3572 27628
rect 3596 27626 3652 27628
rect 3676 27626 3732 27628
rect 3756 27626 3812 27628
rect 3516 27574 3562 27626
rect 3562 27574 3572 27626
rect 3596 27574 3626 27626
rect 3626 27574 3638 27626
rect 3638 27574 3652 27626
rect 3676 27574 3690 27626
rect 3690 27574 3702 27626
rect 3702 27574 3732 27626
rect 3756 27574 3766 27626
rect 3766 27574 3812 27626
rect 3516 27572 3572 27574
rect 3596 27572 3652 27574
rect 3676 27572 3732 27574
rect 3756 27572 3812 27574
rect 3516 26538 3572 26540
rect 3596 26538 3652 26540
rect 3676 26538 3732 26540
rect 3756 26538 3812 26540
rect 3516 26486 3562 26538
rect 3562 26486 3572 26538
rect 3596 26486 3626 26538
rect 3626 26486 3638 26538
rect 3638 26486 3652 26538
rect 3676 26486 3690 26538
rect 3690 26486 3702 26538
rect 3702 26486 3732 26538
rect 3756 26486 3766 26538
rect 3766 26486 3812 26538
rect 3516 26484 3572 26486
rect 3596 26484 3652 26486
rect 3676 26484 3732 26486
rect 3756 26484 3812 26486
rect 2350 25192 2406 25248
rect 3516 25450 3572 25452
rect 3596 25450 3652 25452
rect 3676 25450 3732 25452
rect 3756 25450 3812 25452
rect 3516 25398 3562 25450
rect 3562 25398 3572 25450
rect 3596 25398 3626 25450
rect 3626 25398 3638 25450
rect 3638 25398 3652 25450
rect 3676 25398 3690 25450
rect 3690 25398 3702 25450
rect 3702 25398 3732 25450
rect 3756 25398 3766 25450
rect 3766 25398 3812 25450
rect 3516 25396 3572 25398
rect 3596 25396 3652 25398
rect 3676 25396 3732 25398
rect 3756 25396 3812 25398
rect 3516 24362 3572 24364
rect 3596 24362 3652 24364
rect 3676 24362 3732 24364
rect 3756 24362 3812 24364
rect 3516 24310 3562 24362
rect 3562 24310 3572 24362
rect 3596 24310 3626 24362
rect 3626 24310 3638 24362
rect 3638 24310 3652 24362
rect 3676 24310 3690 24362
rect 3690 24310 3702 24362
rect 3702 24310 3732 24362
rect 3756 24310 3766 24362
rect 3766 24310 3812 24362
rect 3516 24308 3572 24310
rect 3596 24308 3652 24310
rect 3676 24308 3732 24310
rect 3756 24308 3812 24310
rect 3516 23274 3572 23276
rect 3596 23274 3652 23276
rect 3676 23274 3732 23276
rect 3756 23274 3812 23276
rect 3516 23222 3562 23274
rect 3562 23222 3572 23274
rect 3596 23222 3626 23274
rect 3626 23222 3638 23274
rect 3638 23222 3652 23274
rect 3676 23222 3690 23274
rect 3690 23222 3702 23274
rect 3702 23222 3732 23274
rect 3756 23222 3766 23274
rect 3766 23222 3812 23274
rect 3516 23220 3572 23222
rect 3596 23220 3652 23222
rect 3676 23220 3732 23222
rect 3756 23220 3812 23222
rect 3516 22186 3572 22188
rect 3596 22186 3652 22188
rect 3676 22186 3732 22188
rect 3756 22186 3812 22188
rect 3516 22134 3562 22186
rect 3562 22134 3572 22186
rect 3596 22134 3626 22186
rect 3626 22134 3638 22186
rect 3638 22134 3652 22186
rect 3676 22134 3690 22186
rect 3690 22134 3702 22186
rect 3702 22134 3732 22186
rect 3756 22134 3766 22186
rect 3766 22134 3812 22186
rect 3516 22132 3572 22134
rect 3596 22132 3652 22134
rect 3676 22132 3732 22134
rect 3756 22132 3812 22134
rect 3516 21098 3572 21100
rect 3596 21098 3652 21100
rect 3676 21098 3732 21100
rect 3756 21098 3812 21100
rect 3516 21046 3562 21098
rect 3562 21046 3572 21098
rect 3596 21046 3626 21098
rect 3626 21046 3638 21098
rect 3638 21046 3652 21098
rect 3676 21046 3690 21098
rect 3690 21046 3702 21098
rect 3702 21046 3732 21098
rect 3756 21046 3766 21098
rect 3766 21046 3812 21098
rect 3516 21044 3572 21046
rect 3596 21044 3652 21046
rect 3676 21044 3732 21046
rect 3756 21044 3812 21046
rect 4650 22744 4706 22800
rect 3516 20010 3572 20012
rect 3596 20010 3652 20012
rect 3676 20010 3732 20012
rect 3756 20010 3812 20012
rect 3516 19958 3562 20010
rect 3562 19958 3572 20010
rect 3596 19958 3626 20010
rect 3626 19958 3638 20010
rect 3638 19958 3652 20010
rect 3676 19958 3690 20010
rect 3690 19958 3702 20010
rect 3702 19958 3732 20010
rect 3756 19958 3766 20010
rect 3766 19958 3812 20010
rect 3516 19956 3572 19958
rect 3596 19956 3652 19958
rect 3676 19956 3732 19958
rect 3756 19956 3812 19958
rect 1154 16488 1210 16544
rect 3270 19636 3326 19672
rect 3270 19616 3272 19636
rect 3272 19616 3324 19636
rect 3324 19616 3326 19636
rect 3516 18922 3572 18924
rect 3596 18922 3652 18924
rect 3676 18922 3732 18924
rect 3756 18922 3812 18924
rect 3516 18870 3562 18922
rect 3562 18870 3572 18922
rect 3596 18870 3626 18922
rect 3626 18870 3638 18922
rect 3638 18870 3652 18922
rect 3676 18870 3690 18922
rect 3690 18870 3702 18922
rect 3702 18870 3732 18922
rect 3756 18870 3766 18922
rect 3766 18870 3812 18922
rect 3516 18868 3572 18870
rect 3596 18868 3652 18870
rect 3676 18868 3732 18870
rect 3756 18868 3812 18870
rect 3516 17834 3572 17836
rect 3596 17834 3652 17836
rect 3676 17834 3732 17836
rect 3756 17834 3812 17836
rect 3516 17782 3562 17834
rect 3562 17782 3572 17834
rect 3596 17782 3626 17834
rect 3626 17782 3638 17834
rect 3638 17782 3652 17834
rect 3676 17782 3690 17834
rect 3690 17782 3702 17834
rect 3702 17782 3732 17834
rect 3756 17782 3766 17834
rect 3766 17782 3812 17834
rect 3516 17780 3572 17782
rect 3596 17780 3652 17782
rect 3676 17780 3732 17782
rect 3756 17780 3812 17782
rect 3516 16746 3572 16748
rect 3596 16746 3652 16748
rect 3676 16746 3732 16748
rect 3756 16746 3812 16748
rect 3516 16694 3562 16746
rect 3562 16694 3572 16746
rect 3596 16694 3626 16746
rect 3626 16694 3638 16746
rect 3638 16694 3652 16746
rect 3676 16694 3690 16746
rect 3690 16694 3702 16746
rect 3702 16694 3732 16746
rect 3756 16694 3766 16746
rect 3766 16694 3812 16746
rect 3516 16692 3572 16694
rect 3596 16692 3652 16694
rect 3676 16692 3732 16694
rect 3756 16692 3812 16694
rect 4558 17304 4614 17360
rect 3516 15658 3572 15660
rect 3596 15658 3652 15660
rect 3676 15658 3732 15660
rect 3756 15658 3812 15660
rect 3516 15606 3562 15658
rect 3562 15606 3572 15658
rect 3596 15606 3626 15658
rect 3626 15606 3638 15658
rect 3638 15606 3652 15658
rect 3676 15606 3690 15658
rect 3690 15606 3702 15658
rect 3702 15606 3732 15658
rect 3756 15606 3766 15658
rect 3766 15606 3812 15658
rect 3516 15604 3572 15606
rect 3596 15604 3652 15606
rect 3676 15604 3732 15606
rect 3756 15604 3812 15606
rect 2626 14584 2682 14640
rect 970 12680 1026 12736
rect 3516 14570 3572 14572
rect 3596 14570 3652 14572
rect 3676 14570 3732 14572
rect 3756 14570 3812 14572
rect 3516 14518 3562 14570
rect 3562 14518 3572 14570
rect 3596 14518 3626 14570
rect 3626 14518 3638 14570
rect 3638 14518 3652 14570
rect 3676 14518 3690 14570
rect 3690 14518 3702 14570
rect 3702 14518 3732 14570
rect 3756 14518 3766 14570
rect 3766 14518 3812 14570
rect 3516 14516 3572 14518
rect 3596 14516 3652 14518
rect 3676 14516 3732 14518
rect 3756 14516 3812 14518
rect 4926 19616 4982 19672
rect 6122 20704 6178 20760
rect 5110 18664 5166 18720
rect 3516 13482 3572 13484
rect 3596 13482 3652 13484
rect 3676 13482 3732 13484
rect 3756 13482 3812 13484
rect 3516 13430 3562 13482
rect 3562 13430 3572 13482
rect 3596 13430 3626 13482
rect 3626 13430 3638 13482
rect 3638 13430 3652 13482
rect 3676 13430 3690 13482
rect 3690 13430 3702 13482
rect 3702 13430 3732 13482
rect 3756 13430 3766 13482
rect 3766 13430 3812 13482
rect 3516 13428 3572 13430
rect 3596 13428 3652 13430
rect 3676 13428 3732 13430
rect 3756 13428 3812 13430
rect 2074 12680 2130 12736
rect 1246 12408 1302 12464
rect 1338 11612 1394 11648
rect 1338 11592 1340 11612
rect 1340 11592 1392 11612
rect 1392 11592 1394 11612
rect 1430 10504 1486 10560
rect 3516 12394 3572 12396
rect 3596 12394 3652 12396
rect 3676 12394 3732 12396
rect 3756 12394 3812 12396
rect 3516 12342 3562 12394
rect 3562 12342 3572 12394
rect 3596 12342 3626 12394
rect 3626 12342 3638 12394
rect 3638 12342 3652 12394
rect 3676 12342 3690 12394
rect 3690 12342 3702 12394
rect 3702 12342 3732 12394
rect 3756 12342 3766 12394
rect 3766 12342 3812 12394
rect 3516 12340 3572 12342
rect 3596 12340 3652 12342
rect 3676 12340 3732 12342
rect 3756 12340 3812 12342
rect 3516 11306 3572 11308
rect 3596 11306 3652 11308
rect 3676 11306 3732 11308
rect 3756 11306 3812 11308
rect 3516 11254 3562 11306
rect 3562 11254 3572 11306
rect 3596 11254 3626 11306
rect 3626 11254 3638 11306
rect 3638 11254 3652 11306
rect 3676 11254 3690 11306
rect 3690 11254 3702 11306
rect 3702 11254 3732 11306
rect 3756 11254 3766 11306
rect 3766 11254 3812 11306
rect 3516 11252 3572 11254
rect 3596 11252 3652 11254
rect 3676 11252 3732 11254
rect 3756 11252 3812 11254
rect 3516 10218 3572 10220
rect 3596 10218 3652 10220
rect 3676 10218 3732 10220
rect 3756 10218 3812 10220
rect 3516 10166 3562 10218
rect 3562 10166 3572 10218
rect 3596 10166 3626 10218
rect 3626 10166 3638 10218
rect 3638 10166 3652 10218
rect 3676 10166 3690 10218
rect 3690 10166 3702 10218
rect 3702 10166 3732 10218
rect 3756 10166 3766 10218
rect 3766 10166 3812 10218
rect 3516 10164 3572 10166
rect 3596 10164 3652 10166
rect 3676 10164 3732 10166
rect 3756 10164 3812 10166
rect 3516 9130 3572 9132
rect 3596 9130 3652 9132
rect 3676 9130 3732 9132
rect 3756 9130 3812 9132
rect 3516 9078 3562 9130
rect 3562 9078 3572 9130
rect 3596 9078 3626 9130
rect 3626 9078 3638 9130
rect 3638 9078 3652 9130
rect 3676 9078 3690 9130
rect 3690 9078 3702 9130
rect 3702 9078 3732 9130
rect 3756 9078 3766 9130
rect 3766 9078 3812 9130
rect 3516 9076 3572 9078
rect 3596 9076 3652 9078
rect 3676 9076 3732 9078
rect 3756 9076 3812 9078
rect 878 6424 934 6480
rect 3516 8042 3572 8044
rect 3596 8042 3652 8044
rect 3676 8042 3732 8044
rect 3756 8042 3812 8044
rect 3516 7990 3562 8042
rect 3562 7990 3572 8042
rect 3596 7990 3626 8042
rect 3626 7990 3638 8042
rect 3638 7990 3652 8042
rect 3676 7990 3690 8042
rect 3690 7990 3702 8042
rect 3702 7990 3732 8042
rect 3756 7990 3766 8042
rect 3766 7990 3812 8042
rect 3516 7988 3572 7990
rect 3596 7988 3652 7990
rect 3676 7988 3732 7990
rect 3756 7988 3812 7990
rect 3516 6954 3572 6956
rect 3596 6954 3652 6956
rect 3676 6954 3732 6956
rect 3756 6954 3812 6956
rect 3516 6902 3562 6954
rect 3562 6902 3572 6954
rect 3596 6902 3626 6954
rect 3626 6902 3638 6954
rect 3638 6902 3652 6954
rect 3676 6902 3690 6954
rect 3690 6902 3702 6954
rect 3702 6902 3732 6954
rect 3756 6902 3766 6954
rect 3766 6902 3812 6954
rect 3516 6900 3572 6902
rect 3596 6900 3652 6902
rect 3676 6900 3732 6902
rect 3756 6900 3812 6902
rect 6030 9144 6086 9200
rect 4282 6560 4338 6616
rect 4834 6560 4890 6616
rect 1246 4248 1302 4304
rect 3516 5866 3572 5868
rect 3596 5866 3652 5868
rect 3676 5866 3732 5868
rect 3756 5866 3812 5868
rect 3516 5814 3562 5866
rect 3562 5814 3572 5866
rect 3596 5814 3626 5866
rect 3626 5814 3638 5866
rect 3638 5814 3652 5866
rect 3676 5814 3690 5866
rect 3690 5814 3702 5866
rect 3702 5814 3732 5866
rect 3756 5814 3766 5866
rect 3766 5814 3812 5866
rect 3516 5812 3572 5814
rect 3596 5812 3652 5814
rect 3676 5812 3732 5814
rect 3756 5812 3812 5814
rect 3516 4778 3572 4780
rect 3596 4778 3652 4780
rect 3676 4778 3732 4780
rect 3756 4778 3812 4780
rect 3516 4726 3562 4778
rect 3562 4726 3572 4778
rect 3596 4726 3626 4778
rect 3626 4726 3638 4778
rect 3638 4726 3652 4778
rect 3676 4726 3690 4778
rect 3690 4726 3702 4778
rect 3702 4726 3732 4778
rect 3756 4726 3766 4778
rect 3766 4726 3812 4778
rect 3516 4724 3572 4726
rect 3596 4724 3652 4726
rect 3676 4724 3732 4726
rect 3756 4724 3812 4726
rect 3516 3690 3572 3692
rect 3596 3690 3652 3692
rect 3676 3690 3732 3692
rect 3756 3690 3812 3692
rect 3516 3638 3562 3690
rect 3562 3638 3572 3690
rect 3596 3638 3626 3690
rect 3626 3638 3638 3690
rect 3638 3638 3652 3690
rect 3676 3638 3690 3690
rect 3690 3638 3702 3690
rect 3702 3638 3732 3690
rect 3756 3638 3766 3690
rect 3766 3638 3812 3690
rect 3516 3636 3572 3638
rect 3596 3636 3652 3638
rect 3676 3636 3732 3638
rect 3756 3636 3812 3638
rect 1154 2344 1210 2400
rect 3516 2602 3572 2604
rect 3596 2602 3652 2604
rect 3676 2602 3732 2604
rect 3756 2602 3812 2604
rect 3516 2550 3562 2602
rect 3562 2550 3572 2602
rect 3596 2550 3626 2602
rect 3626 2550 3638 2602
rect 3638 2550 3652 2602
rect 3676 2550 3690 2602
rect 3690 2550 3702 2602
rect 3702 2550 3732 2602
rect 3756 2550 3766 2602
rect 3766 2550 3812 2602
rect 3516 2548 3572 2550
rect 3596 2548 3652 2550
rect 3676 2548 3732 2550
rect 3756 2548 3812 2550
rect 418 576 474 632
rect 3516 1514 3572 1516
rect 3596 1514 3652 1516
rect 3676 1514 3732 1516
rect 3756 1514 3812 1516
rect 3516 1462 3562 1514
rect 3562 1462 3572 1514
rect 3596 1462 3626 1514
rect 3626 1462 3638 1514
rect 3638 1462 3652 1514
rect 3676 1462 3690 1514
rect 3690 1462 3702 1514
rect 3702 1462 3732 1514
rect 3756 1462 3766 1514
rect 3766 1462 3812 1514
rect 3516 1460 3572 1462
rect 3596 1460 3652 1462
rect 3676 1460 3732 1462
rect 3756 1460 3812 1462
rect 5846 8056 5902 8112
rect 5938 7920 5994 7976
rect 7410 10504 7466 10560
rect 8422 17304 8478 17360
rect 8238 14196 8294 14232
rect 8238 14176 8240 14196
rect 8240 14176 8292 14196
rect 8292 14176 8294 14196
rect 8054 13632 8110 13688
rect 7686 8328 7742 8384
rect 9618 25192 9674 25248
rect 10262 23832 10318 23888
rect 8606 9416 8662 9472
rect 8882 7240 8938 7296
rect 3516 426 3572 428
rect 3596 426 3652 428
rect 3676 426 3732 428
rect 3756 426 3812 428
rect 3516 374 3562 426
rect 3562 374 3572 426
rect 3596 374 3626 426
rect 3626 374 3638 426
rect 3638 374 3652 426
rect 3676 374 3690 426
rect 3690 374 3702 426
rect 3702 374 3732 426
rect 3756 374 3766 426
rect 3766 374 3812 426
rect 5938 712 5994 768
rect 9894 12680 9950 12736
rect 9986 12000 10042 12056
rect 9710 11320 9766 11376
rect 10170 10912 10226 10968
rect 12010 23832 12066 23888
rect 10814 10096 10870 10152
rect 12562 23868 12564 23888
rect 12564 23868 12616 23888
rect 12616 23868 12618 23888
rect 12562 23832 12618 23868
rect 13298 24648 13354 24704
rect 13666 29680 13722 29736
rect 16518 29408 16574 29464
rect 18876 31434 18932 31436
rect 18956 31434 19012 31436
rect 19036 31434 19092 31436
rect 19116 31434 19172 31436
rect 18876 31382 18922 31434
rect 18922 31382 18932 31434
rect 18956 31382 18986 31434
rect 18986 31382 18998 31434
rect 18998 31382 19012 31434
rect 19036 31382 19050 31434
rect 19050 31382 19062 31434
rect 19062 31382 19092 31434
rect 19116 31382 19126 31434
rect 19126 31382 19172 31434
rect 18876 31380 18932 31382
rect 18956 31380 19012 31382
rect 19036 31380 19092 31382
rect 19116 31380 19172 31382
rect 12746 9824 12802 9880
rect 12010 9280 12066 9336
rect 18876 30346 18932 30348
rect 18956 30346 19012 30348
rect 19036 30346 19092 30348
rect 19116 30346 19172 30348
rect 18876 30294 18922 30346
rect 18922 30294 18932 30346
rect 18956 30294 18986 30346
rect 18986 30294 18998 30346
rect 18998 30294 19012 30346
rect 19036 30294 19050 30346
rect 19050 30294 19062 30346
rect 19062 30294 19092 30346
rect 19116 30294 19126 30346
rect 19126 30294 19172 30346
rect 18876 30292 18932 30294
rect 18956 30292 19012 30294
rect 19036 30292 19092 30294
rect 19116 30292 19172 30294
rect 16518 20704 16574 20760
rect 19554 29680 19610 29736
rect 18876 29258 18932 29260
rect 18956 29258 19012 29260
rect 19036 29258 19092 29260
rect 19116 29258 19172 29260
rect 18876 29206 18922 29258
rect 18922 29206 18932 29258
rect 18956 29206 18986 29258
rect 18986 29206 18998 29258
rect 18998 29206 19012 29258
rect 19036 29206 19050 29258
rect 19050 29206 19062 29258
rect 19062 29206 19092 29258
rect 19116 29206 19126 29258
rect 19126 29206 19172 29258
rect 18876 29204 18932 29206
rect 18956 29204 19012 29206
rect 19036 29204 19092 29206
rect 19116 29204 19172 29206
rect 18876 28170 18932 28172
rect 18956 28170 19012 28172
rect 19036 28170 19092 28172
rect 19116 28170 19172 28172
rect 18876 28118 18922 28170
rect 18922 28118 18932 28170
rect 18956 28118 18986 28170
rect 18986 28118 18998 28170
rect 18998 28118 19012 28170
rect 19036 28118 19050 28170
rect 19050 28118 19062 28170
rect 19062 28118 19092 28170
rect 19116 28118 19126 28170
rect 19126 28118 19172 28170
rect 18876 28116 18932 28118
rect 18956 28116 19012 28118
rect 19036 28116 19092 28118
rect 19116 28116 19172 28118
rect 18876 27082 18932 27084
rect 18956 27082 19012 27084
rect 19036 27082 19092 27084
rect 19116 27082 19172 27084
rect 18876 27030 18922 27082
rect 18922 27030 18932 27082
rect 18956 27030 18986 27082
rect 18986 27030 18998 27082
rect 18998 27030 19012 27082
rect 19036 27030 19050 27082
rect 19050 27030 19062 27082
rect 19062 27030 19092 27082
rect 19116 27030 19126 27082
rect 19126 27030 19172 27082
rect 18876 27028 18932 27030
rect 18956 27028 19012 27030
rect 19036 27028 19092 27030
rect 19116 27028 19172 27030
rect 18876 25994 18932 25996
rect 18956 25994 19012 25996
rect 19036 25994 19092 25996
rect 19116 25994 19172 25996
rect 18876 25942 18922 25994
rect 18922 25942 18932 25994
rect 18956 25942 18986 25994
rect 18986 25942 18998 25994
rect 18998 25942 19012 25994
rect 19036 25942 19050 25994
rect 19050 25942 19062 25994
rect 19062 25942 19092 25994
rect 19116 25942 19126 25994
rect 19126 25942 19172 25994
rect 18876 25940 18932 25942
rect 18956 25940 19012 25942
rect 19036 25940 19092 25942
rect 19116 25940 19172 25942
rect 18876 24906 18932 24908
rect 18956 24906 19012 24908
rect 19036 24906 19092 24908
rect 19116 24906 19172 24908
rect 18876 24854 18922 24906
rect 18922 24854 18932 24906
rect 18956 24854 18986 24906
rect 18986 24854 18998 24906
rect 18998 24854 19012 24906
rect 19036 24854 19050 24906
rect 19050 24854 19062 24906
rect 19062 24854 19092 24906
rect 19116 24854 19126 24906
rect 19126 24854 19172 24906
rect 18876 24852 18932 24854
rect 18956 24852 19012 24854
rect 19036 24852 19092 24854
rect 19116 24852 19172 24854
rect 18876 23818 18932 23820
rect 18956 23818 19012 23820
rect 19036 23818 19092 23820
rect 19116 23818 19172 23820
rect 18876 23766 18922 23818
rect 18922 23766 18932 23818
rect 18956 23766 18986 23818
rect 18986 23766 18998 23818
rect 18998 23766 19012 23818
rect 19036 23766 19050 23818
rect 19050 23766 19062 23818
rect 19062 23766 19092 23818
rect 19116 23766 19126 23818
rect 19126 23766 19172 23818
rect 18876 23764 18932 23766
rect 18956 23764 19012 23766
rect 19036 23764 19092 23766
rect 19116 23764 19172 23766
rect 18876 22730 18932 22732
rect 18956 22730 19012 22732
rect 19036 22730 19092 22732
rect 19116 22730 19172 22732
rect 18876 22678 18922 22730
rect 18922 22678 18932 22730
rect 18956 22678 18986 22730
rect 18986 22678 18998 22730
rect 18998 22678 19012 22730
rect 19036 22678 19050 22730
rect 19050 22678 19062 22730
rect 19062 22678 19092 22730
rect 19116 22678 19126 22730
rect 19126 22678 19172 22730
rect 18876 22676 18932 22678
rect 18956 22676 19012 22678
rect 19036 22676 19092 22678
rect 19116 22676 19172 22678
rect 18876 21642 18932 21644
rect 18956 21642 19012 21644
rect 19036 21642 19092 21644
rect 19116 21642 19172 21644
rect 18876 21590 18922 21642
rect 18922 21590 18932 21642
rect 18956 21590 18986 21642
rect 18986 21590 18998 21642
rect 18998 21590 19012 21642
rect 19036 21590 19050 21642
rect 19050 21590 19062 21642
rect 19062 21590 19092 21642
rect 19116 21590 19126 21642
rect 19126 21590 19172 21642
rect 18876 21588 18932 21590
rect 18956 21588 19012 21590
rect 19036 21588 19092 21590
rect 19116 21588 19172 21590
rect 18876 20554 18932 20556
rect 18956 20554 19012 20556
rect 19036 20554 19092 20556
rect 19116 20554 19172 20556
rect 18876 20502 18922 20554
rect 18922 20502 18932 20554
rect 18956 20502 18986 20554
rect 18986 20502 18998 20554
rect 18998 20502 19012 20554
rect 19036 20502 19050 20554
rect 19050 20502 19062 20554
rect 19062 20502 19092 20554
rect 19116 20502 19126 20554
rect 19126 20502 19172 20554
rect 18876 20500 18932 20502
rect 18956 20500 19012 20502
rect 19036 20500 19092 20502
rect 19116 20500 19172 20502
rect 10998 3296 11054 3352
rect 11734 3704 11790 3760
rect 12562 3432 12618 3488
rect 3516 372 3572 374
rect 3596 372 3652 374
rect 3676 372 3732 374
rect 3756 372 3812 374
rect 12746 384 12802 440
rect 17346 13768 17402 13824
rect 18876 19466 18932 19468
rect 18956 19466 19012 19468
rect 19036 19466 19092 19468
rect 19116 19466 19172 19468
rect 18876 19414 18922 19466
rect 18922 19414 18932 19466
rect 18956 19414 18986 19466
rect 18986 19414 18998 19466
rect 18998 19414 19012 19466
rect 19036 19414 19050 19466
rect 19050 19414 19062 19466
rect 19062 19414 19092 19466
rect 19116 19414 19126 19466
rect 19126 19414 19172 19466
rect 18876 19412 18932 19414
rect 18956 19412 19012 19414
rect 19036 19412 19092 19414
rect 19116 19412 19172 19414
rect 18876 18378 18932 18380
rect 18956 18378 19012 18380
rect 19036 18378 19092 18380
rect 19116 18378 19172 18380
rect 18876 18326 18922 18378
rect 18922 18326 18932 18378
rect 18956 18326 18986 18378
rect 18986 18326 18998 18378
rect 18998 18326 19012 18378
rect 19036 18326 19050 18378
rect 19050 18326 19062 18378
rect 19062 18326 19092 18378
rect 19116 18326 19126 18378
rect 19126 18326 19172 18378
rect 18876 18324 18932 18326
rect 18956 18324 19012 18326
rect 19036 18324 19092 18326
rect 19116 18324 19172 18326
rect 18876 17290 18932 17292
rect 18956 17290 19012 17292
rect 19036 17290 19092 17292
rect 19116 17290 19172 17292
rect 18876 17238 18922 17290
rect 18922 17238 18932 17290
rect 18956 17238 18986 17290
rect 18986 17238 18998 17290
rect 18998 17238 19012 17290
rect 19036 17238 19050 17290
rect 19050 17238 19062 17290
rect 19062 17238 19092 17290
rect 19116 17238 19126 17290
rect 19126 17238 19172 17290
rect 18876 17236 18932 17238
rect 18956 17236 19012 17238
rect 19036 17236 19092 17238
rect 19116 17236 19172 17238
rect 18876 16202 18932 16204
rect 18956 16202 19012 16204
rect 19036 16202 19092 16204
rect 19116 16202 19172 16204
rect 18876 16150 18922 16202
rect 18922 16150 18932 16202
rect 18956 16150 18986 16202
rect 18986 16150 18998 16202
rect 18998 16150 19012 16202
rect 19036 16150 19050 16202
rect 19050 16150 19062 16202
rect 19062 16150 19092 16202
rect 19116 16150 19126 16202
rect 19126 16150 19172 16202
rect 18876 16148 18932 16150
rect 18956 16148 19012 16150
rect 19036 16148 19092 16150
rect 19116 16148 19172 16150
rect 18876 15114 18932 15116
rect 18956 15114 19012 15116
rect 19036 15114 19092 15116
rect 19116 15114 19172 15116
rect 18876 15062 18922 15114
rect 18922 15062 18932 15114
rect 18956 15062 18986 15114
rect 18986 15062 18998 15114
rect 18998 15062 19012 15114
rect 19036 15062 19050 15114
rect 19050 15062 19062 15114
rect 19062 15062 19092 15114
rect 19116 15062 19126 15114
rect 19126 15062 19172 15114
rect 18876 15060 18932 15062
rect 18956 15060 19012 15062
rect 19036 15060 19092 15062
rect 19116 15060 19172 15062
rect 18876 14026 18932 14028
rect 18956 14026 19012 14028
rect 19036 14026 19092 14028
rect 19116 14026 19172 14028
rect 18876 13974 18922 14026
rect 18922 13974 18932 14026
rect 18956 13974 18986 14026
rect 18986 13974 18998 14026
rect 18998 13974 19012 14026
rect 19036 13974 19050 14026
rect 19050 13974 19062 14026
rect 19062 13974 19092 14026
rect 19116 13974 19126 14026
rect 19126 13974 19172 14026
rect 18876 13972 18932 13974
rect 18956 13972 19012 13974
rect 19036 13972 19092 13974
rect 19116 13972 19172 13974
rect 18876 12938 18932 12940
rect 18956 12938 19012 12940
rect 19036 12938 19092 12940
rect 19116 12938 19172 12940
rect 18876 12886 18922 12938
rect 18922 12886 18932 12938
rect 18956 12886 18986 12938
rect 18986 12886 18998 12938
rect 18998 12886 19012 12938
rect 19036 12886 19050 12938
rect 19050 12886 19062 12938
rect 19062 12886 19092 12938
rect 19116 12886 19126 12938
rect 19126 12886 19172 12938
rect 18876 12884 18932 12886
rect 18956 12884 19012 12886
rect 19036 12884 19092 12886
rect 19116 12884 19172 12886
rect 18876 11850 18932 11852
rect 18956 11850 19012 11852
rect 19036 11850 19092 11852
rect 19116 11850 19172 11852
rect 18876 11798 18922 11850
rect 18922 11798 18932 11850
rect 18956 11798 18986 11850
rect 18986 11798 18998 11850
rect 18998 11798 19012 11850
rect 19036 11798 19050 11850
rect 19050 11798 19062 11850
rect 19062 11798 19092 11850
rect 19116 11798 19126 11850
rect 19126 11798 19172 11850
rect 18876 11796 18932 11798
rect 18956 11796 19012 11798
rect 19036 11796 19092 11798
rect 19116 11796 19172 11798
rect 18876 10762 18932 10764
rect 18956 10762 19012 10764
rect 19036 10762 19092 10764
rect 19116 10762 19172 10764
rect 18876 10710 18922 10762
rect 18922 10710 18932 10762
rect 18956 10710 18986 10762
rect 18986 10710 18998 10762
rect 18998 10710 19012 10762
rect 19036 10710 19050 10762
rect 19050 10710 19062 10762
rect 19062 10710 19092 10762
rect 19116 10710 19126 10762
rect 19126 10710 19172 10762
rect 18876 10708 18932 10710
rect 18956 10708 19012 10710
rect 19036 10708 19092 10710
rect 19116 10708 19172 10710
rect 16334 5608 16390 5664
rect 18266 9416 18322 9472
rect 17806 8192 17862 8248
rect 18876 9674 18932 9676
rect 18956 9674 19012 9676
rect 19036 9674 19092 9676
rect 19116 9674 19172 9676
rect 18876 9622 18922 9674
rect 18922 9622 18932 9674
rect 18956 9622 18986 9674
rect 18986 9622 18998 9674
rect 18998 9622 19012 9674
rect 19036 9622 19050 9674
rect 19050 9622 19062 9674
rect 19062 9622 19092 9674
rect 19116 9622 19126 9674
rect 19126 9622 19172 9674
rect 18876 9620 18932 9622
rect 18956 9620 19012 9622
rect 19036 9620 19092 9622
rect 19116 9620 19172 9622
rect 18450 9416 18506 9472
rect 18876 8586 18932 8588
rect 18956 8586 19012 8588
rect 19036 8586 19092 8588
rect 19116 8586 19172 8588
rect 18876 8534 18922 8586
rect 18922 8534 18932 8586
rect 18956 8534 18986 8586
rect 18986 8534 18998 8586
rect 18998 8534 19012 8586
rect 19036 8534 19050 8586
rect 19050 8534 19062 8586
rect 19062 8534 19092 8586
rect 19116 8534 19126 8586
rect 19126 8534 19172 8586
rect 18876 8532 18932 8534
rect 18956 8532 19012 8534
rect 19036 8532 19092 8534
rect 19116 8532 19172 8534
rect 18876 7498 18932 7500
rect 18956 7498 19012 7500
rect 19036 7498 19092 7500
rect 19116 7498 19172 7500
rect 18876 7446 18922 7498
rect 18922 7446 18932 7498
rect 18956 7446 18986 7498
rect 18986 7446 18998 7498
rect 18998 7446 19012 7498
rect 19036 7446 19050 7498
rect 19050 7446 19062 7498
rect 19062 7446 19092 7498
rect 19116 7446 19126 7498
rect 19126 7446 19172 7498
rect 18876 7444 18932 7446
rect 18956 7444 19012 7446
rect 19036 7444 19092 7446
rect 19116 7444 19172 7446
rect 18876 6410 18932 6412
rect 18956 6410 19012 6412
rect 19036 6410 19092 6412
rect 19116 6410 19172 6412
rect 18876 6358 18922 6410
rect 18922 6358 18932 6410
rect 18956 6358 18986 6410
rect 18986 6358 18998 6410
rect 18998 6358 19012 6410
rect 19036 6358 19050 6410
rect 19050 6358 19062 6410
rect 19062 6358 19092 6410
rect 19116 6358 19126 6410
rect 19126 6358 19172 6410
rect 18876 6356 18932 6358
rect 18956 6356 19012 6358
rect 19036 6356 19092 6358
rect 19116 6356 19172 6358
rect 18876 5322 18932 5324
rect 18956 5322 19012 5324
rect 19036 5322 19092 5324
rect 19116 5322 19172 5324
rect 18876 5270 18922 5322
rect 18922 5270 18932 5322
rect 18956 5270 18986 5322
rect 18986 5270 18998 5322
rect 18998 5270 19012 5322
rect 19036 5270 19050 5322
rect 19050 5270 19062 5322
rect 19062 5270 19092 5322
rect 19116 5270 19126 5322
rect 19126 5270 19172 5322
rect 18876 5268 18932 5270
rect 18956 5268 19012 5270
rect 19036 5268 19092 5270
rect 19116 5268 19172 5270
rect 18634 4520 18690 4576
rect 19370 5336 19426 5392
rect 19278 4520 19334 4576
rect 18876 4234 18932 4236
rect 18956 4234 19012 4236
rect 19036 4234 19092 4236
rect 19116 4234 19172 4236
rect 18876 4182 18922 4234
rect 18922 4182 18932 4234
rect 18956 4182 18986 4234
rect 18986 4182 18998 4234
rect 18998 4182 19012 4234
rect 19036 4182 19050 4234
rect 19050 4182 19062 4234
rect 19062 4182 19092 4234
rect 19116 4182 19126 4234
rect 19126 4182 19172 4234
rect 18876 4180 18932 4182
rect 18956 4180 19012 4182
rect 19036 4180 19092 4182
rect 19116 4180 19172 4182
rect 18876 3146 18932 3148
rect 18956 3146 19012 3148
rect 19036 3146 19092 3148
rect 19116 3146 19172 3148
rect 18876 3094 18922 3146
rect 18922 3094 18932 3146
rect 18956 3094 18986 3146
rect 18986 3094 18998 3146
rect 18998 3094 19012 3146
rect 19036 3094 19050 3146
rect 19050 3094 19062 3146
rect 19062 3094 19092 3146
rect 19116 3094 19126 3146
rect 19126 3094 19172 3146
rect 18876 3092 18932 3094
rect 18956 3092 19012 3094
rect 19036 3092 19092 3094
rect 19116 3092 19172 3094
rect 17714 712 17770 768
rect 18876 2058 18932 2060
rect 18956 2058 19012 2060
rect 19036 2058 19092 2060
rect 19116 2058 19172 2060
rect 18876 2006 18922 2058
rect 18922 2006 18932 2058
rect 18956 2006 18986 2058
rect 18986 2006 18998 2058
rect 18998 2006 19012 2058
rect 19036 2006 19050 2058
rect 19050 2006 19062 2058
rect 19062 2006 19092 2058
rect 19116 2006 19126 2058
rect 19126 2006 19172 2058
rect 18876 2004 18932 2006
rect 18956 2004 19012 2006
rect 19036 2004 19092 2006
rect 19116 2004 19172 2006
rect 18876 970 18932 972
rect 18956 970 19012 972
rect 19036 970 19092 972
rect 19116 970 19172 972
rect 18876 918 18922 970
rect 18922 918 18932 970
rect 18956 918 18986 970
rect 18986 918 18998 970
rect 18998 918 19012 970
rect 19036 918 19050 970
rect 19050 918 19062 970
rect 19062 918 19092 970
rect 19116 918 19126 970
rect 19126 918 19172 970
rect 18876 916 18932 918
rect 18956 916 19012 918
rect 19036 916 19092 918
rect 19116 916 19172 918
rect 20382 9824 20438 9880
rect 20566 12000 20622 12056
rect 20658 11320 20714 11376
rect 20658 9824 20714 9880
rect 20658 9144 20714 9200
rect 20566 7240 20622 7296
rect 19646 3704 19702 3760
rect 20474 3704 20530 3760
rect 19554 712 19610 768
rect 25350 29408 25406 29464
rect 23050 12680 23106 12736
rect 23970 10912 24026 10968
rect 22958 10504 23014 10560
rect 23142 9280 23198 9336
rect 24062 9824 24118 9880
rect 23786 8056 23842 8112
rect 23878 7920 23934 7976
rect 24338 9416 24394 9472
rect 21486 4520 21542 4576
rect 22222 5200 22278 5256
rect 23418 3296 23474 3352
rect 25534 15264 25590 15320
rect 27098 21384 27154 21440
rect 26914 17304 26970 17360
rect 23786 3296 23842 3352
rect 25718 10096 25774 10152
rect 26270 13632 26326 13688
rect 25902 8228 25904 8248
rect 25904 8228 25956 8248
rect 25956 8228 25958 8248
rect 25902 8192 25958 8228
rect 28754 26688 28810 26744
rect 27834 15264 27890 15320
rect 28570 14176 28626 14232
rect 29950 29544 30006 29600
rect 30042 27640 30098 27696
rect 30042 25464 30098 25520
rect 28846 11456 28902 11512
rect 20934 576 20990 632
rect 20566 440 20622 496
rect 20750 440 20806 496
rect 26546 5608 26602 5664
rect 25442 3432 25498 3488
rect 30134 23560 30190 23616
rect 30502 19480 30558 19536
rect 30502 15400 30558 15456
rect 30502 13768 30558 13824
rect 29950 9144 30006 9200
rect 30502 7240 30558 7296
rect 28754 5336 28810 5392
rect 30502 5200 30558 5256
rect 30502 3160 30558 3216
rect 28018 712 28074 768
<< metal3 >>
rect 18864 31440 19184 31456
rect 18864 31376 18872 31440
rect 18936 31376 18952 31440
rect 19016 31376 19032 31440
rect 19096 31376 19112 31440
rect 19176 31376 19184 31440
rect 18864 31360 19184 31376
rect 0 30965 440 31052
rect 0 30962 479 30965
rect 0 30960 580 30962
rect 0 30904 418 30960
rect 474 30904 580 30960
rect 0 30902 580 30904
rect 0 30899 479 30902
rect 0 30812 440 30899
rect 3504 30896 3824 30912
rect 3504 30832 3512 30896
rect 3576 30832 3592 30896
rect 3656 30832 3672 30896
rect 3736 30832 3752 30896
rect 3816 30832 3824 30896
rect 3504 30816 3824 30832
rect 18864 30352 19184 30368
rect 18864 30288 18872 30352
rect 18936 30288 18952 30352
rect 19016 30288 19032 30352
rect 19096 30288 19112 30352
rect 19176 30288 19184 30352
rect 18864 30272 19184 30288
rect 3504 29808 3824 29824
rect 3504 29744 3512 29808
rect 3576 29744 3592 29808
rect 3656 29744 3672 29808
rect 3736 29744 3752 29808
rect 3816 29744 3824 29808
rect 3504 29728 3824 29744
rect 13661 29738 13727 29741
rect 19549 29738 19615 29741
rect 13661 29736 19615 29738
rect 13661 29680 13666 29736
rect 13722 29680 19554 29736
rect 19610 29680 19615 29736
rect 13661 29678 19615 29680
rect 13661 29675 13727 29678
rect 19549 29675 19615 29678
rect 29945 29602 30011 29605
rect 31648 29602 32088 29692
rect 29945 29600 32088 29602
rect 29945 29544 29950 29600
rect 30006 29544 32088 29600
rect 29945 29542 32088 29544
rect 29945 29539 30011 29542
rect 16513 29466 16579 29469
rect 25345 29466 25411 29469
rect 16513 29464 25411 29466
rect 16513 29408 16518 29464
rect 16574 29408 25350 29464
rect 25406 29408 25411 29464
rect 31648 29452 32088 29542
rect 16513 29406 25411 29408
rect 16513 29403 16579 29406
rect 25345 29403 25411 29406
rect 18864 29264 19184 29280
rect 18864 29200 18872 29264
rect 18936 29200 18952 29264
rect 19016 29200 19032 29264
rect 19096 29200 19112 29264
rect 19176 29200 19184 29264
rect 18864 29184 19184 29200
rect 0 28786 440 28876
rect 1609 28786 1675 28789
rect 0 28784 1675 28786
rect 0 28728 1614 28784
rect 1670 28728 1675 28784
rect 0 28726 1675 28728
rect 0 28636 440 28726
rect 1609 28723 1675 28726
rect 3504 28720 3824 28736
rect 3504 28656 3512 28720
rect 3576 28656 3592 28720
rect 3656 28656 3672 28720
rect 3736 28656 3752 28720
rect 3816 28656 3824 28720
rect 3504 28640 3824 28656
rect 18864 28176 19184 28192
rect 18864 28112 18872 28176
rect 18936 28112 18952 28176
rect 19016 28112 19032 28176
rect 19096 28112 19112 28176
rect 19176 28112 19184 28176
rect 18864 28096 19184 28112
rect 30037 27698 30103 27701
rect 31648 27698 32088 27788
rect 30037 27696 32088 27698
rect 3504 27632 3824 27648
rect 30037 27640 30042 27696
rect 30098 27640 32088 27696
rect 30037 27638 32088 27640
rect 30037 27635 30103 27638
rect 3504 27568 3512 27632
rect 3576 27568 3592 27632
rect 3656 27568 3672 27632
rect 3736 27568 3752 27632
rect 3816 27568 3824 27632
rect 3504 27552 3824 27568
rect 31648 27548 32088 27638
rect 18864 27088 19184 27104
rect 18864 27024 18872 27088
rect 18936 27024 18952 27088
rect 19016 27024 19032 27088
rect 19096 27024 19112 27088
rect 19176 27024 19184 27088
rect 18864 27008 19184 27024
rect 0 26882 440 26972
rect 0 26822 4570 26882
rect 0 26732 440 26822
rect 4510 26746 4570 26822
rect 28749 26746 28815 26749
rect 4510 26744 28815 26746
rect 4510 26688 28754 26744
rect 28810 26688 28815 26744
rect 4510 26686 28815 26688
rect 28749 26683 28815 26686
rect 3504 26544 3824 26560
rect 3504 26480 3512 26544
rect 3576 26480 3592 26544
rect 3656 26480 3672 26544
rect 3736 26480 3752 26544
rect 3816 26480 3824 26544
rect 3504 26464 3824 26480
rect 18864 26000 19184 26016
rect 18864 25936 18872 26000
rect 18936 25936 18952 26000
rect 19016 25936 19032 26000
rect 19096 25936 19112 26000
rect 19176 25936 19184 26000
rect 18864 25920 19184 25936
rect 30037 25522 30103 25525
rect 31648 25522 32088 25612
rect 30037 25520 32088 25522
rect 3504 25456 3824 25472
rect 30037 25464 30042 25520
rect 30098 25464 32088 25520
rect 30037 25462 32088 25464
rect 30037 25459 30103 25462
rect 3504 25392 3512 25456
rect 3576 25392 3592 25456
rect 3656 25392 3672 25456
rect 3736 25392 3752 25456
rect 3816 25392 3824 25456
rect 3504 25376 3824 25392
rect 31648 25372 32088 25462
rect 2345 25250 2411 25253
rect 9613 25250 9679 25253
rect 2345 25248 9679 25250
rect 2345 25192 2350 25248
rect 2406 25192 9618 25248
rect 9674 25192 9679 25248
rect 2345 25190 9679 25192
rect 2345 25187 2411 25190
rect 9613 25187 9679 25190
rect 18864 24912 19184 24928
rect 18864 24848 18872 24912
rect 18936 24848 18952 24912
rect 19016 24848 19032 24912
rect 19096 24848 19112 24912
rect 19176 24848 19184 24912
rect 18864 24832 19184 24848
rect 0 24706 440 24796
rect 13293 24706 13359 24709
rect 0 24704 13359 24706
rect 0 24648 13298 24704
rect 13354 24648 13359 24704
rect 0 24646 13359 24648
rect 0 24556 440 24646
rect 13293 24643 13359 24646
rect 3504 24368 3824 24384
rect 3504 24304 3512 24368
rect 3576 24304 3592 24368
rect 3656 24304 3672 24368
rect 3736 24304 3752 24368
rect 3816 24304 3824 24368
rect 3504 24288 3824 24304
rect 10257 23890 10323 23893
rect 12005 23890 12071 23893
rect 12557 23890 12623 23893
rect 10257 23888 12623 23890
rect 10257 23832 10262 23888
rect 10318 23832 12010 23888
rect 12066 23832 12562 23888
rect 12618 23832 12623 23888
rect 10257 23830 12623 23832
rect 10257 23827 10323 23830
rect 12005 23827 12071 23830
rect 12557 23827 12623 23830
rect 18864 23824 19184 23840
rect 18864 23760 18872 23824
rect 18936 23760 18952 23824
rect 19016 23760 19032 23824
rect 19096 23760 19112 23824
rect 19176 23760 19184 23824
rect 18864 23744 19184 23760
rect 30129 23618 30195 23621
rect 31648 23618 32088 23708
rect 30129 23616 32088 23618
rect 30129 23560 30134 23616
rect 30190 23560 32088 23616
rect 30129 23558 32088 23560
rect 30129 23555 30195 23558
rect 31648 23468 32088 23558
rect 3504 23280 3824 23296
rect 3504 23216 3512 23280
rect 3576 23216 3592 23280
rect 3656 23216 3672 23280
rect 3736 23216 3752 23280
rect 3816 23216 3824 23280
rect 3504 23200 3824 23216
rect 0 22802 440 22892
rect 4645 22802 4711 22805
rect 0 22800 4711 22802
rect 0 22744 4650 22800
rect 4706 22744 4711 22800
rect 0 22742 4711 22744
rect 0 22652 440 22742
rect 4645 22739 4711 22742
rect 18864 22736 19184 22752
rect 18864 22672 18872 22736
rect 18936 22672 18952 22736
rect 19016 22672 19032 22736
rect 19096 22672 19112 22736
rect 19176 22672 19184 22736
rect 18864 22656 19184 22672
rect 3504 22192 3824 22208
rect 3504 22128 3512 22192
rect 3576 22128 3592 22192
rect 3656 22128 3672 22192
rect 3736 22128 3752 22192
rect 3816 22128 3824 22192
rect 3504 22112 3824 22128
rect 18864 21648 19184 21664
rect 18864 21584 18872 21648
rect 18936 21584 18952 21648
rect 19016 21584 19032 21648
rect 19096 21584 19112 21648
rect 19176 21584 19184 21648
rect 18864 21568 19184 21584
rect 27093 21442 27159 21445
rect 31648 21442 32088 21532
rect 27093 21440 32088 21442
rect 27093 21384 27098 21440
rect 27154 21384 32088 21440
rect 27093 21382 32088 21384
rect 27093 21379 27159 21382
rect 31648 21292 32088 21382
rect 3504 21104 3824 21120
rect 3504 21040 3512 21104
rect 3576 21040 3592 21104
rect 3656 21040 3672 21104
rect 3736 21040 3752 21104
rect 3816 21040 3824 21104
rect 3504 21024 3824 21040
rect 6117 20762 6183 20765
rect 16513 20762 16579 20765
rect 6117 20760 16579 20762
rect 0 20626 440 20716
rect 6117 20704 6122 20760
rect 6178 20704 16518 20760
rect 16574 20704 16579 20760
rect 6117 20702 16579 20704
rect 6117 20699 6183 20702
rect 16513 20699 16579 20702
rect 1149 20626 1215 20629
rect 0 20624 1215 20626
rect 0 20568 1154 20624
rect 1210 20568 1215 20624
rect 0 20566 1215 20568
rect 0 20476 440 20566
rect 1149 20563 1215 20566
rect 18864 20560 19184 20576
rect 18864 20496 18872 20560
rect 18936 20496 18952 20560
rect 19016 20496 19032 20560
rect 19096 20496 19112 20560
rect 19176 20496 19184 20560
rect 18864 20480 19184 20496
rect 3504 20016 3824 20032
rect 3504 19952 3512 20016
rect 3576 19952 3592 20016
rect 3656 19952 3672 20016
rect 3736 19952 3752 20016
rect 3816 19952 3824 20016
rect 3504 19936 3824 19952
rect 3265 19674 3331 19677
rect 4921 19674 4987 19677
rect 3265 19672 4987 19674
rect 3265 19616 3270 19672
rect 3326 19616 4926 19672
rect 4982 19616 4987 19672
rect 3265 19614 4987 19616
rect 3265 19611 3331 19614
rect 4921 19611 4987 19614
rect 30497 19538 30563 19541
rect 31648 19538 32088 19628
rect 30497 19536 32088 19538
rect 18864 19472 19184 19488
rect 30497 19480 30502 19536
rect 30558 19480 32088 19536
rect 30497 19478 32088 19480
rect 30497 19475 30563 19478
rect 18864 19408 18872 19472
rect 18936 19408 18952 19472
rect 19016 19408 19032 19472
rect 19096 19408 19112 19472
rect 19176 19408 19184 19472
rect 18864 19392 19184 19408
rect 31648 19388 32088 19478
rect 3504 18928 3824 18944
rect 3504 18864 3512 18928
rect 3576 18864 3592 18928
rect 3656 18864 3672 18928
rect 3736 18864 3752 18928
rect 3816 18864 3824 18928
rect 3504 18848 3824 18864
rect 0 18722 440 18812
rect 5105 18722 5171 18725
rect 0 18720 5171 18722
rect 0 18664 5110 18720
rect 5166 18664 5171 18720
rect 0 18662 5171 18664
rect 0 18572 440 18662
rect 5105 18659 5171 18662
rect 18864 18384 19184 18400
rect 18864 18320 18872 18384
rect 18936 18320 18952 18384
rect 19016 18320 19032 18384
rect 19096 18320 19112 18384
rect 19176 18320 19184 18384
rect 18864 18304 19184 18320
rect 3504 17840 3824 17856
rect 3504 17776 3512 17840
rect 3576 17776 3592 17840
rect 3656 17776 3672 17840
rect 3736 17776 3752 17840
rect 3816 17776 3824 17840
rect 3504 17760 3824 17776
rect 4553 17362 4619 17365
rect 8417 17362 8483 17365
rect 4553 17360 8483 17362
rect 4553 17304 4558 17360
rect 4614 17304 8422 17360
rect 8478 17304 8483 17360
rect 26909 17362 26975 17365
rect 31648 17362 32088 17452
rect 26909 17360 32088 17362
rect 4553 17302 8483 17304
rect 4553 17299 4619 17302
rect 8417 17299 8483 17302
rect 18864 17296 19184 17312
rect 26909 17304 26914 17360
rect 26970 17304 32088 17360
rect 26909 17302 32088 17304
rect 26909 17299 26975 17302
rect 18864 17232 18872 17296
rect 18936 17232 18952 17296
rect 19016 17232 19032 17296
rect 19096 17232 19112 17296
rect 19176 17232 19184 17296
rect 18864 17216 19184 17232
rect 31648 17212 32088 17302
rect 3504 16752 3824 16768
rect 3504 16688 3512 16752
rect 3576 16688 3592 16752
rect 3656 16688 3672 16752
rect 3736 16688 3752 16752
rect 3816 16688 3824 16752
rect 3504 16672 3824 16688
rect 0 16546 440 16636
rect 1149 16546 1215 16549
rect 0 16544 1215 16546
rect 0 16488 1154 16544
rect 1210 16488 1215 16544
rect 0 16486 1215 16488
rect 0 16396 440 16486
rect 1149 16483 1215 16486
rect 18864 16208 19184 16224
rect 18864 16144 18872 16208
rect 18936 16144 18952 16208
rect 19016 16144 19032 16208
rect 19096 16144 19112 16208
rect 19176 16144 19184 16208
rect 18864 16128 19184 16144
rect 3504 15664 3824 15680
rect 3504 15600 3512 15664
rect 3576 15600 3592 15664
rect 3656 15600 3672 15664
rect 3736 15600 3752 15664
rect 3816 15600 3824 15664
rect 3504 15584 3824 15600
rect 30497 15458 30563 15461
rect 31648 15458 32088 15548
rect 30497 15456 32088 15458
rect 30497 15400 30502 15456
rect 30558 15400 32088 15456
rect 30497 15398 32088 15400
rect 30497 15395 30563 15398
rect 25529 15322 25595 15325
rect 27829 15322 27895 15325
rect 25529 15320 27895 15322
rect 25529 15264 25534 15320
rect 25590 15264 27834 15320
rect 27890 15264 27895 15320
rect 31648 15308 32088 15398
rect 25529 15262 27895 15264
rect 25529 15259 25595 15262
rect 27829 15259 27895 15262
rect 18864 15120 19184 15136
rect 18864 15056 18872 15120
rect 18936 15056 18952 15120
rect 19016 15056 19032 15120
rect 19096 15056 19112 15120
rect 19176 15056 19184 15120
rect 18864 15040 19184 15056
rect 0 14642 440 14732
rect 2621 14642 2687 14645
rect 0 14640 2687 14642
rect 0 14584 2626 14640
rect 2682 14584 2687 14640
rect 0 14582 2687 14584
rect 0 14492 440 14582
rect 2621 14579 2687 14582
rect 3504 14576 3824 14592
rect 3504 14512 3512 14576
rect 3576 14512 3592 14576
rect 3656 14512 3672 14576
rect 3736 14512 3752 14576
rect 3816 14512 3824 14576
rect 3504 14496 3824 14512
rect 8233 14234 8299 14237
rect 28565 14234 28631 14237
rect 8233 14232 28631 14234
rect 8233 14176 8238 14232
rect 8294 14176 28570 14232
rect 28626 14176 28631 14232
rect 8233 14174 28631 14176
rect 8233 14171 8299 14174
rect 28565 14171 28631 14174
rect 18864 14032 19184 14048
rect 18864 13968 18872 14032
rect 18936 13968 18952 14032
rect 19016 13968 19032 14032
rect 19096 13968 19112 14032
rect 19176 13968 19184 14032
rect 18864 13952 19184 13968
rect 17341 13826 17407 13829
rect 30497 13826 30563 13829
rect 17341 13824 30563 13826
rect 17341 13768 17346 13824
rect 17402 13768 30502 13824
rect 30558 13768 30563 13824
rect 17341 13766 30563 13768
rect 17341 13763 17407 13766
rect 30497 13763 30563 13766
rect 8049 13690 8115 13693
rect 26265 13690 26331 13693
rect 8049 13688 26331 13690
rect 8049 13632 8054 13688
rect 8110 13632 26270 13688
rect 26326 13632 26331 13688
rect 8049 13630 26331 13632
rect 8049 13627 8115 13630
rect 26265 13627 26331 13630
rect 3504 13488 3824 13504
rect 3504 13424 3512 13488
rect 3576 13424 3592 13488
rect 3656 13424 3672 13488
rect 3736 13424 3752 13488
rect 3816 13424 3824 13488
rect 3504 13408 3824 13424
rect 31648 13282 32088 13372
rect 31604 13132 32088 13282
rect 31604 13086 31698 13132
rect 18864 12944 19184 12960
rect 18864 12880 18872 12944
rect 18936 12880 18952 12944
rect 19016 12880 19032 12944
rect 19096 12880 19112 12944
rect 19176 12880 19184 12944
rect 18864 12864 19184 12880
rect 965 12738 1031 12741
rect 2069 12738 2135 12741
rect 9889 12738 9955 12741
rect 965 12736 9955 12738
rect 965 12680 970 12736
rect 1026 12680 2074 12736
rect 2130 12680 9894 12736
rect 9950 12680 9955 12736
rect 965 12678 9955 12680
rect 965 12675 1031 12678
rect 2069 12675 2135 12678
rect 9889 12675 9955 12678
rect 23045 12738 23111 12741
rect 31638 12738 31698 13086
rect 23045 12736 31698 12738
rect 23045 12680 23050 12736
rect 23106 12680 31698 12736
rect 23045 12678 31698 12680
rect 23045 12675 23111 12678
rect 0 12466 440 12556
rect 1241 12466 1307 12469
rect 0 12464 1307 12466
rect 0 12408 1246 12464
rect 1302 12408 1307 12464
rect 0 12406 1307 12408
rect 0 12316 440 12406
rect 1241 12403 1307 12406
rect 3504 12400 3824 12416
rect 3504 12336 3512 12400
rect 3576 12336 3592 12400
rect 3656 12336 3672 12400
rect 3736 12336 3752 12400
rect 3816 12336 3824 12400
rect 3504 12320 3824 12336
rect 9981 12058 10047 12061
rect 20561 12058 20627 12061
rect 9981 12056 20627 12058
rect 9981 12000 9986 12056
rect 10042 12000 20566 12056
rect 20622 12000 20627 12056
rect 9981 11998 20627 12000
rect 9981 11995 10047 11998
rect 20561 11995 20627 11998
rect 18864 11856 19184 11872
rect 18864 11792 18872 11856
rect 18936 11792 18952 11856
rect 19016 11792 19032 11856
rect 19096 11792 19112 11856
rect 19176 11792 19184 11856
rect 18864 11776 19184 11792
rect 1333 11650 1399 11653
rect 1333 11648 14230 11650
rect 1333 11592 1338 11648
rect 1394 11592 14230 11648
rect 1333 11590 14230 11592
rect 1333 11587 1399 11590
rect 14170 11514 14230 11590
rect 28841 11514 28907 11517
rect 14170 11512 29410 11514
rect 14170 11456 28846 11512
rect 28902 11456 29410 11512
rect 14170 11454 29410 11456
rect 28841 11451 28907 11454
rect 9705 11378 9771 11381
rect 20653 11378 20719 11381
rect 9705 11376 20719 11378
rect 3504 11312 3824 11328
rect 9705 11320 9710 11376
rect 9766 11320 20658 11376
rect 20714 11320 20719 11376
rect 9705 11318 20719 11320
rect 29350 11378 29410 11454
rect 31648 11378 32088 11468
rect 29350 11318 32088 11378
rect 9705 11315 9771 11318
rect 20653 11315 20719 11318
rect 3504 11248 3512 11312
rect 3576 11248 3592 11312
rect 3656 11248 3672 11312
rect 3736 11248 3752 11312
rect 3816 11248 3824 11312
rect 3504 11232 3824 11248
rect 31648 11228 32088 11318
rect 10165 10970 10231 10973
rect 23965 10970 24031 10973
rect 10165 10968 24031 10970
rect 10165 10912 10170 10968
rect 10226 10912 23970 10968
rect 24026 10912 24031 10968
rect 10165 10910 24031 10912
rect 10165 10907 10231 10910
rect 23965 10907 24031 10910
rect 18864 10768 19184 10784
rect 18864 10704 18872 10768
rect 18936 10704 18952 10768
rect 19016 10704 19032 10768
rect 19096 10704 19112 10768
rect 19176 10704 19184 10768
rect 18864 10688 19184 10704
rect 0 10562 440 10652
rect 1425 10562 1491 10565
rect 0 10560 1491 10562
rect 0 10504 1430 10560
rect 1486 10504 1491 10560
rect 0 10502 1491 10504
rect 0 10412 440 10502
rect 1425 10499 1491 10502
rect 7405 10562 7471 10565
rect 22953 10562 23019 10565
rect 7405 10560 23019 10562
rect 7405 10504 7410 10560
rect 7466 10504 22958 10560
rect 23014 10504 23019 10560
rect 7405 10502 23019 10504
rect 7405 10499 7471 10502
rect 22953 10499 23019 10502
rect 3504 10224 3824 10240
rect 3504 10160 3512 10224
rect 3576 10160 3592 10224
rect 3656 10160 3672 10224
rect 3736 10160 3752 10224
rect 3816 10160 3824 10224
rect 3504 10144 3824 10160
rect 10809 10154 10875 10157
rect 25713 10154 25779 10157
rect 10809 10152 25779 10154
rect 10809 10096 10814 10152
rect 10870 10096 25718 10152
rect 25774 10096 25779 10152
rect 10809 10094 25779 10096
rect 10809 10091 10875 10094
rect 25713 10091 25779 10094
rect 12741 9882 12807 9885
rect 20377 9882 20443 9885
rect 12741 9880 20443 9882
rect 12741 9824 12746 9880
rect 12802 9824 20382 9880
rect 20438 9824 20443 9880
rect 12741 9822 20443 9824
rect 12741 9819 12807 9822
rect 20377 9819 20443 9822
rect 20653 9882 20719 9885
rect 24057 9882 24123 9885
rect 20653 9880 24123 9882
rect 20653 9824 20658 9880
rect 20714 9824 24062 9880
rect 24118 9824 24123 9880
rect 20653 9822 24123 9824
rect 20653 9819 20719 9822
rect 24057 9819 24123 9822
rect 18864 9680 19184 9696
rect 18864 9616 18872 9680
rect 18936 9616 18952 9680
rect 19016 9616 19032 9680
rect 19096 9616 19112 9680
rect 19176 9616 19184 9680
rect 18864 9600 19184 9616
rect 8601 9474 8667 9477
rect 18261 9474 18327 9477
rect 8601 9472 18327 9474
rect 8601 9416 8606 9472
rect 8662 9416 18266 9472
rect 18322 9416 18327 9472
rect 8601 9414 18327 9416
rect 8601 9411 8667 9414
rect 18261 9411 18327 9414
rect 18445 9474 18511 9477
rect 24333 9474 24399 9477
rect 18445 9472 24399 9474
rect 18445 9416 18450 9472
rect 18506 9416 24338 9472
rect 24394 9416 24399 9472
rect 18445 9414 24399 9416
rect 18445 9411 18511 9414
rect 24333 9411 24399 9414
rect 12005 9338 12071 9341
rect 23137 9338 23203 9341
rect 12005 9336 23203 9338
rect 12005 9280 12010 9336
rect 12066 9280 23142 9336
rect 23198 9280 23203 9336
rect 12005 9278 23203 9280
rect 12005 9275 12071 9278
rect 23137 9275 23203 9278
rect 6025 9202 6091 9205
rect 20653 9202 20719 9205
rect 6025 9200 20719 9202
rect 3504 9136 3824 9152
rect 6025 9144 6030 9200
rect 6086 9144 20658 9200
rect 20714 9144 20719 9200
rect 6025 9142 20719 9144
rect 6025 9139 6091 9142
rect 20653 9139 20719 9142
rect 29945 9202 30011 9205
rect 31648 9202 32088 9292
rect 29945 9200 32088 9202
rect 29945 9144 29950 9200
rect 30006 9144 32088 9200
rect 29945 9142 32088 9144
rect 29945 9139 30011 9142
rect 3504 9072 3512 9136
rect 3576 9072 3592 9136
rect 3656 9072 3672 9136
rect 3736 9072 3752 9136
rect 3816 9072 3824 9136
rect 3504 9056 3824 9072
rect 31648 9052 32088 9142
rect 18864 8592 19184 8608
rect 18864 8528 18872 8592
rect 18936 8528 18952 8592
rect 19016 8528 19032 8592
rect 19096 8528 19112 8592
rect 19176 8528 19184 8592
rect 18864 8512 19184 8528
rect 0 8386 440 8476
rect 7681 8386 7747 8389
rect 0 8384 7747 8386
rect 0 8328 7686 8384
rect 7742 8328 7747 8384
rect 0 8326 7747 8328
rect 0 8236 440 8326
rect 7681 8323 7747 8326
rect 17801 8250 17867 8253
rect 25897 8250 25963 8253
rect 17801 8248 25963 8250
rect 17801 8192 17806 8248
rect 17862 8192 25902 8248
rect 25958 8192 25963 8248
rect 17801 8190 25963 8192
rect 17801 8187 17867 8190
rect 25897 8187 25963 8190
rect 5841 8114 5907 8117
rect 23781 8114 23847 8117
rect 5841 8112 23847 8114
rect 3504 8048 3824 8064
rect 5841 8056 5846 8112
rect 5902 8056 23786 8112
rect 23842 8056 23847 8112
rect 5841 8054 23847 8056
rect 5841 8051 5907 8054
rect 23781 8051 23847 8054
rect 3504 7984 3512 8048
rect 3576 7984 3592 8048
rect 3656 7984 3672 8048
rect 3736 7984 3752 8048
rect 3816 7984 3824 8048
rect 3504 7968 3824 7984
rect 5933 7978 5999 7981
rect 23873 7978 23939 7981
rect 5933 7976 23939 7978
rect 5933 7920 5938 7976
rect 5994 7920 23878 7976
rect 23934 7920 23939 7976
rect 5933 7918 23939 7920
rect 5933 7915 5999 7918
rect 23873 7915 23939 7918
rect 18864 7504 19184 7520
rect 18864 7440 18872 7504
rect 18936 7440 18952 7504
rect 19016 7440 19032 7504
rect 19096 7440 19112 7504
rect 19176 7440 19184 7504
rect 18864 7424 19184 7440
rect 8877 7298 8943 7301
rect 20561 7298 20627 7301
rect 8877 7296 20627 7298
rect 8877 7240 8882 7296
rect 8938 7240 20566 7296
rect 20622 7240 20627 7296
rect 8877 7238 20627 7240
rect 8877 7235 8943 7238
rect 20561 7235 20627 7238
rect 30497 7298 30563 7301
rect 31648 7298 32088 7388
rect 30497 7296 32088 7298
rect 30497 7240 30502 7296
rect 30558 7240 32088 7296
rect 30497 7238 32088 7240
rect 30497 7235 30563 7238
rect 31648 7148 32088 7238
rect 3504 6960 3824 6976
rect 3504 6896 3512 6960
rect 3576 6896 3592 6960
rect 3656 6896 3672 6960
rect 3736 6896 3752 6960
rect 3816 6896 3824 6960
rect 3504 6880 3824 6896
rect 4277 6618 4343 6621
rect 4829 6618 4895 6621
rect 4277 6616 4895 6618
rect 0 6482 440 6572
rect 4277 6560 4282 6616
rect 4338 6560 4834 6616
rect 4890 6560 4895 6616
rect 4277 6558 4895 6560
rect 4277 6555 4343 6558
rect 4829 6555 4895 6558
rect 873 6482 939 6485
rect 0 6480 939 6482
rect 0 6424 878 6480
rect 934 6424 939 6480
rect 0 6422 939 6424
rect 0 6332 440 6422
rect 873 6419 939 6422
rect 18864 6416 19184 6432
rect 18864 6352 18872 6416
rect 18936 6352 18952 6416
rect 19016 6352 19032 6416
rect 19096 6352 19112 6416
rect 19176 6352 19184 6416
rect 18864 6336 19184 6352
rect 3504 5872 3824 5888
rect 3504 5808 3512 5872
rect 3576 5808 3592 5872
rect 3656 5808 3672 5872
rect 3736 5808 3752 5872
rect 3816 5808 3824 5872
rect 3504 5792 3824 5808
rect 16329 5666 16395 5669
rect 26541 5666 26607 5669
rect 16329 5664 26607 5666
rect 16329 5608 16334 5664
rect 16390 5608 26546 5664
rect 26602 5608 26607 5664
rect 16329 5606 26607 5608
rect 16329 5603 16395 5606
rect 26541 5603 26607 5606
rect 19365 5394 19431 5397
rect 28749 5394 28815 5397
rect 19365 5392 28815 5394
rect 18864 5328 19184 5344
rect 19365 5336 19370 5392
rect 19426 5336 28754 5392
rect 28810 5336 28815 5392
rect 19365 5334 28815 5336
rect 19365 5331 19431 5334
rect 28749 5331 28815 5334
rect 18864 5264 18872 5328
rect 18936 5264 18952 5328
rect 19016 5264 19032 5328
rect 19096 5264 19112 5328
rect 19176 5264 19184 5328
rect 18864 5248 19184 5264
rect 22217 5258 22283 5261
rect 30497 5258 30563 5261
rect 22217 5256 30563 5258
rect 22217 5200 22222 5256
rect 22278 5200 30502 5256
rect 30558 5200 30563 5256
rect 22217 5198 30563 5200
rect 22217 5195 22283 5198
rect 30497 5195 30563 5198
rect 31648 5122 32088 5212
rect 31604 4972 32088 5122
rect 31604 4926 31698 4972
rect 3504 4784 3824 4800
rect 3504 4720 3512 4784
rect 3576 4720 3592 4784
rect 3656 4720 3672 4784
rect 3736 4720 3752 4784
rect 3816 4720 3824 4784
rect 3504 4704 3824 4720
rect 18629 4578 18695 4581
rect 19273 4578 19339 4581
rect 18629 4576 19339 4578
rect 18629 4520 18634 4576
rect 18690 4520 19278 4576
rect 19334 4520 19339 4576
rect 18629 4518 19339 4520
rect 18629 4515 18695 4518
rect 19273 4515 19339 4518
rect 21481 4578 21547 4581
rect 31638 4578 31698 4926
rect 21481 4576 31698 4578
rect 21481 4520 21486 4576
rect 21542 4520 31698 4576
rect 21481 4518 31698 4520
rect 21481 4515 21547 4518
rect 0 4306 440 4396
rect 1241 4306 1307 4309
rect 0 4304 1307 4306
rect 0 4248 1246 4304
rect 1302 4248 1307 4304
rect 0 4246 1307 4248
rect 0 4156 440 4246
rect 1241 4243 1307 4246
rect 18864 4240 19184 4256
rect 18864 4176 18872 4240
rect 18936 4176 18952 4240
rect 19016 4176 19032 4240
rect 19096 4176 19112 4240
rect 19176 4176 19184 4240
rect 18864 4160 19184 4176
rect 11729 3762 11795 3765
rect 19641 3762 19707 3765
rect 20469 3762 20535 3765
rect 11729 3760 20535 3762
rect 3504 3696 3824 3712
rect 11729 3704 11734 3760
rect 11790 3704 19646 3760
rect 19702 3704 20474 3760
rect 20530 3704 20535 3760
rect 11729 3702 20535 3704
rect 11729 3699 11795 3702
rect 19641 3699 19707 3702
rect 20469 3699 20535 3702
rect 3504 3632 3512 3696
rect 3576 3632 3592 3696
rect 3656 3632 3672 3696
rect 3736 3632 3752 3696
rect 3816 3632 3824 3696
rect 3504 3616 3824 3632
rect 12557 3490 12623 3493
rect 25437 3490 25503 3493
rect 12557 3488 25503 3490
rect 12557 3432 12562 3488
rect 12618 3432 25442 3488
rect 25498 3432 25503 3488
rect 12557 3430 25503 3432
rect 12557 3427 12623 3430
rect 25437 3427 25503 3430
rect 10993 3354 11059 3357
rect 23413 3354 23479 3357
rect 23781 3354 23847 3357
rect 10993 3352 23847 3354
rect 10993 3296 10998 3352
rect 11054 3296 23418 3352
rect 23474 3296 23786 3352
rect 23842 3296 23847 3352
rect 10993 3294 23847 3296
rect 10993 3291 11059 3294
rect 23413 3291 23479 3294
rect 23781 3291 23847 3294
rect 30497 3218 30563 3221
rect 31648 3218 32088 3308
rect 30497 3216 32088 3218
rect 18864 3152 19184 3168
rect 30497 3160 30502 3216
rect 30558 3160 32088 3216
rect 30497 3158 32088 3160
rect 30497 3155 30563 3158
rect 18864 3088 18872 3152
rect 18936 3088 18952 3152
rect 19016 3088 19032 3152
rect 19096 3088 19112 3152
rect 19176 3088 19184 3152
rect 18864 3072 19184 3088
rect 31648 3068 32088 3158
rect 3504 2608 3824 2624
rect 3504 2544 3512 2608
rect 3576 2544 3592 2608
rect 3656 2544 3672 2608
rect 3736 2544 3752 2608
rect 3816 2544 3824 2608
rect 3504 2528 3824 2544
rect 0 2402 440 2492
rect 1149 2402 1215 2405
rect 0 2400 1215 2402
rect 0 2344 1154 2400
rect 1210 2344 1215 2400
rect 0 2342 1215 2344
rect 0 2252 440 2342
rect 1149 2339 1215 2342
rect 18864 2064 19184 2080
rect 18864 2000 18872 2064
rect 18936 2000 18952 2064
rect 19016 2000 19032 2064
rect 19096 2000 19112 2064
rect 19176 2000 19184 2064
rect 18864 1984 19184 2000
rect 3504 1520 3824 1536
rect 3504 1456 3512 1520
rect 3576 1456 3592 1520
rect 3656 1456 3672 1520
rect 3736 1456 3752 1520
rect 3816 1456 3824 1520
rect 3504 1440 3824 1456
rect 31648 1044 32088 1132
rect 31630 1042 31636 1044
rect 18864 976 19184 992
rect 31508 982 31636 1042
rect 31630 980 31636 982
rect 31700 980 32088 1044
rect 18864 912 18872 976
rect 18936 912 18952 976
rect 19016 912 19032 976
rect 19096 912 19112 976
rect 19176 912 19184 976
rect 18864 896 19184 912
rect 31648 892 32088 980
rect 5933 770 5999 773
rect 17709 770 17775 773
rect 5933 768 17775 770
rect 5933 712 5938 768
rect 5994 712 17714 768
rect 17770 712 17775 768
rect 5933 710 17775 712
rect 5933 707 5999 710
rect 17709 707 17775 710
rect 19549 770 19615 773
rect 28013 770 28079 773
rect 19549 768 28079 770
rect 19549 712 19554 768
rect 19610 712 28018 768
rect 28074 712 28079 768
rect 19549 710 28079 712
rect 19549 707 19615 710
rect 28013 707 28079 710
rect 31630 708 31636 772
rect 31700 708 31706 772
rect 413 634 479 637
rect 20929 634 20995 637
rect 413 632 20995 634
rect 413 576 418 632
rect 474 576 20934 632
rect 20990 576 20995 632
rect 413 574 20995 576
rect 413 571 479 574
rect 20929 571 20995 574
rect 20561 498 20627 501
rect 12744 496 20627 498
rect 3504 432 3824 448
rect 12744 445 20566 496
rect 3504 368 3512 432
rect 3576 368 3592 432
rect 3656 368 3672 432
rect 3736 368 3752 432
rect 3816 368 3824 432
rect 12741 440 20566 445
rect 20622 440 20627 496
rect 12741 384 12746 440
rect 12802 438 20627 440
rect 12802 384 12807 438
rect 20561 435 20627 438
rect 20745 498 20811 501
rect 31638 498 31698 708
rect 20745 496 31698 498
rect 20745 440 20750 496
rect 20806 440 31698 496
rect 20745 438 31698 440
rect 20745 435 20811 438
rect 12741 379 12807 384
rect 3504 352 3824 368
<< via3 >>
rect 18872 31436 18936 31440
rect 18872 31380 18876 31436
rect 18876 31380 18932 31436
rect 18932 31380 18936 31436
rect 18872 31376 18936 31380
rect 18952 31436 19016 31440
rect 18952 31380 18956 31436
rect 18956 31380 19012 31436
rect 19012 31380 19016 31436
rect 18952 31376 19016 31380
rect 19032 31436 19096 31440
rect 19032 31380 19036 31436
rect 19036 31380 19092 31436
rect 19092 31380 19096 31436
rect 19032 31376 19096 31380
rect 19112 31436 19176 31440
rect 19112 31380 19116 31436
rect 19116 31380 19172 31436
rect 19172 31380 19176 31436
rect 19112 31376 19176 31380
rect 3512 30892 3576 30896
rect 3512 30836 3516 30892
rect 3516 30836 3572 30892
rect 3572 30836 3576 30892
rect 3512 30832 3576 30836
rect 3592 30892 3656 30896
rect 3592 30836 3596 30892
rect 3596 30836 3652 30892
rect 3652 30836 3656 30892
rect 3592 30832 3656 30836
rect 3672 30892 3736 30896
rect 3672 30836 3676 30892
rect 3676 30836 3732 30892
rect 3732 30836 3736 30892
rect 3672 30832 3736 30836
rect 3752 30892 3816 30896
rect 3752 30836 3756 30892
rect 3756 30836 3812 30892
rect 3812 30836 3816 30892
rect 3752 30832 3816 30836
rect 18872 30348 18936 30352
rect 18872 30292 18876 30348
rect 18876 30292 18932 30348
rect 18932 30292 18936 30348
rect 18872 30288 18936 30292
rect 18952 30348 19016 30352
rect 18952 30292 18956 30348
rect 18956 30292 19012 30348
rect 19012 30292 19016 30348
rect 18952 30288 19016 30292
rect 19032 30348 19096 30352
rect 19032 30292 19036 30348
rect 19036 30292 19092 30348
rect 19092 30292 19096 30348
rect 19032 30288 19096 30292
rect 19112 30348 19176 30352
rect 19112 30292 19116 30348
rect 19116 30292 19172 30348
rect 19172 30292 19176 30348
rect 19112 30288 19176 30292
rect 3512 29804 3576 29808
rect 3512 29748 3516 29804
rect 3516 29748 3572 29804
rect 3572 29748 3576 29804
rect 3512 29744 3576 29748
rect 3592 29804 3656 29808
rect 3592 29748 3596 29804
rect 3596 29748 3652 29804
rect 3652 29748 3656 29804
rect 3592 29744 3656 29748
rect 3672 29804 3736 29808
rect 3672 29748 3676 29804
rect 3676 29748 3732 29804
rect 3732 29748 3736 29804
rect 3672 29744 3736 29748
rect 3752 29804 3816 29808
rect 3752 29748 3756 29804
rect 3756 29748 3812 29804
rect 3812 29748 3816 29804
rect 3752 29744 3816 29748
rect 18872 29260 18936 29264
rect 18872 29204 18876 29260
rect 18876 29204 18932 29260
rect 18932 29204 18936 29260
rect 18872 29200 18936 29204
rect 18952 29260 19016 29264
rect 18952 29204 18956 29260
rect 18956 29204 19012 29260
rect 19012 29204 19016 29260
rect 18952 29200 19016 29204
rect 19032 29260 19096 29264
rect 19032 29204 19036 29260
rect 19036 29204 19092 29260
rect 19092 29204 19096 29260
rect 19032 29200 19096 29204
rect 19112 29260 19176 29264
rect 19112 29204 19116 29260
rect 19116 29204 19172 29260
rect 19172 29204 19176 29260
rect 19112 29200 19176 29204
rect 3512 28716 3576 28720
rect 3512 28660 3516 28716
rect 3516 28660 3572 28716
rect 3572 28660 3576 28716
rect 3512 28656 3576 28660
rect 3592 28716 3656 28720
rect 3592 28660 3596 28716
rect 3596 28660 3652 28716
rect 3652 28660 3656 28716
rect 3592 28656 3656 28660
rect 3672 28716 3736 28720
rect 3672 28660 3676 28716
rect 3676 28660 3732 28716
rect 3732 28660 3736 28716
rect 3672 28656 3736 28660
rect 3752 28716 3816 28720
rect 3752 28660 3756 28716
rect 3756 28660 3812 28716
rect 3812 28660 3816 28716
rect 3752 28656 3816 28660
rect 18872 28172 18936 28176
rect 18872 28116 18876 28172
rect 18876 28116 18932 28172
rect 18932 28116 18936 28172
rect 18872 28112 18936 28116
rect 18952 28172 19016 28176
rect 18952 28116 18956 28172
rect 18956 28116 19012 28172
rect 19012 28116 19016 28172
rect 18952 28112 19016 28116
rect 19032 28172 19096 28176
rect 19032 28116 19036 28172
rect 19036 28116 19092 28172
rect 19092 28116 19096 28172
rect 19032 28112 19096 28116
rect 19112 28172 19176 28176
rect 19112 28116 19116 28172
rect 19116 28116 19172 28172
rect 19172 28116 19176 28172
rect 19112 28112 19176 28116
rect 3512 27628 3576 27632
rect 3512 27572 3516 27628
rect 3516 27572 3572 27628
rect 3572 27572 3576 27628
rect 3512 27568 3576 27572
rect 3592 27628 3656 27632
rect 3592 27572 3596 27628
rect 3596 27572 3652 27628
rect 3652 27572 3656 27628
rect 3592 27568 3656 27572
rect 3672 27628 3736 27632
rect 3672 27572 3676 27628
rect 3676 27572 3732 27628
rect 3732 27572 3736 27628
rect 3672 27568 3736 27572
rect 3752 27628 3816 27632
rect 3752 27572 3756 27628
rect 3756 27572 3812 27628
rect 3812 27572 3816 27628
rect 3752 27568 3816 27572
rect 18872 27084 18936 27088
rect 18872 27028 18876 27084
rect 18876 27028 18932 27084
rect 18932 27028 18936 27084
rect 18872 27024 18936 27028
rect 18952 27084 19016 27088
rect 18952 27028 18956 27084
rect 18956 27028 19012 27084
rect 19012 27028 19016 27084
rect 18952 27024 19016 27028
rect 19032 27084 19096 27088
rect 19032 27028 19036 27084
rect 19036 27028 19092 27084
rect 19092 27028 19096 27084
rect 19032 27024 19096 27028
rect 19112 27084 19176 27088
rect 19112 27028 19116 27084
rect 19116 27028 19172 27084
rect 19172 27028 19176 27084
rect 19112 27024 19176 27028
rect 3512 26540 3576 26544
rect 3512 26484 3516 26540
rect 3516 26484 3572 26540
rect 3572 26484 3576 26540
rect 3512 26480 3576 26484
rect 3592 26540 3656 26544
rect 3592 26484 3596 26540
rect 3596 26484 3652 26540
rect 3652 26484 3656 26540
rect 3592 26480 3656 26484
rect 3672 26540 3736 26544
rect 3672 26484 3676 26540
rect 3676 26484 3732 26540
rect 3732 26484 3736 26540
rect 3672 26480 3736 26484
rect 3752 26540 3816 26544
rect 3752 26484 3756 26540
rect 3756 26484 3812 26540
rect 3812 26484 3816 26540
rect 3752 26480 3816 26484
rect 18872 25996 18936 26000
rect 18872 25940 18876 25996
rect 18876 25940 18932 25996
rect 18932 25940 18936 25996
rect 18872 25936 18936 25940
rect 18952 25996 19016 26000
rect 18952 25940 18956 25996
rect 18956 25940 19012 25996
rect 19012 25940 19016 25996
rect 18952 25936 19016 25940
rect 19032 25996 19096 26000
rect 19032 25940 19036 25996
rect 19036 25940 19092 25996
rect 19092 25940 19096 25996
rect 19032 25936 19096 25940
rect 19112 25996 19176 26000
rect 19112 25940 19116 25996
rect 19116 25940 19172 25996
rect 19172 25940 19176 25996
rect 19112 25936 19176 25940
rect 3512 25452 3576 25456
rect 3512 25396 3516 25452
rect 3516 25396 3572 25452
rect 3572 25396 3576 25452
rect 3512 25392 3576 25396
rect 3592 25452 3656 25456
rect 3592 25396 3596 25452
rect 3596 25396 3652 25452
rect 3652 25396 3656 25452
rect 3592 25392 3656 25396
rect 3672 25452 3736 25456
rect 3672 25396 3676 25452
rect 3676 25396 3732 25452
rect 3732 25396 3736 25452
rect 3672 25392 3736 25396
rect 3752 25452 3816 25456
rect 3752 25396 3756 25452
rect 3756 25396 3812 25452
rect 3812 25396 3816 25452
rect 3752 25392 3816 25396
rect 18872 24908 18936 24912
rect 18872 24852 18876 24908
rect 18876 24852 18932 24908
rect 18932 24852 18936 24908
rect 18872 24848 18936 24852
rect 18952 24908 19016 24912
rect 18952 24852 18956 24908
rect 18956 24852 19012 24908
rect 19012 24852 19016 24908
rect 18952 24848 19016 24852
rect 19032 24908 19096 24912
rect 19032 24852 19036 24908
rect 19036 24852 19092 24908
rect 19092 24852 19096 24908
rect 19032 24848 19096 24852
rect 19112 24908 19176 24912
rect 19112 24852 19116 24908
rect 19116 24852 19172 24908
rect 19172 24852 19176 24908
rect 19112 24848 19176 24852
rect 3512 24364 3576 24368
rect 3512 24308 3516 24364
rect 3516 24308 3572 24364
rect 3572 24308 3576 24364
rect 3512 24304 3576 24308
rect 3592 24364 3656 24368
rect 3592 24308 3596 24364
rect 3596 24308 3652 24364
rect 3652 24308 3656 24364
rect 3592 24304 3656 24308
rect 3672 24364 3736 24368
rect 3672 24308 3676 24364
rect 3676 24308 3732 24364
rect 3732 24308 3736 24364
rect 3672 24304 3736 24308
rect 3752 24364 3816 24368
rect 3752 24308 3756 24364
rect 3756 24308 3812 24364
rect 3812 24308 3816 24364
rect 3752 24304 3816 24308
rect 18872 23820 18936 23824
rect 18872 23764 18876 23820
rect 18876 23764 18932 23820
rect 18932 23764 18936 23820
rect 18872 23760 18936 23764
rect 18952 23820 19016 23824
rect 18952 23764 18956 23820
rect 18956 23764 19012 23820
rect 19012 23764 19016 23820
rect 18952 23760 19016 23764
rect 19032 23820 19096 23824
rect 19032 23764 19036 23820
rect 19036 23764 19092 23820
rect 19092 23764 19096 23820
rect 19032 23760 19096 23764
rect 19112 23820 19176 23824
rect 19112 23764 19116 23820
rect 19116 23764 19172 23820
rect 19172 23764 19176 23820
rect 19112 23760 19176 23764
rect 3512 23276 3576 23280
rect 3512 23220 3516 23276
rect 3516 23220 3572 23276
rect 3572 23220 3576 23276
rect 3512 23216 3576 23220
rect 3592 23276 3656 23280
rect 3592 23220 3596 23276
rect 3596 23220 3652 23276
rect 3652 23220 3656 23276
rect 3592 23216 3656 23220
rect 3672 23276 3736 23280
rect 3672 23220 3676 23276
rect 3676 23220 3732 23276
rect 3732 23220 3736 23276
rect 3672 23216 3736 23220
rect 3752 23276 3816 23280
rect 3752 23220 3756 23276
rect 3756 23220 3812 23276
rect 3812 23220 3816 23276
rect 3752 23216 3816 23220
rect 18872 22732 18936 22736
rect 18872 22676 18876 22732
rect 18876 22676 18932 22732
rect 18932 22676 18936 22732
rect 18872 22672 18936 22676
rect 18952 22732 19016 22736
rect 18952 22676 18956 22732
rect 18956 22676 19012 22732
rect 19012 22676 19016 22732
rect 18952 22672 19016 22676
rect 19032 22732 19096 22736
rect 19032 22676 19036 22732
rect 19036 22676 19092 22732
rect 19092 22676 19096 22732
rect 19032 22672 19096 22676
rect 19112 22732 19176 22736
rect 19112 22676 19116 22732
rect 19116 22676 19172 22732
rect 19172 22676 19176 22732
rect 19112 22672 19176 22676
rect 3512 22188 3576 22192
rect 3512 22132 3516 22188
rect 3516 22132 3572 22188
rect 3572 22132 3576 22188
rect 3512 22128 3576 22132
rect 3592 22188 3656 22192
rect 3592 22132 3596 22188
rect 3596 22132 3652 22188
rect 3652 22132 3656 22188
rect 3592 22128 3656 22132
rect 3672 22188 3736 22192
rect 3672 22132 3676 22188
rect 3676 22132 3732 22188
rect 3732 22132 3736 22188
rect 3672 22128 3736 22132
rect 3752 22188 3816 22192
rect 3752 22132 3756 22188
rect 3756 22132 3812 22188
rect 3812 22132 3816 22188
rect 3752 22128 3816 22132
rect 18872 21644 18936 21648
rect 18872 21588 18876 21644
rect 18876 21588 18932 21644
rect 18932 21588 18936 21644
rect 18872 21584 18936 21588
rect 18952 21644 19016 21648
rect 18952 21588 18956 21644
rect 18956 21588 19012 21644
rect 19012 21588 19016 21644
rect 18952 21584 19016 21588
rect 19032 21644 19096 21648
rect 19032 21588 19036 21644
rect 19036 21588 19092 21644
rect 19092 21588 19096 21644
rect 19032 21584 19096 21588
rect 19112 21644 19176 21648
rect 19112 21588 19116 21644
rect 19116 21588 19172 21644
rect 19172 21588 19176 21644
rect 19112 21584 19176 21588
rect 3512 21100 3576 21104
rect 3512 21044 3516 21100
rect 3516 21044 3572 21100
rect 3572 21044 3576 21100
rect 3512 21040 3576 21044
rect 3592 21100 3656 21104
rect 3592 21044 3596 21100
rect 3596 21044 3652 21100
rect 3652 21044 3656 21100
rect 3592 21040 3656 21044
rect 3672 21100 3736 21104
rect 3672 21044 3676 21100
rect 3676 21044 3732 21100
rect 3732 21044 3736 21100
rect 3672 21040 3736 21044
rect 3752 21100 3816 21104
rect 3752 21044 3756 21100
rect 3756 21044 3812 21100
rect 3812 21044 3816 21100
rect 3752 21040 3816 21044
rect 18872 20556 18936 20560
rect 18872 20500 18876 20556
rect 18876 20500 18932 20556
rect 18932 20500 18936 20556
rect 18872 20496 18936 20500
rect 18952 20556 19016 20560
rect 18952 20500 18956 20556
rect 18956 20500 19012 20556
rect 19012 20500 19016 20556
rect 18952 20496 19016 20500
rect 19032 20556 19096 20560
rect 19032 20500 19036 20556
rect 19036 20500 19092 20556
rect 19092 20500 19096 20556
rect 19032 20496 19096 20500
rect 19112 20556 19176 20560
rect 19112 20500 19116 20556
rect 19116 20500 19172 20556
rect 19172 20500 19176 20556
rect 19112 20496 19176 20500
rect 3512 20012 3576 20016
rect 3512 19956 3516 20012
rect 3516 19956 3572 20012
rect 3572 19956 3576 20012
rect 3512 19952 3576 19956
rect 3592 20012 3656 20016
rect 3592 19956 3596 20012
rect 3596 19956 3652 20012
rect 3652 19956 3656 20012
rect 3592 19952 3656 19956
rect 3672 20012 3736 20016
rect 3672 19956 3676 20012
rect 3676 19956 3732 20012
rect 3732 19956 3736 20012
rect 3672 19952 3736 19956
rect 3752 20012 3816 20016
rect 3752 19956 3756 20012
rect 3756 19956 3812 20012
rect 3812 19956 3816 20012
rect 3752 19952 3816 19956
rect 18872 19468 18936 19472
rect 18872 19412 18876 19468
rect 18876 19412 18932 19468
rect 18932 19412 18936 19468
rect 18872 19408 18936 19412
rect 18952 19468 19016 19472
rect 18952 19412 18956 19468
rect 18956 19412 19012 19468
rect 19012 19412 19016 19468
rect 18952 19408 19016 19412
rect 19032 19468 19096 19472
rect 19032 19412 19036 19468
rect 19036 19412 19092 19468
rect 19092 19412 19096 19468
rect 19032 19408 19096 19412
rect 19112 19468 19176 19472
rect 19112 19412 19116 19468
rect 19116 19412 19172 19468
rect 19172 19412 19176 19468
rect 19112 19408 19176 19412
rect 3512 18924 3576 18928
rect 3512 18868 3516 18924
rect 3516 18868 3572 18924
rect 3572 18868 3576 18924
rect 3512 18864 3576 18868
rect 3592 18924 3656 18928
rect 3592 18868 3596 18924
rect 3596 18868 3652 18924
rect 3652 18868 3656 18924
rect 3592 18864 3656 18868
rect 3672 18924 3736 18928
rect 3672 18868 3676 18924
rect 3676 18868 3732 18924
rect 3732 18868 3736 18924
rect 3672 18864 3736 18868
rect 3752 18924 3816 18928
rect 3752 18868 3756 18924
rect 3756 18868 3812 18924
rect 3812 18868 3816 18924
rect 3752 18864 3816 18868
rect 18872 18380 18936 18384
rect 18872 18324 18876 18380
rect 18876 18324 18932 18380
rect 18932 18324 18936 18380
rect 18872 18320 18936 18324
rect 18952 18380 19016 18384
rect 18952 18324 18956 18380
rect 18956 18324 19012 18380
rect 19012 18324 19016 18380
rect 18952 18320 19016 18324
rect 19032 18380 19096 18384
rect 19032 18324 19036 18380
rect 19036 18324 19092 18380
rect 19092 18324 19096 18380
rect 19032 18320 19096 18324
rect 19112 18380 19176 18384
rect 19112 18324 19116 18380
rect 19116 18324 19172 18380
rect 19172 18324 19176 18380
rect 19112 18320 19176 18324
rect 3512 17836 3576 17840
rect 3512 17780 3516 17836
rect 3516 17780 3572 17836
rect 3572 17780 3576 17836
rect 3512 17776 3576 17780
rect 3592 17836 3656 17840
rect 3592 17780 3596 17836
rect 3596 17780 3652 17836
rect 3652 17780 3656 17836
rect 3592 17776 3656 17780
rect 3672 17836 3736 17840
rect 3672 17780 3676 17836
rect 3676 17780 3732 17836
rect 3732 17780 3736 17836
rect 3672 17776 3736 17780
rect 3752 17836 3816 17840
rect 3752 17780 3756 17836
rect 3756 17780 3812 17836
rect 3812 17780 3816 17836
rect 3752 17776 3816 17780
rect 18872 17292 18936 17296
rect 18872 17236 18876 17292
rect 18876 17236 18932 17292
rect 18932 17236 18936 17292
rect 18872 17232 18936 17236
rect 18952 17292 19016 17296
rect 18952 17236 18956 17292
rect 18956 17236 19012 17292
rect 19012 17236 19016 17292
rect 18952 17232 19016 17236
rect 19032 17292 19096 17296
rect 19032 17236 19036 17292
rect 19036 17236 19092 17292
rect 19092 17236 19096 17292
rect 19032 17232 19096 17236
rect 19112 17292 19176 17296
rect 19112 17236 19116 17292
rect 19116 17236 19172 17292
rect 19172 17236 19176 17292
rect 19112 17232 19176 17236
rect 3512 16748 3576 16752
rect 3512 16692 3516 16748
rect 3516 16692 3572 16748
rect 3572 16692 3576 16748
rect 3512 16688 3576 16692
rect 3592 16748 3656 16752
rect 3592 16692 3596 16748
rect 3596 16692 3652 16748
rect 3652 16692 3656 16748
rect 3592 16688 3656 16692
rect 3672 16748 3736 16752
rect 3672 16692 3676 16748
rect 3676 16692 3732 16748
rect 3732 16692 3736 16748
rect 3672 16688 3736 16692
rect 3752 16748 3816 16752
rect 3752 16692 3756 16748
rect 3756 16692 3812 16748
rect 3812 16692 3816 16748
rect 3752 16688 3816 16692
rect 18872 16204 18936 16208
rect 18872 16148 18876 16204
rect 18876 16148 18932 16204
rect 18932 16148 18936 16204
rect 18872 16144 18936 16148
rect 18952 16204 19016 16208
rect 18952 16148 18956 16204
rect 18956 16148 19012 16204
rect 19012 16148 19016 16204
rect 18952 16144 19016 16148
rect 19032 16204 19096 16208
rect 19032 16148 19036 16204
rect 19036 16148 19092 16204
rect 19092 16148 19096 16204
rect 19032 16144 19096 16148
rect 19112 16204 19176 16208
rect 19112 16148 19116 16204
rect 19116 16148 19172 16204
rect 19172 16148 19176 16204
rect 19112 16144 19176 16148
rect 3512 15660 3576 15664
rect 3512 15604 3516 15660
rect 3516 15604 3572 15660
rect 3572 15604 3576 15660
rect 3512 15600 3576 15604
rect 3592 15660 3656 15664
rect 3592 15604 3596 15660
rect 3596 15604 3652 15660
rect 3652 15604 3656 15660
rect 3592 15600 3656 15604
rect 3672 15660 3736 15664
rect 3672 15604 3676 15660
rect 3676 15604 3732 15660
rect 3732 15604 3736 15660
rect 3672 15600 3736 15604
rect 3752 15660 3816 15664
rect 3752 15604 3756 15660
rect 3756 15604 3812 15660
rect 3812 15604 3816 15660
rect 3752 15600 3816 15604
rect 18872 15116 18936 15120
rect 18872 15060 18876 15116
rect 18876 15060 18932 15116
rect 18932 15060 18936 15116
rect 18872 15056 18936 15060
rect 18952 15116 19016 15120
rect 18952 15060 18956 15116
rect 18956 15060 19012 15116
rect 19012 15060 19016 15116
rect 18952 15056 19016 15060
rect 19032 15116 19096 15120
rect 19032 15060 19036 15116
rect 19036 15060 19092 15116
rect 19092 15060 19096 15116
rect 19032 15056 19096 15060
rect 19112 15116 19176 15120
rect 19112 15060 19116 15116
rect 19116 15060 19172 15116
rect 19172 15060 19176 15116
rect 19112 15056 19176 15060
rect 3512 14572 3576 14576
rect 3512 14516 3516 14572
rect 3516 14516 3572 14572
rect 3572 14516 3576 14572
rect 3512 14512 3576 14516
rect 3592 14572 3656 14576
rect 3592 14516 3596 14572
rect 3596 14516 3652 14572
rect 3652 14516 3656 14572
rect 3592 14512 3656 14516
rect 3672 14572 3736 14576
rect 3672 14516 3676 14572
rect 3676 14516 3732 14572
rect 3732 14516 3736 14572
rect 3672 14512 3736 14516
rect 3752 14572 3816 14576
rect 3752 14516 3756 14572
rect 3756 14516 3812 14572
rect 3812 14516 3816 14572
rect 3752 14512 3816 14516
rect 18872 14028 18936 14032
rect 18872 13972 18876 14028
rect 18876 13972 18932 14028
rect 18932 13972 18936 14028
rect 18872 13968 18936 13972
rect 18952 14028 19016 14032
rect 18952 13972 18956 14028
rect 18956 13972 19012 14028
rect 19012 13972 19016 14028
rect 18952 13968 19016 13972
rect 19032 14028 19096 14032
rect 19032 13972 19036 14028
rect 19036 13972 19092 14028
rect 19092 13972 19096 14028
rect 19032 13968 19096 13972
rect 19112 14028 19176 14032
rect 19112 13972 19116 14028
rect 19116 13972 19172 14028
rect 19172 13972 19176 14028
rect 19112 13968 19176 13972
rect 3512 13484 3576 13488
rect 3512 13428 3516 13484
rect 3516 13428 3572 13484
rect 3572 13428 3576 13484
rect 3512 13424 3576 13428
rect 3592 13484 3656 13488
rect 3592 13428 3596 13484
rect 3596 13428 3652 13484
rect 3652 13428 3656 13484
rect 3592 13424 3656 13428
rect 3672 13484 3736 13488
rect 3672 13428 3676 13484
rect 3676 13428 3732 13484
rect 3732 13428 3736 13484
rect 3672 13424 3736 13428
rect 3752 13484 3816 13488
rect 3752 13428 3756 13484
rect 3756 13428 3812 13484
rect 3812 13428 3816 13484
rect 3752 13424 3816 13428
rect 18872 12940 18936 12944
rect 18872 12884 18876 12940
rect 18876 12884 18932 12940
rect 18932 12884 18936 12940
rect 18872 12880 18936 12884
rect 18952 12940 19016 12944
rect 18952 12884 18956 12940
rect 18956 12884 19012 12940
rect 19012 12884 19016 12940
rect 18952 12880 19016 12884
rect 19032 12940 19096 12944
rect 19032 12884 19036 12940
rect 19036 12884 19092 12940
rect 19092 12884 19096 12940
rect 19032 12880 19096 12884
rect 19112 12940 19176 12944
rect 19112 12884 19116 12940
rect 19116 12884 19172 12940
rect 19172 12884 19176 12940
rect 19112 12880 19176 12884
rect 3512 12396 3576 12400
rect 3512 12340 3516 12396
rect 3516 12340 3572 12396
rect 3572 12340 3576 12396
rect 3512 12336 3576 12340
rect 3592 12396 3656 12400
rect 3592 12340 3596 12396
rect 3596 12340 3652 12396
rect 3652 12340 3656 12396
rect 3592 12336 3656 12340
rect 3672 12396 3736 12400
rect 3672 12340 3676 12396
rect 3676 12340 3732 12396
rect 3732 12340 3736 12396
rect 3672 12336 3736 12340
rect 3752 12396 3816 12400
rect 3752 12340 3756 12396
rect 3756 12340 3812 12396
rect 3812 12340 3816 12396
rect 3752 12336 3816 12340
rect 18872 11852 18936 11856
rect 18872 11796 18876 11852
rect 18876 11796 18932 11852
rect 18932 11796 18936 11852
rect 18872 11792 18936 11796
rect 18952 11852 19016 11856
rect 18952 11796 18956 11852
rect 18956 11796 19012 11852
rect 19012 11796 19016 11852
rect 18952 11792 19016 11796
rect 19032 11852 19096 11856
rect 19032 11796 19036 11852
rect 19036 11796 19092 11852
rect 19092 11796 19096 11852
rect 19032 11792 19096 11796
rect 19112 11852 19176 11856
rect 19112 11796 19116 11852
rect 19116 11796 19172 11852
rect 19172 11796 19176 11852
rect 19112 11792 19176 11796
rect 3512 11308 3576 11312
rect 3512 11252 3516 11308
rect 3516 11252 3572 11308
rect 3572 11252 3576 11308
rect 3512 11248 3576 11252
rect 3592 11308 3656 11312
rect 3592 11252 3596 11308
rect 3596 11252 3652 11308
rect 3652 11252 3656 11308
rect 3592 11248 3656 11252
rect 3672 11308 3736 11312
rect 3672 11252 3676 11308
rect 3676 11252 3732 11308
rect 3732 11252 3736 11308
rect 3672 11248 3736 11252
rect 3752 11308 3816 11312
rect 3752 11252 3756 11308
rect 3756 11252 3812 11308
rect 3812 11252 3816 11308
rect 3752 11248 3816 11252
rect 18872 10764 18936 10768
rect 18872 10708 18876 10764
rect 18876 10708 18932 10764
rect 18932 10708 18936 10764
rect 18872 10704 18936 10708
rect 18952 10764 19016 10768
rect 18952 10708 18956 10764
rect 18956 10708 19012 10764
rect 19012 10708 19016 10764
rect 18952 10704 19016 10708
rect 19032 10764 19096 10768
rect 19032 10708 19036 10764
rect 19036 10708 19092 10764
rect 19092 10708 19096 10764
rect 19032 10704 19096 10708
rect 19112 10764 19176 10768
rect 19112 10708 19116 10764
rect 19116 10708 19172 10764
rect 19172 10708 19176 10764
rect 19112 10704 19176 10708
rect 3512 10220 3576 10224
rect 3512 10164 3516 10220
rect 3516 10164 3572 10220
rect 3572 10164 3576 10220
rect 3512 10160 3576 10164
rect 3592 10220 3656 10224
rect 3592 10164 3596 10220
rect 3596 10164 3652 10220
rect 3652 10164 3656 10220
rect 3592 10160 3656 10164
rect 3672 10220 3736 10224
rect 3672 10164 3676 10220
rect 3676 10164 3732 10220
rect 3732 10164 3736 10220
rect 3672 10160 3736 10164
rect 3752 10220 3816 10224
rect 3752 10164 3756 10220
rect 3756 10164 3812 10220
rect 3812 10164 3816 10220
rect 3752 10160 3816 10164
rect 18872 9676 18936 9680
rect 18872 9620 18876 9676
rect 18876 9620 18932 9676
rect 18932 9620 18936 9676
rect 18872 9616 18936 9620
rect 18952 9676 19016 9680
rect 18952 9620 18956 9676
rect 18956 9620 19012 9676
rect 19012 9620 19016 9676
rect 18952 9616 19016 9620
rect 19032 9676 19096 9680
rect 19032 9620 19036 9676
rect 19036 9620 19092 9676
rect 19092 9620 19096 9676
rect 19032 9616 19096 9620
rect 19112 9676 19176 9680
rect 19112 9620 19116 9676
rect 19116 9620 19172 9676
rect 19172 9620 19176 9676
rect 19112 9616 19176 9620
rect 3512 9132 3576 9136
rect 3512 9076 3516 9132
rect 3516 9076 3572 9132
rect 3572 9076 3576 9132
rect 3512 9072 3576 9076
rect 3592 9132 3656 9136
rect 3592 9076 3596 9132
rect 3596 9076 3652 9132
rect 3652 9076 3656 9132
rect 3592 9072 3656 9076
rect 3672 9132 3736 9136
rect 3672 9076 3676 9132
rect 3676 9076 3732 9132
rect 3732 9076 3736 9132
rect 3672 9072 3736 9076
rect 3752 9132 3816 9136
rect 3752 9076 3756 9132
rect 3756 9076 3812 9132
rect 3812 9076 3816 9132
rect 3752 9072 3816 9076
rect 18872 8588 18936 8592
rect 18872 8532 18876 8588
rect 18876 8532 18932 8588
rect 18932 8532 18936 8588
rect 18872 8528 18936 8532
rect 18952 8588 19016 8592
rect 18952 8532 18956 8588
rect 18956 8532 19012 8588
rect 19012 8532 19016 8588
rect 18952 8528 19016 8532
rect 19032 8588 19096 8592
rect 19032 8532 19036 8588
rect 19036 8532 19092 8588
rect 19092 8532 19096 8588
rect 19032 8528 19096 8532
rect 19112 8588 19176 8592
rect 19112 8532 19116 8588
rect 19116 8532 19172 8588
rect 19172 8532 19176 8588
rect 19112 8528 19176 8532
rect 3512 8044 3576 8048
rect 3512 7988 3516 8044
rect 3516 7988 3572 8044
rect 3572 7988 3576 8044
rect 3512 7984 3576 7988
rect 3592 8044 3656 8048
rect 3592 7988 3596 8044
rect 3596 7988 3652 8044
rect 3652 7988 3656 8044
rect 3592 7984 3656 7988
rect 3672 8044 3736 8048
rect 3672 7988 3676 8044
rect 3676 7988 3732 8044
rect 3732 7988 3736 8044
rect 3672 7984 3736 7988
rect 3752 8044 3816 8048
rect 3752 7988 3756 8044
rect 3756 7988 3812 8044
rect 3812 7988 3816 8044
rect 3752 7984 3816 7988
rect 18872 7500 18936 7504
rect 18872 7444 18876 7500
rect 18876 7444 18932 7500
rect 18932 7444 18936 7500
rect 18872 7440 18936 7444
rect 18952 7500 19016 7504
rect 18952 7444 18956 7500
rect 18956 7444 19012 7500
rect 19012 7444 19016 7500
rect 18952 7440 19016 7444
rect 19032 7500 19096 7504
rect 19032 7444 19036 7500
rect 19036 7444 19092 7500
rect 19092 7444 19096 7500
rect 19032 7440 19096 7444
rect 19112 7500 19176 7504
rect 19112 7444 19116 7500
rect 19116 7444 19172 7500
rect 19172 7444 19176 7500
rect 19112 7440 19176 7444
rect 3512 6956 3576 6960
rect 3512 6900 3516 6956
rect 3516 6900 3572 6956
rect 3572 6900 3576 6956
rect 3512 6896 3576 6900
rect 3592 6956 3656 6960
rect 3592 6900 3596 6956
rect 3596 6900 3652 6956
rect 3652 6900 3656 6956
rect 3592 6896 3656 6900
rect 3672 6956 3736 6960
rect 3672 6900 3676 6956
rect 3676 6900 3732 6956
rect 3732 6900 3736 6956
rect 3672 6896 3736 6900
rect 3752 6956 3816 6960
rect 3752 6900 3756 6956
rect 3756 6900 3812 6956
rect 3812 6900 3816 6956
rect 3752 6896 3816 6900
rect 18872 6412 18936 6416
rect 18872 6356 18876 6412
rect 18876 6356 18932 6412
rect 18932 6356 18936 6412
rect 18872 6352 18936 6356
rect 18952 6412 19016 6416
rect 18952 6356 18956 6412
rect 18956 6356 19012 6412
rect 19012 6356 19016 6412
rect 18952 6352 19016 6356
rect 19032 6412 19096 6416
rect 19032 6356 19036 6412
rect 19036 6356 19092 6412
rect 19092 6356 19096 6412
rect 19032 6352 19096 6356
rect 19112 6412 19176 6416
rect 19112 6356 19116 6412
rect 19116 6356 19172 6412
rect 19172 6356 19176 6412
rect 19112 6352 19176 6356
rect 3512 5868 3576 5872
rect 3512 5812 3516 5868
rect 3516 5812 3572 5868
rect 3572 5812 3576 5868
rect 3512 5808 3576 5812
rect 3592 5868 3656 5872
rect 3592 5812 3596 5868
rect 3596 5812 3652 5868
rect 3652 5812 3656 5868
rect 3592 5808 3656 5812
rect 3672 5868 3736 5872
rect 3672 5812 3676 5868
rect 3676 5812 3732 5868
rect 3732 5812 3736 5868
rect 3672 5808 3736 5812
rect 3752 5868 3816 5872
rect 3752 5812 3756 5868
rect 3756 5812 3812 5868
rect 3812 5812 3816 5868
rect 3752 5808 3816 5812
rect 18872 5324 18936 5328
rect 18872 5268 18876 5324
rect 18876 5268 18932 5324
rect 18932 5268 18936 5324
rect 18872 5264 18936 5268
rect 18952 5324 19016 5328
rect 18952 5268 18956 5324
rect 18956 5268 19012 5324
rect 19012 5268 19016 5324
rect 18952 5264 19016 5268
rect 19032 5324 19096 5328
rect 19032 5268 19036 5324
rect 19036 5268 19092 5324
rect 19092 5268 19096 5324
rect 19032 5264 19096 5268
rect 19112 5324 19176 5328
rect 19112 5268 19116 5324
rect 19116 5268 19172 5324
rect 19172 5268 19176 5324
rect 19112 5264 19176 5268
rect 3512 4780 3576 4784
rect 3512 4724 3516 4780
rect 3516 4724 3572 4780
rect 3572 4724 3576 4780
rect 3512 4720 3576 4724
rect 3592 4780 3656 4784
rect 3592 4724 3596 4780
rect 3596 4724 3652 4780
rect 3652 4724 3656 4780
rect 3592 4720 3656 4724
rect 3672 4780 3736 4784
rect 3672 4724 3676 4780
rect 3676 4724 3732 4780
rect 3732 4724 3736 4780
rect 3672 4720 3736 4724
rect 3752 4780 3816 4784
rect 3752 4724 3756 4780
rect 3756 4724 3812 4780
rect 3812 4724 3816 4780
rect 3752 4720 3816 4724
rect 18872 4236 18936 4240
rect 18872 4180 18876 4236
rect 18876 4180 18932 4236
rect 18932 4180 18936 4236
rect 18872 4176 18936 4180
rect 18952 4236 19016 4240
rect 18952 4180 18956 4236
rect 18956 4180 19012 4236
rect 19012 4180 19016 4236
rect 18952 4176 19016 4180
rect 19032 4236 19096 4240
rect 19032 4180 19036 4236
rect 19036 4180 19092 4236
rect 19092 4180 19096 4236
rect 19032 4176 19096 4180
rect 19112 4236 19176 4240
rect 19112 4180 19116 4236
rect 19116 4180 19172 4236
rect 19172 4180 19176 4236
rect 19112 4176 19176 4180
rect 3512 3692 3576 3696
rect 3512 3636 3516 3692
rect 3516 3636 3572 3692
rect 3572 3636 3576 3692
rect 3512 3632 3576 3636
rect 3592 3692 3656 3696
rect 3592 3636 3596 3692
rect 3596 3636 3652 3692
rect 3652 3636 3656 3692
rect 3592 3632 3656 3636
rect 3672 3692 3736 3696
rect 3672 3636 3676 3692
rect 3676 3636 3732 3692
rect 3732 3636 3736 3692
rect 3672 3632 3736 3636
rect 3752 3692 3816 3696
rect 3752 3636 3756 3692
rect 3756 3636 3812 3692
rect 3812 3636 3816 3692
rect 3752 3632 3816 3636
rect 18872 3148 18936 3152
rect 18872 3092 18876 3148
rect 18876 3092 18932 3148
rect 18932 3092 18936 3148
rect 18872 3088 18936 3092
rect 18952 3148 19016 3152
rect 18952 3092 18956 3148
rect 18956 3092 19012 3148
rect 19012 3092 19016 3148
rect 18952 3088 19016 3092
rect 19032 3148 19096 3152
rect 19032 3092 19036 3148
rect 19036 3092 19092 3148
rect 19092 3092 19096 3148
rect 19032 3088 19096 3092
rect 19112 3148 19176 3152
rect 19112 3092 19116 3148
rect 19116 3092 19172 3148
rect 19172 3092 19176 3148
rect 19112 3088 19176 3092
rect 3512 2604 3576 2608
rect 3512 2548 3516 2604
rect 3516 2548 3572 2604
rect 3572 2548 3576 2604
rect 3512 2544 3576 2548
rect 3592 2604 3656 2608
rect 3592 2548 3596 2604
rect 3596 2548 3652 2604
rect 3652 2548 3656 2604
rect 3592 2544 3656 2548
rect 3672 2604 3736 2608
rect 3672 2548 3676 2604
rect 3676 2548 3732 2604
rect 3732 2548 3736 2604
rect 3672 2544 3736 2548
rect 3752 2604 3816 2608
rect 3752 2548 3756 2604
rect 3756 2548 3812 2604
rect 3812 2548 3816 2604
rect 3752 2544 3816 2548
rect 18872 2060 18936 2064
rect 18872 2004 18876 2060
rect 18876 2004 18932 2060
rect 18932 2004 18936 2060
rect 18872 2000 18936 2004
rect 18952 2060 19016 2064
rect 18952 2004 18956 2060
rect 18956 2004 19012 2060
rect 19012 2004 19016 2060
rect 18952 2000 19016 2004
rect 19032 2060 19096 2064
rect 19032 2004 19036 2060
rect 19036 2004 19092 2060
rect 19092 2004 19096 2060
rect 19032 2000 19096 2004
rect 19112 2060 19176 2064
rect 19112 2004 19116 2060
rect 19116 2004 19172 2060
rect 19172 2004 19176 2060
rect 19112 2000 19176 2004
rect 3512 1516 3576 1520
rect 3512 1460 3516 1516
rect 3516 1460 3572 1516
rect 3572 1460 3576 1516
rect 3512 1456 3576 1460
rect 3592 1516 3656 1520
rect 3592 1460 3596 1516
rect 3596 1460 3652 1516
rect 3652 1460 3656 1516
rect 3592 1456 3656 1460
rect 3672 1516 3736 1520
rect 3672 1460 3676 1516
rect 3676 1460 3732 1516
rect 3732 1460 3736 1516
rect 3672 1456 3736 1460
rect 3752 1516 3816 1520
rect 3752 1460 3756 1516
rect 3756 1460 3812 1516
rect 3812 1460 3816 1516
rect 3752 1456 3816 1460
rect 31636 980 31700 1044
rect 18872 972 18936 976
rect 18872 916 18876 972
rect 18876 916 18932 972
rect 18932 916 18936 972
rect 18872 912 18936 916
rect 18952 972 19016 976
rect 18952 916 18956 972
rect 18956 916 19012 972
rect 19012 916 19016 972
rect 18952 912 19016 916
rect 19032 972 19096 976
rect 19032 916 19036 972
rect 19036 916 19092 972
rect 19092 916 19096 972
rect 19032 912 19096 916
rect 19112 972 19176 976
rect 19112 916 19116 972
rect 19116 916 19172 972
rect 19172 916 19176 972
rect 19112 912 19176 916
rect 31636 708 31700 772
rect 3512 428 3576 432
rect 3512 372 3516 428
rect 3516 372 3572 428
rect 3572 372 3576 428
rect 3512 368 3576 372
rect 3592 428 3656 432
rect 3592 372 3596 428
rect 3596 372 3652 428
rect 3652 372 3656 428
rect 3592 368 3656 372
rect 3672 428 3736 432
rect 3672 372 3676 428
rect 3676 372 3732 428
rect 3732 372 3736 428
rect 3672 368 3736 372
rect 3752 428 3816 432
rect 3752 372 3756 428
rect 3756 372 3812 428
rect 3812 372 3816 428
rect 3752 368 3816 372
<< metal4 >>
rect 18864 31440 19184 31456
rect 3504 30896 3824 31408
rect 3504 30832 3512 30896
rect 3576 30832 3592 30896
rect 3656 30832 3672 30896
rect 3736 30832 3752 30896
rect 3816 30832 3824 30896
rect 3504 29808 3824 30832
rect 3504 29744 3512 29808
rect 3576 29744 3592 29808
rect 3656 29744 3672 29808
rect 3736 29744 3752 29808
rect 3816 29744 3824 29808
rect 3504 28720 3824 29744
rect 3504 28656 3512 28720
rect 3576 28656 3592 28720
rect 3656 28656 3672 28720
rect 3736 28656 3752 28720
rect 3816 28656 3824 28720
rect 3504 27632 3824 28656
rect 3504 27568 3512 27632
rect 3576 27568 3592 27632
rect 3656 27568 3672 27632
rect 3736 27568 3752 27632
rect 3816 27568 3824 27632
rect 3504 26544 3824 27568
rect 3504 26480 3512 26544
rect 3576 26480 3592 26544
rect 3656 26480 3672 26544
rect 3736 26480 3752 26544
rect 3816 26480 3824 26544
rect 3504 25456 3824 26480
rect 3504 25392 3512 25456
rect 3576 25392 3592 25456
rect 3656 25392 3672 25456
rect 3736 25392 3752 25456
rect 3816 25392 3824 25456
rect 3504 24368 3824 25392
rect 3504 24304 3512 24368
rect 3576 24304 3592 24368
rect 3656 24304 3672 24368
rect 3736 24304 3752 24368
rect 3816 24304 3824 24368
rect 3504 23280 3824 24304
rect 3504 23216 3512 23280
rect 3576 23216 3592 23280
rect 3656 23216 3672 23280
rect 3736 23216 3752 23280
rect 3816 23216 3824 23280
rect 3504 22192 3824 23216
rect 3504 22128 3512 22192
rect 3576 22128 3592 22192
rect 3656 22128 3672 22192
rect 3736 22128 3752 22192
rect 3816 22128 3824 22192
rect 3504 21104 3824 22128
rect 3504 21040 3512 21104
rect 3576 21040 3592 21104
rect 3656 21040 3672 21104
rect 3736 21040 3752 21104
rect 3816 21040 3824 21104
rect 3504 20016 3824 21040
rect 3504 19952 3512 20016
rect 3576 19952 3592 20016
rect 3656 19952 3672 20016
rect 3736 19952 3752 20016
rect 3816 19952 3824 20016
rect 3504 18928 3824 19952
rect 3504 18864 3512 18928
rect 3576 18864 3592 18928
rect 3656 18864 3672 18928
rect 3736 18864 3752 18928
rect 3816 18864 3824 18928
rect 3504 17840 3824 18864
rect 3504 17776 3512 17840
rect 3576 17776 3592 17840
rect 3656 17776 3672 17840
rect 3736 17776 3752 17840
rect 3816 17776 3824 17840
rect 3504 16752 3824 17776
rect 3504 16688 3512 16752
rect 3576 16688 3592 16752
rect 3656 16688 3672 16752
rect 3736 16688 3752 16752
rect 3816 16688 3824 16752
rect 3504 15664 3824 16688
rect 3504 15600 3512 15664
rect 3576 15600 3592 15664
rect 3656 15600 3672 15664
rect 3736 15600 3752 15664
rect 3816 15600 3824 15664
rect 3504 14576 3824 15600
rect 3504 14512 3512 14576
rect 3576 14512 3592 14576
rect 3656 14512 3672 14576
rect 3736 14512 3752 14576
rect 3816 14512 3824 14576
rect 3504 13488 3824 14512
rect 3504 13424 3512 13488
rect 3576 13424 3592 13488
rect 3656 13424 3672 13488
rect 3736 13424 3752 13488
rect 3816 13424 3824 13488
rect 3504 12400 3824 13424
rect 3504 12336 3512 12400
rect 3576 12336 3592 12400
rect 3656 12336 3672 12400
rect 3736 12336 3752 12400
rect 3816 12336 3824 12400
rect 3504 11312 3824 12336
rect 3504 11248 3512 11312
rect 3576 11248 3592 11312
rect 3656 11248 3672 11312
rect 3736 11248 3752 11312
rect 3816 11248 3824 11312
rect 3504 10224 3824 11248
rect 3504 10160 3512 10224
rect 3576 10160 3592 10224
rect 3656 10160 3672 10224
rect 3736 10160 3752 10224
rect 3816 10160 3824 10224
rect 3504 9136 3824 10160
rect 3504 9072 3512 9136
rect 3576 9072 3592 9136
rect 3656 9072 3672 9136
rect 3736 9072 3752 9136
rect 3816 9072 3824 9136
rect 3504 8048 3824 9072
rect 3504 7984 3512 8048
rect 3576 7984 3592 8048
rect 3656 7984 3672 8048
rect 3736 7984 3752 8048
rect 3816 7984 3824 8048
rect 3504 6960 3824 7984
rect 3504 6896 3512 6960
rect 3576 6896 3592 6960
rect 3656 6896 3672 6960
rect 3736 6896 3752 6960
rect 3816 6896 3824 6960
rect 3504 5872 3824 6896
rect 3504 5808 3512 5872
rect 3576 5808 3592 5872
rect 3656 5808 3672 5872
rect 3736 5808 3752 5872
rect 3816 5808 3824 5872
rect 3504 4784 3824 5808
rect 3504 4720 3512 4784
rect 3576 4720 3592 4784
rect 3656 4720 3672 4784
rect 3736 4720 3752 4784
rect 3816 4720 3824 4784
rect 3504 3848 3824 4720
rect 3504 3696 3546 3848
rect 3782 3696 3824 3848
rect 3504 3632 3512 3696
rect 3816 3632 3824 3696
rect 3504 3612 3546 3632
rect 3782 3612 3824 3632
rect 3504 2608 3824 3612
rect 3504 2544 3512 2608
rect 3576 2544 3592 2608
rect 3656 2544 3672 2608
rect 3736 2544 3752 2608
rect 3816 2544 3824 2608
rect 3504 1520 3824 2544
rect 3504 1456 3512 1520
rect 3576 1456 3592 1520
rect 3656 1456 3672 1520
rect 3736 1456 3752 1520
rect 3816 1456 3824 1520
rect 3504 432 3824 1456
rect 3504 368 3512 432
rect 3576 368 3592 432
rect 3656 368 3672 432
rect 3736 368 3752 432
rect 3816 368 3824 432
rect 18864 31376 18872 31440
rect 18936 31376 18952 31440
rect 19016 31376 19032 31440
rect 19096 31376 19112 31440
rect 19176 31376 19184 31440
rect 18864 30352 19184 31376
rect 18864 30288 18872 30352
rect 18936 30288 18952 30352
rect 19016 30288 19032 30352
rect 19096 30288 19112 30352
rect 19176 30288 19184 30352
rect 18864 29264 19184 30288
rect 18864 29200 18872 29264
rect 18936 29200 18952 29264
rect 19016 29200 19032 29264
rect 19096 29200 19112 29264
rect 19176 29200 19184 29264
rect 18864 28176 19184 29200
rect 18864 28112 18872 28176
rect 18936 28112 18952 28176
rect 19016 28112 19032 28176
rect 19096 28112 19112 28176
rect 19176 28112 19184 28176
rect 18864 27088 19184 28112
rect 18864 27024 18872 27088
rect 18936 27024 18952 27088
rect 19016 27024 19032 27088
rect 19096 27024 19112 27088
rect 19176 27024 19184 27088
rect 18864 26000 19184 27024
rect 18864 25936 18872 26000
rect 18936 25936 18952 26000
rect 19016 25936 19032 26000
rect 19096 25936 19112 26000
rect 19176 25936 19184 26000
rect 18864 24912 19184 25936
rect 18864 24848 18872 24912
rect 18936 24848 18952 24912
rect 19016 24848 19032 24912
rect 19096 24848 19112 24912
rect 19176 24848 19184 24912
rect 18864 23824 19184 24848
rect 18864 23760 18872 23824
rect 18936 23760 18952 23824
rect 19016 23760 19032 23824
rect 19096 23760 19112 23824
rect 19176 23760 19184 23824
rect 18864 22736 19184 23760
rect 18864 22672 18872 22736
rect 18936 22672 18952 22736
rect 19016 22672 19032 22736
rect 19096 22672 19112 22736
rect 19176 22672 19184 22736
rect 18864 21648 19184 22672
rect 18864 21584 18872 21648
rect 18936 21584 18952 21648
rect 19016 21584 19032 21648
rect 19096 21584 19112 21648
rect 19176 21584 19184 21648
rect 18864 20560 19184 21584
rect 18864 20496 18872 20560
rect 18936 20496 18952 20560
rect 19016 20496 19032 20560
rect 19096 20496 19112 20560
rect 19176 20496 19184 20560
rect 18864 19472 19184 20496
rect 18864 19408 18872 19472
rect 18936 19408 18952 19472
rect 19016 19408 19032 19472
rect 19096 19408 19112 19472
rect 19176 19408 19184 19472
rect 18864 19166 19184 19408
rect 18864 18930 18906 19166
rect 19142 18930 19184 19166
rect 18864 18384 19184 18930
rect 18864 18320 18872 18384
rect 18936 18320 18952 18384
rect 19016 18320 19032 18384
rect 19096 18320 19112 18384
rect 19176 18320 19184 18384
rect 18864 17296 19184 18320
rect 18864 17232 18872 17296
rect 18936 17232 18952 17296
rect 19016 17232 19032 17296
rect 19096 17232 19112 17296
rect 19176 17232 19184 17296
rect 18864 16208 19184 17232
rect 18864 16144 18872 16208
rect 18936 16144 18952 16208
rect 19016 16144 19032 16208
rect 19096 16144 19112 16208
rect 19176 16144 19184 16208
rect 18864 15120 19184 16144
rect 18864 15056 18872 15120
rect 18936 15056 18952 15120
rect 19016 15056 19032 15120
rect 19096 15056 19112 15120
rect 19176 15056 19184 15120
rect 18864 14032 19184 15056
rect 18864 13968 18872 14032
rect 18936 13968 18952 14032
rect 19016 13968 19032 14032
rect 19096 13968 19112 14032
rect 19176 13968 19184 14032
rect 18864 12944 19184 13968
rect 18864 12880 18872 12944
rect 18936 12880 18952 12944
rect 19016 12880 19032 12944
rect 19096 12880 19112 12944
rect 19176 12880 19184 12944
rect 18864 11856 19184 12880
rect 18864 11792 18872 11856
rect 18936 11792 18952 11856
rect 19016 11792 19032 11856
rect 19096 11792 19112 11856
rect 19176 11792 19184 11856
rect 18864 10768 19184 11792
rect 18864 10704 18872 10768
rect 18936 10704 18952 10768
rect 19016 10704 19032 10768
rect 19096 10704 19112 10768
rect 19176 10704 19184 10768
rect 18864 9680 19184 10704
rect 18864 9616 18872 9680
rect 18936 9616 18952 9680
rect 19016 9616 19032 9680
rect 19096 9616 19112 9680
rect 19176 9616 19184 9680
rect 18864 8592 19184 9616
rect 18864 8528 18872 8592
rect 18936 8528 18952 8592
rect 19016 8528 19032 8592
rect 19096 8528 19112 8592
rect 19176 8528 19184 8592
rect 18864 7504 19184 8528
rect 18864 7440 18872 7504
rect 18936 7440 18952 7504
rect 19016 7440 19032 7504
rect 19096 7440 19112 7504
rect 19176 7440 19184 7504
rect 18864 6416 19184 7440
rect 18864 6352 18872 6416
rect 18936 6352 18952 6416
rect 19016 6352 19032 6416
rect 19096 6352 19112 6416
rect 19176 6352 19184 6416
rect 18864 5328 19184 6352
rect 18864 5264 18872 5328
rect 18936 5264 18952 5328
rect 19016 5264 19032 5328
rect 19096 5264 19112 5328
rect 19176 5264 19184 5328
rect 18864 4240 19184 5264
rect 18864 4176 18872 4240
rect 18936 4176 18952 4240
rect 19016 4176 19032 4240
rect 19096 4176 19112 4240
rect 19176 4176 19184 4240
rect 18864 3152 19184 4176
rect 18864 3088 18872 3152
rect 18936 3088 18952 3152
rect 19016 3088 19032 3152
rect 19096 3088 19112 3152
rect 19176 3088 19184 3152
rect 18864 2064 19184 3088
rect 18864 2000 18872 2064
rect 18936 2000 18952 2064
rect 19016 2000 19032 2064
rect 19096 2000 19112 2064
rect 19176 2000 19184 2064
rect 18864 976 19184 2000
rect 31635 1044 31701 1045
rect 31635 980 31636 1044
rect 31700 980 31701 1044
rect 31635 979 31701 980
rect 18864 912 18872 976
rect 18936 912 18952 976
rect 19016 912 19032 976
rect 19096 912 19112 976
rect 19176 912 19184 976
rect 18864 400 19184 912
rect 31638 773 31698 979
rect 31635 772 31701 773
rect 31635 708 31636 772
rect 31700 708 31701 772
rect 31635 707 31701 708
rect 3504 352 3824 368
<< via4 >>
rect 3546 3696 3782 3848
rect 3546 3632 3576 3696
rect 3576 3632 3592 3696
rect 3592 3632 3656 3696
rect 3656 3632 3672 3696
rect 3672 3632 3736 3696
rect 3736 3632 3752 3696
rect 3752 3632 3782 3696
rect 3546 3612 3782 3632
rect 18906 18930 19142 19166
<< metal5 >>
rect 400 19166 31680 19208
rect 400 18930 18906 19166
rect 19142 18930 31680 19166
rect 400 18888 31680 18930
rect 400 3848 31680 3890
rect 400 3612 3546 3848
rect 3782 3612 31680 3848
rect 400 3570 31680 3612
use sky130_fd_sc_hd__decap_12  FILL1380x0 ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 676 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_2 ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 400 0 1 944
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL1380x2720
timestamp 1586547711
transform 1 0 676 0 1 944
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1586547711
transform 1 0 400 0 -1 944
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL3680x2720 ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 1136 0 1 944
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_175 ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 952 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL8740x2720
timestamp 1586547711
transform 1 0 2148 0 1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL6900x0
timestamp 1586547711
transform 1 0 1780 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_183
timestamp 1586547711
transform 1 0 1964 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL7360x2720 ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 1872 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL14720x0
timestamp 1586547711
transform 1 0 3344 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_184
timestamp 1586547711
transform 1 0 3620 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL14260x2720
timestamp 1586547711
transform 1 0 3252 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114 ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 3252 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL12420x0 ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 2884 0 -1 944
box 0 -48 368 592
use sky130_fd_sc_hd__conb_1  _847_ ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 3344 0 1 944
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL21160x2720
timestamp 1586547711
transform 1 0 4632 0 1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL20240x0
timestamp 1586547711
transform 1 0 4448 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_288
timestamp 1586547711
transform 1 0 3896 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_467
timestamp 1586547711
transform 1 0 4080 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1491
timestamp 1586547711
transform 1 0 4264 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1667
timestamp 1586547711
transform 1 0 4448 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL17020x2720
timestamp 1586547711
transform 1 0 3804 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL28980x0
timestamp 1586547711
transform 1 0 6196 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL26680x2720
timestamp 1586547711
transform 1 0 5736 0 1 944
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1490
timestamp 1586547711
transform 1 0 6748 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1587
timestamp 1586547711
transform 1 0 6932 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL31280x2720
timestamp 1586547711
transform 1 0 6656 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1586547711
transform 1 0 6012 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1586547711
transform 1 0 6104 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL28520x2720 ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 6104 0 1 944
box 0 -48 552 592
use sky130_fd_sc_hd__decap_6  FILL25760x0
timestamp 1586547711
transform 1 0 5552 0 -1 944
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL33580x2720
timestamp 1586547711
transform 1 0 7116 0 1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL39100x2720
timestamp 1586547711
transform 1 0 8220 0 1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL34500x0
timestamp 1586547711
transform 1 0 7300 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL43240x0
timestamp 1586547711
transform 1 0 9048 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1586547711
transform 1 0 8956 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL40020x0
timestamp 1586547711
transform 1 0 8404 0 -1 944
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL50140x2720
timestamp 1586547711
transform 1 0 10428 0 1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL48760x0
timestamp 1586547711
transform 1 0 10152 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1586547711
transform 1 0 9692 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_78
timestamp 1586547711
transform 1 0 9876 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_349
timestamp 1586547711
transform 1 0 10060 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1654
timestamp 1586547711
transform 1 0 10244 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL44620x2720
timestamp 1586547711
transform 1 0 9324 0 1 944
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILL54280x0
timestamp 1586547711
transform 1 0 11256 0 -1 944
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL61640x2720
timestamp 1586547711
transform 1 0 12728 0 1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL57500x0
timestamp 1586547711
transform 1 0 11900 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL63020x0
timestamp 1586547711
transform 1 0 13004 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL56580x2720
timestamp 1586547711
transform 1 0 11716 0 1 944
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_177
timestamp 1586547711
transform 1 0 12544 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL55660x2720
timestamp 1586547711
transform 1 0 11532 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL60260x2720
timestamp 1586547711
transform 1 0 12452 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1586547711
transform 1 0 11624 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1586547711
transform 1 0 11808 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL67160x2720
timestamp 1586547711
transform 1 0 13832 0 1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL73600x2720
timestamp 1586547711
transform 1 0 15120 0 1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL71760x0
timestamp 1586547711
transform 1 0 14752 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL77280x0
timestamp 1586547711
transform 1 0 15856 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_187
timestamp 1586547711
transform 1 0 14936 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1586547711
transform 1 0 14660 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL68540x0
timestamp 1586547711
transform 1 0 14108 0 -1 944
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILL79120x2720
timestamp 1586547711
transform 1 0 16224 0 1 944
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_171
timestamp 1586547711
transform 1 0 16500 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL81420x2720
timestamp 1586547711
transform 1 0 16684 0 1 944
box 0 -48 552 592
use sky130_fd_sc_hd__decap_6  FILL82800x0
timestamp 1586547711
transform 1 0 16960 0 -1 944
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL86020x0
timestamp 1586547711
transform 1 0 17604 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1501
timestamp 1586547711
transform 1 0 17880 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_86
timestamp 1586547711
transform 1 0 18064 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1586547711
transform 1 0 17236 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1586547711
transform 1 0 17512 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL84640x2720
timestamp 1586547711
transform 1 0 17328 0 1 944
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_384
timestamp 1586547711
transform 1 0 18248 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_927
timestamp 1586547711
transform 1 0 18432 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1023
timestamp 1586547711
transform 1 0 18616 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_386
timestamp 1586547711
transform 1 0 18800 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_83
timestamp 1586547711
transform 1 0 18984 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_784
timestamp 1586547711
transform 1 0 19168 0 -1 944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL93380x0
timestamp 1586547711
transform 1 0 19076 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL91540x0
timestamp 1586547711
transform 1 0 18708 0 -1 944
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILL95680x0
timestamp 1586547711
transform 1 0 19536 0 -1 944
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1502
timestamp 1586547711
transform 1 0 19352 0 -1 944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL99360x0
timestamp 1586547711
transform 1 0 20272 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _762_ ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 19168 0 1 944
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL103960x2720
timestamp 1586547711
transform 1 0 21192 0 1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL100280x0
timestamp 1586547711
transform 1 0 20456 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1586547711
transform 1 0 20456 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_84
timestamp 1586547711
transform 1 0 20640 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_387
timestamp 1586547711
transform 1 0 20824 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1652
timestamp 1586547711
transform 1 0 21008 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1586547711
transform 1 0 20364 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL105800x0
timestamp 1586547711
transform 1 0 21560 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_884
timestamp 1586547711
transform 1 0 22296 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_802
timestamp 1586547711
transform 1 0 22480 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_342
timestamp 1586547711
transform 1 0 22664 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_61
timestamp 1586547711
transform 1 0 23032 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL112700x2720
timestamp 1586547711
transform 1 0 22940 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1586547711
transform 1 0 22848 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL111320x0
timestamp 1586547711
transform 1 0 22664 0 -1 944
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1586547711
transform 1 0 23216 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_63
timestamp 1586547711
transform 1 0 23400 0 -1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_343
timestamp 1586547711
transform 1 0 23584 0 -1 944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL114540x0
timestamp 1586547711
transform 1 0 23308 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1586547711
transform 1 0 23216 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL118680x0
timestamp 1586547711
transform 1 0 24136 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_890
timestamp 1586547711
transform 1 0 23768 0 -1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1660
timestamp 1586547711
transform 1 0 23952 0 -1 944
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _888_ ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 23400 0 1 944
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_12  FILL127880x2720
timestamp 1586547711
transform 1 0 25976 0 1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL128800x0
timestamp 1586547711
transform 1 0 26160 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL125580x2720
timestamp 1586547711
transform 1 0 25516 0 1 944
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL124200x0
timestamp 1586547711
transform 1 0 25240 0 -1 944
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_185
timestamp 1586547711
transform 1 0 25792 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL127880x0
timestamp 1586547711
transform 1 0 25976 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1586547711
transform 1 0 26068 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL134320x0
timestamp 1586547711
transform 1 0 27264 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1586547711
transform 1 0 27448 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_102
timestamp 1586547711
transform 1 0 27632 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_373
timestamp 1586547711
transform 1 0 27816 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1646
timestamp 1586547711
transform 1 0 28000 0 1 944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL133400x2720
timestamp 1586547711
transform 1 0 27080 0 1 944
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL140760x2720
timestamp 1586547711
transform 1 0 28552 0 1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL143060x0
timestamp 1586547711
transform 1 0 29012 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL138920x2720
timestamp 1586547711
transform 1 0 28184 0 1 944
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1586547711
transform 1 0 28460 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1586547711
transform 1 0 28920 0 -1 944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL139840x0
timestamp 1586547711
transform 1 0 28368 0 -1 944
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL146280x2720
timestamp 1586547711
transform 1 0 29656 0 1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL148580x0
timestamp 1586547711
transform 1 0 30116 0 -1 944
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL154560x2720
timestamp 1586547711
transform 1 0 31312 0 1 944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL151800x2720
timestamp 1586547711
transform 1 0 30760 0 1 944
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILL154100x0 ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 31220 0 -1 944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1586547711
transform 1 0 31404 0 1 944
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1586547711
transform 1 0 31404 0 -1 944
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1586547711
transform 1 0 400 0 -1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL1380x5440
timestamp 1586547711
transform 1 0 676 0 -1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL9200x5440
timestamp 1586547711
transform 1 0 2240 0 -1 2032
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1668
timestamp 1586547711
transform 1 0 1228 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__conb_1  _839_
timestamp 1586547711
transform 1 0 952 0 -1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__conb_1  _848_
timestamp 1586547711
transform 1 0 1964 0 -1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILL5060x5440
timestamp 1586547711
transform 1 0 1412 0 -1 2032
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILL12880x5440
timestamp 1586547711
transform 1 0 2976 0 -1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1586547711
transform 1 0 3252 0 -1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL14720x5440
timestamp 1586547711
transform 1 0 3344 0 -1 2032
box 0 -48 552 592
use sky130_fd_sc_hd__dfrtp_4  _905_
timestamp 1586547711
transform 1 0 3896 0 -1 2032
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_8  FILL28060x5440
timestamp 1586547711
transform 1 0 6012 0 -1 2032
box 0 -48 736 592
use sky130_fd_sc_hd__buf_4  _802_ ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 6748 0 -1 2032
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL34500x5440
timestamp 1586547711
transform 1 0 7300 0 -1 2032
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL42780x5440
timestamp 1586547711
transform 1 0 8956 0 -1 2032
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1645
timestamp 1586547711
transform 1 0 8036 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL41860x5440
timestamp 1586547711
transform 1 0 8772 0 -1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1586547711
transform 1 0 8864 0 -1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL39100x5440
timestamp 1586547711
transform 1 0 8220 0 -1 2032
box 0 -48 552 592
use sky130_fd_sc_hd__dfrtp_4  _883_
timestamp 1586547711
transform 1 0 9692 0 -1 2032
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_3  FILL62100x5440
timestamp 1586547711
transform 1 0 12820 0 -1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL57040x5440
timestamp 1586547711
transform 1 0 11808 0 -1 2032
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL66240x5440
timestamp 1586547711
transform 1 0 13648 0 -1 2032
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_81
timestamp 1586547711
transform 1 0 13096 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_909
timestamp 1586547711
transform 1 0 13280 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1653
timestamp 1586547711
transform 1 0 13464 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__conb_1  _838_
timestamp 1586547711
transform 1 0 12544 0 -1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL74060x5440
timestamp 1586547711
transform 1 0 15212 0 -1 2032
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL69920x5440
timestamp 1586547711
transform 1 0 14384 0 -1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1586547711
transform 1 0 14476 0 -1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL70840x5440
timestamp 1586547711
transform 1 0 14568 0 -1 2032
box 0 -48 368 592
use sky130_fd_sc_hd__conb_1  _844_
timestamp 1586547711
transform 1 0 14936 0 -1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL83260x5440
timestamp 1586547711
transform 1 0 17052 0 -1 2032
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1039
timestamp 1586547711
transform 1 0 16868 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1095
timestamp 1586547711
transform 1 0 17880 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL81880x5440
timestamp 1586547711
transform 1 0 16776 0 -1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL86940x5440
timestamp 1586547711
transform 1 0 17788 0 -1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__conb_1  _842_
timestamp 1586547711
transform 1 0 16500 0 -1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__o22a_4  _761_
timestamp 1586547711
transform 1 0 18064 0 -1 2032
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILL79580x5440
timestamp 1586547711
transform 1 0 16316 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1024
timestamp 1586547711
transform 1 0 19352 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL98900x5440
timestamp 1586547711
transform 1 0 20180 0 -1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1586547711
transform 1 0 20088 0 -1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL95680x5440
timestamp 1586547711
transform 1 0 19536 0 -1 2032
box 0 -48 552 592
use sky130_fd_sc_hd__dfstp_4  _881_ ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 20272 0 -1 2032
box 0 -48 2208 592
use sky130_fd_sc_hd__decap_8  FILL110400x5440
timestamp 1586547711
transform 1 0 22480 0 -1 2032
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILL120520x5440
timestamp 1586547711
transform 1 0 24504 0 -1 2032
box 0 -48 1104 592
use sky130_fd_sc_hd__o22a_4  _528_
timestamp 1586547711
transform 1 0 23216 0 -1 2032
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_3  FILL128340x5440
timestamp 1586547711
transform 1 0 26068 0 -1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL130640x5440
timestamp 1586547711
transform 1 0 26528 0 -1 2032
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1520
timestamp 1586547711
transform 1 0 26344 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL126040x5440
timestamp 1586547711
transform 1 0 25608 0 -1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1586547711
transform 1 0 25700 0 -1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__conb_1  _846_
timestamp 1586547711
transform 1 0 25792 0 -1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILL134320x5440
timestamp 1586547711
transform 1 0 27264 0 -1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__dfstp_4  _875_
timestamp 1586547711
transform 1 0 27448 0 -1 2032
box 0 -48 2208 592
use sky130_fd_sc_hd__decap_12  FILL146280x5440
timestamp 1586547711
transform 1 0 29656 0 -1 2032
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1586547711
transform 1 0 31312 0 -1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL151800x5440
timestamp 1586547711
transform 1 0 30760 0 -1 2032
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1586547711
transform 1 0 31404 0 -1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1586547711
transform 1 0 400 0 1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_292
timestamp 1586547711
transform 1 0 768 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL1380x8160
timestamp 1586547711
transform 1 0 676 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _906_
timestamp 1586547711
transform 1 0 952 0 1 2032
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_8  FILL21620x8160
timestamp 1586547711
transform 1 0 4724 0 1 2032
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1588
timestamp 1586547711
transform 1 0 3068 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1471
timestamp 1586547711
transform 1 0 3252 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1445
timestamp 1586547711
transform 1 0 3436 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_283
timestamp 1586547711
transform 1 0 3620 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_466
timestamp 1586547711
transform 1 0 4356 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1492
timestamp 1586547711
transform 1 0 4540 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _803_
timestamp 1586547711
transform 1 0 3804 0 1 2032
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_284
timestamp 1586547711
transform 1 0 5460 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_465
timestamp 1586547711
transform 1 0 5644 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1487
timestamp 1586547711
transform 1 0 5828 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1666
timestamp 1586547711
transform 1 0 6104 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1486
timestamp 1586547711
transform 1 0 6932 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL29440x8160
timestamp 1586547711
transform 1 0 6288 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1586547711
transform 1 0 6012 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _801_
timestamp 1586547711
transform 1 0 6380 0 1 2032
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1586
timestamp 1586547711
transform 1 0 7116 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_105
timestamp 1586547711
transform 1 0 7668 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1586547711
transform 1 0 7852 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL34500x8160
timestamp 1586547711
transform 1 0 7300 0 1 2032
box 0 -48 368 592
use sky130_fd_sc_hd__dfstp_4  _874_
timestamp 1586547711
transform 1 0 8036 0 1 2032
box 0 -48 2208 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1586547711
transform 1 0 10244 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_75
timestamp 1586547711
transform 1 0 10428 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_351
timestamp 1586547711
transform 1 0 10612 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1655
timestamp 1586547711
transform 1 0 10796 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL52900x8160
timestamp 1586547711
transform 1 0 10980 0 1 2032
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1093
timestamp 1586547711
transform 1 0 12360 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_347
timestamp 1586547711
transform 1 0 12544 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_77
timestamp 1586547711
transform 1 0 12728 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1586547711
transform 1 0 12912 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL55660x8160
timestamp 1586547711
transform 1 0 11532 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL59340x8160
timestamp 1586547711
transform 1 0 12268 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1586547711
transform 1 0 11624 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL56580x8160
timestamp 1586547711
transform 1 0 11716 0 1 2032
box 0 -48 552 592
use sky130_fd_sc_hd__dfrtp_4  _882_
timestamp 1586547711
transform 1 0 13096 0 1 2032
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_3  FILL74060x8160
timestamp 1586547711
transform 1 0 15212 0 1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_80
timestamp 1586547711
transform 1 0 15488 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_895
timestamp 1586547711
transform 1 0 15672 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1037
timestamp 1586547711
transform 1 0 15856 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL78200x8160
timestamp 1586547711
transform 1 0 16040 0 1 2032
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1038
timestamp 1586547711
transform 1 0 16500 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1036
timestamp 1586547711
transform 1 0 16684 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL80040x8160
timestamp 1586547711
transform 1 0 16408 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1021
timestamp 1586547711
transform 1 0 16868 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1025
timestamp 1586547711
transform 1 0 17052 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1586547711
transform 1 0 17236 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL84640x8160
timestamp 1586547711
transform 1 0 17328 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _571_ ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 17420 0 1 2032
box 0 -48 460 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1020
timestamp 1586547711
transform 1 0 17880 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_385
timestamp 1586547711
transform 1 0 18064 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_87
timestamp 1586547711
transform 1 0 18248 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1586547711
transform 1 0 18432 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__dfstp_4  _880_
timestamp 1586547711
transform 1 0 18616 0 1 2032
box 0 -48 2208 592
use sky130_fd_sc_hd__decap_3  FILL102120x8160
timestamp 1586547711
transform 1 0 20824 0 1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL107180x8160
timestamp 1586547711
transform 1 0 21836 0 1 2032
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1586547711
transform 1 0 21100 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_69
timestamp 1586547711
transform 1 0 21284 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_339
timestamp 1586547711
transform 1 0 21468 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1658
timestamp 1586547711
transform 1 0 21652 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILL110860x8160
timestamp 1586547711
transform 1 0 22572 0 1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1661
timestamp 1586547711
transform 1 0 22940 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_60
timestamp 1586547711
transform 1 0 23124 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp 1586547711
transform 1 0 23308 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1586547711
transform 1 0 22848 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _889_
timestamp 1586547711
transform 1 0 23492 0 1 2032
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1528
timestamp 1586547711
transform 1 0 25792 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_372
timestamp 1586547711
transform 1 0 25976 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_101
timestamp 1586547711
transform 1 0 26160 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _769_
timestamp 1586547711
transform 1 0 26344 0 1 2032
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILL126040x8160
timestamp 1586547711
transform 1 0 25608 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL142600x8160
timestamp 1586547711
transform 1 0 28920 0 1 2032
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1586547711
transform 1 0 28000 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_114
timestamp 1586547711
transform 1 0 28184 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_365
timestamp 1586547711
transform 1 0 28552 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1642
timestamp 1586547711
transform 1 0 28736 0 1 2032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL139840x8160
timestamp 1586547711
transform 1 0 28368 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1586547711
transform 1 0 28460 0 1 2032
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL136160x8160
timestamp 1586547711
transform 1 0 27632 0 1 2032
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL148120x8160
timestamp 1586547711
transform 1 0 30024 0 1 2032
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL153640x8160
timestamp 1586547711
transform 1 0 31128 0 1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1586547711
transform 1 0 31404 0 1 2032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1586547711
transform 1 0 400 0 -1 3120
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL1380x10880
timestamp 1586547711
transform 1 0 676 0 -1 3120
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL4600x10880
timestamp 1586547711
transform 1 0 1320 0 -1 3120
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL10120x10880
timestamp 1586547711
transform 1 0 2424 0 -1 3120
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_469
timestamp 1586547711
transform 1 0 952 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1493
timestamp 1586547711
transform 1 0 1136 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1477
timestamp 1586547711
transform 1 0 2240 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL8280x10880
timestamp 1586547711
transform 1 0 2056 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1476
timestamp 1586547711
transform 1 0 3344 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL13800x10880
timestamp 1586547711
transform 1 0 3160 0 -1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL15640x10880
timestamp 1586547711
transform 1 0 3528 0 -1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1586547711
transform 1 0 3252 0 -1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL21620x10880
timestamp 1586547711
transform 1 0 4724 0 -1 3120
box 0 -48 368 592
use sky130_fd_sc_hd__a21o_4  _751_ ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 3620 0 -1 3120
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1465
timestamp 1586547711
transform 1 0 5092 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _904_
timestamp 1586547711
transform 1 0 5460 0 -1 3120
box 0 -48 2116 592
use sky130_fd_sc_hd__fill_2  FILL24380x10880
timestamp 1586547711
transform 1 0 5276 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_371
timestamp 1586547711
transform 1 0 8036 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL37720x10880
timestamp 1586547711
transform 1 0 7944 0 -1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL41860x10880
timestamp 1586547711
transform 1 0 8772 0 -1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1586547711
transform 1 0 8864 0 -1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL35880x10880
timestamp 1586547711
transform 1 0 7576 0 -1 3120
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILL42780x10880
timestamp 1586547711
transform 1 0 8956 0 -1 3120
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILL39100x10880
timestamp 1586547711
transform 1 0 8220 0 -1 3120
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1519
timestamp 1586547711
transform 1 0 9324 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _884_
timestamp 1586547711
transform 1 0 9692 0 -1 3120
box 0 -48 2116 592
use sky130_fd_sc_hd__fill_2  FILL45540x10880
timestamp 1586547711
transform 1 0 9508 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL59800x10880
timestamp 1586547711
transform 1 0 12360 0 -1 3120
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_350
timestamp 1586547711
transform 1 0 11808 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_791
timestamp 1586547711
transform 1 0 11992 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_904
timestamp 1586547711
transform 1 0 12176 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _596_ ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 13096 0 -1 3120
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL70840x10880
timestamp 1586547711
transform 1 0 14568 0 -1 3120
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_902
timestamp 1586547711
transform 1 0 13740 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1586547711
transform 1 0 14476 0 -1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL67620x10880
timestamp 1586547711
transform 1 0 13924 0 -1 3120
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILL74520x10880
timestamp 1586547711
transform 1 0 15304 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _574_
timestamp 1586547711
transform 1 0 15488 0 -1 3120
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL78660x10880
timestamp 1586547711
transform 1 0 16132 0 -1 3120
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1094
timestamp 1586547711
transform 1 0 17880 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1031
timestamp 1586547711
transform 1 0 18064 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL86480x10880
timestamp 1586547711
transform 1 0 17696 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__and3_4  _575_ ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 16868 0 -1 3120
box 0 -48 828 592
use sky130_fd_sc_hd__decap_8  FILL98900x10880
timestamp 1586547711
transform 1 0 20180 0 -1 3120
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1092
timestamp 1586547711
transform 1 0 18248 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1022
timestamp 1586547711
transform 1 0 19260 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1651
timestamp 1586547711
transform 1 0 19444 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL97980x10880
timestamp 1586547711
transform 1 0 19996 0 -1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1586547711
transform 1 0 20088 0 -1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL96140x10880
timestamp 1586547711
transform 1 0 19628 0 -1 3120
box 0 -48 368 592
use sky130_fd_sc_hd__and3_4  _597_
timestamp 1586547711
transform 1 0 18432 0 -1 3120
box 0 -48 828 592
use sky130_fd_sc_hd__dfrtp_4  _886_
timestamp 1586547711
transform 1 0 21100 0 -1 3120
box 0 -48 2116 592
use sky130_fd_sc_hd__fill_2  FILL102580x10880
timestamp 1586547711
transform 1 0 20916 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL116380x10880
timestamp 1586547711
transform 1 0 23676 0 -1 3120
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL114080x10880
timestamp 1586547711
transform 1 0 23216 0 -1 3120
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_345
timestamp 1586547711
transform 1 0 23492 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1013
timestamp 1586547711
transform 1 0 24872 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_59
timestamp 1586547711
transform 1 0 25792 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL121900x10880
timestamp 1586547711
transform 1 0 24780 0 -1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL126040x10880
timestamp 1586547711
transform 1 0 25608 0 -1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1586547711
transform 1 0 25700 0 -1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL123280x10880
timestamp 1586547711
transform 1 0 25056 0 -1 3120
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL130640x10880
timestamp 1586547711
transform 1 0 26528 0 -1 3120
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_877
timestamp 1586547711
transform 1 0 25976 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1188
timestamp 1586547711
transform 1 0 26160 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_803
timestamp 1586547711
transform 1 0 26344 0 -1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL136160x10880
timestamp 1586547711
transform 1 0 27632 0 -1 3120
box 0 -48 368 592
use sky130_fd_sc_hd__dfstp_4  _871_
timestamp 1586547711
transform 1 0 28000 0 -1 3120
box 0 -48 2208 592
use sky130_fd_sc_hd__decap_12  FILL149040x10880
timestamp 1586547711
transform 1 0 30208 0 -1 3120
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1586547711
transform 1 0 31312 0 -1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1586547711
transform 1 0 31404 0 -1 3120
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1586547711
transform 1 0 400 0 1 3120
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_180
timestamp 1586547711
transform 1 0 1228 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_468
timestamp 1586547711
transform 1 0 1872 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_287
timestamp 1586547711
transform 1 0 2056 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL6900x13600
timestamp 1586547711
transform 1 0 1780 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL5060x13600
timestamp 1586547711
transform 1 0 1412 0 1 3120
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILL1380x13600
timestamp 1586547711
transform 1 0 676 0 1 3120
box 0 -48 552 592
use sky130_fd_sc_hd__a21o_4  _753_
timestamp 1586547711
transform 1 0 2240 0 1 3120
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_290
timestamp 1586547711
transform 1 0 3344 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1454
timestamp 1586547711
transform 1 0 3528 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1470
timestamp 1586547711
transform 1 0 3804 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1453
timestamp 1586547711
transform 1 0 3988 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_286
timestamp 1586547711
transform 1 0 4816 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL16560x13600
timestamp 1586547711
transform 1 0 3712 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _750_ ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 4172 0 1 3120
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_279
timestamp 1586547711
transform 1 0 5092 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_464
timestamp 1586547711
transform 1 0 5276 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1444
timestamp 1586547711
transform 1 0 5460 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL23000x13600
timestamp 1586547711
transform 1 0 5000 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1464
timestamp 1586547711
transform 1 0 5644 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1452
timestamp 1586547711
transform 1 0 5828 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1586547711
transform 1 0 6012 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _748_
timestamp 1586547711
transform 1 0 6104 0 1 3120
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_282
timestamp 1586547711
transform 1 0 6748 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_285
timestamp 1586547711
transform 1 0 6932 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL35420x13600
timestamp 1586547711
transform 1 0 7484 0 1 3120
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_795
timestamp 1586547711
transform 1 0 7116 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_800
timestamp 1586547711
transform 1 0 7300 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1527
timestamp 1586547711
transform 1 0 8772 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_370
timestamp 1586547711
transform 1 0 8956 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_104
timestamp 1586547711
transform 1 0 9140 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL40940x13600
timestamp 1586547711
transform 1 0 8588 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_903
timestamp 1586547711
transform 1 0 10612 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_782
timestamp 1586547711
transform 1 0 10796 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_76
timestamp 1586547711
transform 1 0 10980 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_348
timestamp 1586547711
transform 1 0 11164 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_73
timestamp 1586547711
transform 1 0 11440 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL54740x13600
timestamp 1586547711
transform 1 0 11348 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _768_
timestamp 1586547711
transform 1 0 9324 0 1 3120
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA_906
timestamp 1586547711
transform 1 0 13188 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_346
timestamp 1586547711
transform 1 0 13372 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_79
timestamp 1586547711
transform 1 0 13556 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1586547711
transform 1 0 11624 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _536_
timestamp 1586547711
transform 1 0 11716 0 1 3120
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILL63020x13600
timestamp 1586547711
transform 1 0 13004 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_894
timestamp 1586547711
transform 1 0 15028 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_905
timestamp 1586547711
transform 1 0 15212 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_893
timestamp 1586547711
transform 1 0 15856 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL76820x13600
timestamp 1586547711
transform 1 0 15764 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL74980x13600
timestamp 1586547711
transform 1 0 15396 0 1 3120
box 0 -48 368 592
use sky130_fd_sc_hd__o22a_4  _534_
timestamp 1586547711
transform 1 0 13740 0 1 3120
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA_896
timestamp 1586547711
transform 1 0 16040 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1041
timestamp 1586547711
transform 1 0 16684 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1040
timestamp 1586547711
transform 1 0 16868 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL80960x13600
timestamp 1586547711
transform 1 0 16592 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL79120x13600
timestamp 1586547711
transform 1 0 16224 0 1 3120
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1030
timestamp 1586547711
transform 1 0 17052 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_85
timestamp 1586547711
transform 1 0 17328 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1026
timestamp 1586547711
transform 1 0 17512 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1027
timestamp 1586547711
transform 1 0 17696 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_82
timestamp 1586547711
transform 1 0 17880 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1586547711
transform 1 0 17236 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__a211o_4  _598_ ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 18064 0 1 3120
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1096
timestamp 1586547711
transform 1 0 19352 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1500
timestamp 1586547711
transform 1 0 19720 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1028
timestamp 1586547711
transform 1 0 19904 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL95680x13600
timestamp 1586547711
transform 1 0 19536 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _760_
timestamp 1586547711
transform 1 0 20088 0 1 3120
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL107640x13600
timestamp 1586547711
transform 1 0 21928 0 1 3120
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_827
timestamp 1586547711
transform 1 0 20732 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_67
timestamp 1586547711
transform 1 0 21008 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_338
timestamp 1586547711
transform 1 0 21192 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_781
timestamp 1586547711
transform 1 0 21376 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_882
timestamp 1586547711
transform 1 0 21560 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_888
timestamp 1586547711
transform 1 0 21744 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL102580x13600
timestamp 1586547711
transform 1 0 20916 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1586547711
transform 1 0 22848 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL111320x13600
timestamp 1586547711
transform 1 0 22664 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_58
timestamp 1586547711
transform 1 0 23032 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_344
timestamp 1586547711
transform 1 0 23216 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL112700x13600
timestamp 1586547711
transform 1 0 22940 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_807
timestamp 1586547711
transform 1 0 23400 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_885
timestamp 1586547711
transform 1 0 23584 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_891
timestamp 1586547711
transform 1 0 23768 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL117760x13600
timestamp 1586547711
transform 1 0 23952 0 1 3120
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1033
timestamp 1586547711
transform 1 0 24320 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_100
timestamp 1586547711
transform 1 0 24504 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_62
timestamp 1586547711
transform 1 0 24688 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL132480x13600
timestamp 1586547711
transform 1 0 26896 0 1 3120
box 0 -48 552 592
use sky130_fd_sc_hd__a32oi_4  _619_ ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 24872 0 1 3120
box 0 -48 2024 592
use sky130_fd_sc_hd__diode_2  ANTENNA_377
timestamp 1586547711
transform 1 0 27540 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_376
timestamp 1586547711
transform 1 0 27724 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_99
timestamp 1586547711
transform 1 0 27908 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_98
timestamp 1586547711
transform 1 0 28092 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1586547711
transform 1 0 28276 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL135240x13600
timestamp 1586547711
transform 1 0 27448 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1586547711
transform 1 0 28460 0 1 3120
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _770_
timestamp 1586547711
transform 1 0 28552 0 1 3120
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_3  FILL153640x13600
timestamp 1586547711
transform 1 0 31128 0 1 3120
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL149960x13600
timestamp 1586547711
transform 1 0 30392 0 1 3120
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_808
timestamp 1586547711
transform 1 0 29840 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1521
timestamp 1586547711
transform 1 0 30024 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1529
timestamp 1586547711
transform 1 0 30208 0 1 3120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1586547711
transform 1 0 31404 0 1 3120
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1586547711
transform 1 0 400 0 1 4208
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1586547711
transform 1 0 400 0 -1 4208
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL1380x19040
timestamp 1586547711
transform 1 0 676 0 1 4208
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL5520x16320
timestamp 1586547711
transform 1 0 1504 0 -1 4208
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_291
timestamp 1586547711
transform 1 0 1412 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__conb_1  _830_
timestamp 1586547711
transform 1 0 1228 0 -1 4208
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILL1380x16320
timestamp 1586547711
transform 1 0 676 0 -1 4208
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL8740x19040
timestamp 1586547711
transform 1 0 2148 0 1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL10120x16320
timestamp 1586547711
transform 1 0 2424 0 -1 4208
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_470
timestamp 1586547711
transform 1 0 1596 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1447
timestamp 1586547711
transform 1 0 1780 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1483
timestamp 1586547711
transform 1 0 1964 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1446
timestamp 1586547711
transform 1 0 2240 0 -1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL14260x19040
timestamp 1586547711
transform 1 0 3252 0 1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL17940x16320
timestamp 1586547711
transform 1 0 3988 0 -1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_278
timestamp 1586547711
transform 1 0 4540 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1451
timestamp 1586547711
transform 1 0 4724 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL13800x16320
timestamp 1586547711
transform 1 0 3160 0 -1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1586547711
transform 1 0 3252 0 -1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL19780x19040
timestamp 1586547711
transform 1 0 4356 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _752_
timestamp 1586547711
transform 1 0 3344 0 -1 4208
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL23460x19040
timestamp 1586547711
transform 1 0 5092 0 1 4208
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1458
timestamp 1586547711
transform 1 0 4908 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_805
timestamp 1586547711
transform 1 0 5828 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _749_
timestamp 1586547711
transform 1 0 5092 0 -1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL28980x16320
timestamp 1586547711
transform 1 0 6196 0 -1 4208
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_289
timestamp 1586547711
transform 1 0 6748 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_796
timestamp 1586547711
transform 1 0 6932 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1586547711
transform 1 0 6012 0 1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _497_
timestamp 1586547711
transform 1 0 6104 0 1 4208
box 0 -48 644 592
use sky130_fd_sc_hd__or2_4  _495_
timestamp 1586547711
transform 1 0 6932 0 -1 4208
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL35880x16320
timestamp 1586547711
transform 1 0 7576 0 -1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL37260x19040
timestamp 1586547711
transform 1 0 7852 0 1 4208
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_281
timestamp 1586547711
transform 1 0 7300 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_764
timestamp 1586547711
transform 1 0 7484 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_785
timestamp 1586547711
transform 1 0 7668 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL33580x19040
timestamp 1586547711
transform 1 0 7116 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_788
timestamp 1586547711
transform 1 0 8680 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL40940x19040
timestamp 1586547711
transform 1 0 8588 0 1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1586547711
transform 1 0 8864 0 -1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL42780x16320
timestamp 1586547711
transform 1 0 8956 0 -1 4208
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL41400x16320
timestamp 1586547711
transform 1 0 8680 0 -1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _489_
timestamp 1586547711
transform 1 0 8864 0 1 4208
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL45540x16320
timestamp 1586547711
transform 1 0 9508 0 -1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_776
timestamp 1586547711
transform 1 0 9416 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_779
timestamp 1586547711
transform 1 0 9600 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_786
timestamp 1586547711
transform 1 0 9784 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_793
timestamp 1586547711
transform 1 0 9324 0 -1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL47840x19040
timestamp 1586547711
transform 1 0 9968 0 1 4208
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1586547711
transform 1 0 10520 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_111
timestamp 1586547711
transform 1 0 10704 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_367
timestamp 1586547711
transform 1 0 10888 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1643
timestamp 1586547711
transform 1 0 11072 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_907
timestamp 1586547711
transform 1 0 10796 0 -1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL54280x19040
timestamp 1586547711
transform 1 0 11256 0 1 4208
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL51060x16320
timestamp 1586547711
transform 1 0 10612 0 -1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _535_
timestamp 1586547711
transform 1 0 10980 0 -1 4208
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL56580x19040
timestamp 1586547711
transform 1 0 11716 0 1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL60260x16320
timestamp 1586547711
transform 1 0 12452 0 -1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_901
timestamp 1586547711
transform 1 0 13464 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_908
timestamp 1586547711
transform 1 0 12268 0 -1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL64860x19040
timestamp 1586547711
transform 1 0 13372 0 1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1586547711
transform 1 0 11624 0 1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL62100x19040
timestamp 1586547711
transform 1 0 12820 0 1 4208
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILL65780x16320
timestamp 1586547711
transform 1 0 13556 0 -1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _532_
timestamp 1586547711
transform 1 0 13648 0 1 4208
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_825
timestamp 1586547711
transform 1 0 14292 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_897
timestamp 1586547711
transform 1 0 14476 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_774
timestamp 1586547711
transform 1 0 13740 0 -1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1586547711
transform 1 0 14476 0 -1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL67620x16320
timestamp 1586547711
transform 1 0 13924 0 -1 4208
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILL73600x16320
timestamp 1586547711
transform 1 0 15120 0 -1 4208
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1114
timestamp 1586547711
transform 1 0 14660 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1012
timestamp 1586547711
transform 1 0 14844 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_875
timestamp 1586547711
transform 1 0 15028 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_103
timestamp 1586547711
transform 1 0 15212 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _533_
timestamp 1586547711
transform 1 0 14568 0 -1 4208
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_910
timestamp 1586547711
transform 1 0 15396 0 -1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1032
timestamp 1586547711
transform 1 0 15580 0 -1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL76820x16320
timestamp 1586547711
transform 1 0 15764 0 -1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _531_
timestamp 1586547711
transform 1 0 15856 0 -1 4208
box 0 -48 460 592
use sky130_fd_sc_hd__and3_4  _606_
timestamp 1586547711
transform 1 0 15396 0 1 4208
box 0 -48 828 592
use sky130_fd_sc_hd__decap_8  FILL79580x16320
timestamp 1586547711
transform 1 0 16316 0 -1 4208
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_65
timestamp 1586547711
transform 1 0 16224 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1115
timestamp 1586547711
transform 1 0 16408 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1116
timestamp 1586547711
transform 1 0 16592 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1117
timestamp 1586547711
transform 1 0 16776 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL82800x19040
timestamp 1586547711
transform 1 0 16960 0 1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_874
timestamp 1586547711
transform 1 0 17052 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_871
timestamp 1586547711
transform 1 0 17328 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_71
timestamp 1586547711
transform 1 0 17512 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_68
timestamp 1586547711
transform 1 0 17696 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1586547711
transform 1 0 17236 0 1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL83260x16320
timestamp 1586547711
transform 1 0 17052 0 -1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _595_
timestamp 1586547711
transform 1 0 17880 0 1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__a211o_4  _576_
timestamp 1586547711
transform 1 0 17236 0 -1 4208
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_8  FILL93380x16320
timestamp 1586547711
transform 1 0 19076 0 -1 4208
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_898
timestamp 1586547711
transform 1 0 18984 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1035
timestamp 1586547711
transform 1 0 19168 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_899
timestamp 1586547711
transform 1 0 18524 0 -1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1091
timestamp 1586547711
transform 1 0 18708 0 -1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1097
timestamp 1586547711
transform 1 0 18892 0 -1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL94760x19040
timestamp 1586547711
transform 1 0 19352 0 1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL97060x16320
timestamp 1586547711
transform 1 0 19812 0 -1 4208
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL98900x16320
timestamp 1586547711
transform 1 0 20180 0 -1 4208
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1586547711
transform 1 0 20088 0 -1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL100280x19040
timestamp 1586547711
transform 1 0 20456 0 1 4208
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1586547711
transform 1 0 21376 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL102580x16320
timestamp 1586547711
transform 1 0 20916 0 -1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL103960x19040
timestamp 1586547711
transform 1 0 21192 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL108560x19040
timestamp 1586547711
transform 1 0 22112 0 1 4208
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL109480x16320
timestamp 1586547711
transform 1 0 22296 0 -1 4208
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_72
timestamp 1586547711
transform 1 0 21560 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_337
timestamp 1586547711
transform 1 0 21744 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1657
timestamp 1586547711
transform 1 0 21928 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _526_
timestamp 1586547711
transform 1 0 21008 0 -1 4208
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL112700x19040
timestamp 1586547711
transform 1 0 22940 0 1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL120980x19040
timestamp 1586547711
transform 1 0 24596 0 1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_879
timestamp 1586547711
transform 1 0 24228 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_880
timestamp 1586547711
transform 1 0 24412 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1586547711
transform 1 0 22848 0 1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL119600x16320
timestamp 1586547711
transform 1 0 24320 0 -1 4208
box 0 -48 552 592
use sky130_fd_sc_hd__o22a_4  _529_
timestamp 1586547711
transform 1 0 23032 0 -1 4208
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILL118220x19040
timestamp 1586547711
transform 1 0 24044 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL126500x19040
timestamp 1586547711
transform 1 0 25700 0 1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL130180x16320
timestamp 1586547711
transform 1 0 26436 0 -1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL132020x19040
timestamp 1586547711
transform 1 0 26804 0 1 4208
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_876
timestamp 1586547711
transform 1 0 24872 0 -1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1151
timestamp 1586547711
transform 1 0 25056 0 -1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL126040x16320
timestamp 1586547711
transform 1 0 25608 0 -1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1586547711
transform 1 0 25700 0 -1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL124200x16320
timestamp 1586547711
transform 1 0 25240 0 -1 4208
box 0 -48 368 592
use sky130_fd_sc_hd__and2_4  _633_
timestamp 1586547711
transform 1 0 25792 0 -1 4208
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL135240x19040
timestamp 1586547711
transform 1 0 27448 0 1 4208
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1192
timestamp 1586547711
transform 1 0 27080 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1524
timestamp 1586547711
transform 1 0 27264 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL135700x16320
timestamp 1586547711
transform 1 0 27540 0 -1 4208
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILL138920x19040
timestamp 1586547711
transform 1 0 28184 0 1 4208
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1586547711
transform 1 0 28552 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_120
timestamp 1586547711
transform 1 0 28736 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_361
timestamp 1586547711
transform 1 0 28920 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1640
timestamp 1586547711
transform 1 0 29104 0 1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1647
timestamp 1586547711
transform 1 0 28184 0 -1 4208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL138460x16320
timestamp 1586547711
transform 1 0 28092 0 -1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1586547711
transform 1 0 28460 0 1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__dfstp_4  _876_
timestamp 1586547711
transform 1 0 28368 0 -1 4208
box 0 -48 2208 592
use sky130_fd_sc_hd__decap_12  FILL144440x19040
timestamp 1586547711
transform 1 0 29288 0 1 4208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL153640x19040
timestamp 1586547711
transform 1 0 31128 0 1 4208
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL149960x19040
timestamp 1586547711
transform 1 0 30392 0 1 4208
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL150880x16320
timestamp 1586547711
transform 1 0 30576 0 -1 4208
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1586547711
transform 1 0 31312 0 -1 4208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1586547711
transform 1 0 31404 0 1 4208
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1586547711
transform 1 0 31404 0 -1 4208
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1586547711
transform 1 0 400 0 -1 5296
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL10580x21760
timestamp 1586547711
transform 1 0 2516 0 -1 5296
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_471
timestamp 1586547711
transform 1 0 676 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_172
timestamp 1586547711
transform 1 0 860 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1497
timestamp 1586547711
transform 1 0 1044 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL4140x21760
timestamp 1586547711
transform 1 0 1228 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _755_
timestamp 1586547711
transform 1 0 1412 0 -1 5296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL14720x21760
timestamp 1586547711
transform 1 0 3344 0 -1 5296
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1485
timestamp 1586547711
transform 1 0 3620 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1665
timestamp 1586547711
transform 1 0 3804 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_760
timestamp 1586547711
transform 1 0 3988 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1443
timestamp 1586547711
transform 1 0 4172 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1586547711
transform 1 0 3252 0 -1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL19780x21760
timestamp 1586547711
transform 1 0 4356 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _746_
timestamp 1586547711
transform 1 0 4540 0 -1 5296
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL23920x21760
timestamp 1586547711
transform 1 0 5184 0 -1 5296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL33120x21760
timestamp 1586547711
transform 1 0 7024 0 -1 5296
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL29440x21760
timestamp 1586547711
transform 1 0 6288 0 -1 5296
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL37720x21760
timestamp 1586547711
transform 1 0 7944 0 -1 5296
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1586547711
transform 1 0 8864 0 -1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL41400x21760
timestamp 1586547711
transform 1 0 8680 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _492_
timestamp 1586547711
transform 1 0 8956 0 -1 5296
box 0 -48 552 592
use sky130_fd_sc_hd__or2_4  _491_
timestamp 1586547711
transform 1 0 7300 0 -1 5296
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_368
timestamp 1586547711
transform 1 0 9508 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_777
timestamp 1586547711
transform 1 0 9692 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1526
timestamp 1586547711
transform 1 0 9876 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL50140x21760
timestamp 1586547711
transform 1 0 10428 0 -1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL48300x21760
timestamp 1586547711
transform 1 0 10060 0 -1 5296
box 0 -48 368 592
use sky130_fd_sc_hd__dfstp_4  _872_
timestamp 1586547711
transform 1 0 10520 0 -1 5296
box 0 -48 2208 592
use sky130_fd_sc_hd__decap_12  FILL61640x21760
timestamp 1586547711
transform 1 0 12728 0 -1 5296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL70840x21760
timestamp 1586547711
transform 1 0 14568 0 -1 5296
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL69920x21760
timestamp 1586547711
transform 1 0 14384 0 -1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL74520x21760
timestamp 1586547711
transform 1 0 15304 0 -1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1586547711
transform 1 0 14476 0 -1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL67160x21760
timestamp 1586547711
transform 1 0 13832 0 -1 5296
box 0 -48 552 592
use sky130_fd_sc_hd__o32a_4  _607_ ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 15396 0 -1 5296
box 0 -48 1656 592
use sky130_fd_sc_hd__decap_8  FILL83260x21760
timestamp 1586547711
transform 1 0 17052 0 -1 5296
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL86940x21760
timestamp 1586547711
transform 1 0 17788 0 -1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__a21o_4  _573_
timestamp 1586547711
transform 1 0 17880 0 -1 5296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL92920x21760
timestamp 1586547711
transform 1 0 18984 0 -1 5296
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1586547711
transform 1 0 20088 0 -1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL98900x21760
timestamp 1586547711
transform 1 0 20180 0 -1 5296
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_336
timestamp 1586547711
transform 1 0 20824 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_773
timestamp 1586547711
transform 1 0 21008 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_881
timestamp 1586547711
transform 1 0 21192 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL101660x21760
timestamp 1586547711
transform 1 0 20732 0 -1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _885_
timestamp 1586547711
transform 1 0 21376 0 -1 5296
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_8  FILL115460x21760
timestamp 1586547711
transform 1 0 23492 0 -1 5296
box 0 -48 736 592
use sky130_fd_sc_hd__buf_4  _523_
timestamp 1586547711
transform 1 0 24228 0 -1 5296
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL126960x21760
timestamp 1586547711
transform 1 0 25792 0 -1 5296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL121900x21760
timestamp 1586547711
transform 1 0 24780 0 -1 5296
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1586547711
transform 1 0 25700 0 -1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL125580x21760
timestamp 1586547711
transform 1 0 25516 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL132480x21760
timestamp 1586547711
transform 1 0 26896 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1196
timestamp 1586547711
transform 1 0 27632 0 -1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL137080x21760
timestamp 1586547711
transform 1 0 27816 0 -1 5296
box 0 -48 552 592
use sky130_fd_sc_hd__buf_4  _765_
timestamp 1586547711
transform 1 0 27080 0 -1 5296
box 0 -48 552 592
use sky130_fd_sc_hd__dfstp_4  _869_
timestamp 1586547711
transform 1 0 28368 0 -1 5296
box 0 -48 2208 592
use sky130_fd_sc_hd__decap_8  FILL150880x21760
timestamp 1586547711
transform 1 0 30576 0 -1 5296
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1586547711
transform 1 0 31312 0 -1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1586547711
transform 1 0 31404 0 -1 5296
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1586547711
transform 1 0 400 0 1 5296
box 0 -48 276 592
use sky130_fd_sc_hd__dfrtp_4  _907_
timestamp 1586547711
transform 1 0 676 0 1 5296
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA_294
timestamp 1586547711
transform 1 0 2792 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1455
timestamp 1586547711
transform 1 0 2976 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1459
timestamp 1586547711
transform 1 0 3252 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_463
timestamp 1586547711
transform 1 0 3436 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_280
timestamp 1586547711
transform 1 0 3620 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_462
timestamp 1586547711
transform 1 0 3804 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL13800x24480
timestamp 1586547711
transform 1 0 3160 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__a21o_4  _747_
timestamp 1586547711
transform 1 0 3988 0 1 5296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL23460x24480
timestamp 1586547711
transform 1 0 5092 0 1 5296
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_794
timestamp 1586547711
transform 1 0 6564 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_765
timestamp 1586547711
transform 1 0 6748 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_775
timestamp 1586547711
transform 1 0 7024 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL30360x24480
timestamp 1586547711
transform 1 0 6472 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL32660x24480
timestamp 1586547711
transform 1 0 6932 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1586547711
transform 1 0 6012 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL28520x24480
timestamp 1586547711
transform 1 0 6104 0 1 5296
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL27140x24480
timestamp 1586547711
transform 1 0 5828 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _488_
timestamp 1586547711
transform 1 0 7208 0 1 5296
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_277
timestamp 1586547711
transform 1 0 7852 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_763
timestamp 1586547711
transform 1 0 8036 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1644
timestamp 1586547711
transform 1 0 8312 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL39100x24480
timestamp 1586547711
transform 1 0 8220 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1518
timestamp 1586547711
transform 1 0 8496 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_369
timestamp 1586547711
transform 1 0 8680 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_108
timestamp 1586547711
transform 1 0 8864 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1586547711
transform 1 0 9048 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_107
timestamp 1586547711
transform 1 0 9232 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1517
timestamp 1586547711
transform 1 0 11072 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_366
timestamp 1586547711
transform 1 0 11256 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_110
timestamp 1586547711
transform 1 0 11440 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL51520x24480
timestamp 1586547711
transform 1 0 10704 0 1 5296
box 0 -48 368 592
use sky130_fd_sc_hd__o22a_4  _767_
timestamp 1586547711
transform 1 0 9416 0 1 5296
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA_767
timestamp 1586547711
transform 1 0 13188 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_769
timestamp 1586547711
transform 1 0 13372 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1113
timestamp 1586547711
transform 1 0 13648 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL65780x24480
timestamp 1586547711
transform 1 0 13556 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1586547711
transform 1 0 11624 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _766_
timestamp 1586547711
transform 1 0 11716 0 1 5296
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILL63020x24480
timestamp 1586547711
transform 1 0 13004 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILL72220x24480
timestamp 1586547711
transform 1 0 14844 0 1 5296
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_74
timestamp 1586547711
transform 1 0 14476 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_900
timestamp 1586547711
transform 1 0 14660 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1029
timestamp 1586547711
transform 1 0 15120 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1008
timestamp 1586547711
transform 1 0 15764 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _572_
timestamp 1586547711
transform 1 0 15304 0 1 5296
box 0 -48 460 592
use sky130_fd_sc_hd__and2_4  _605_
timestamp 1586547711
transform 1 0 13832 0 1 5296
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL79580x24480
timestamp 1586547711
transform 1 0 16316 0 1 5296
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL84640x24480
timestamp 1586547711
transform 1 0 17328 0 1 5296
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1018
timestamp 1586547711
transform 1 0 15948 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1019
timestamp 1586547711
transform 1 0 16132 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1586547711
transform 1 0 17236 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL83260x24480
timestamp 1586547711
transform 1 0 17052 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL88320x24480
timestamp 1586547711
transform 1 0 18064 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_867
timestamp 1586547711
transform 1 0 18248 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_869
timestamp 1586547711
transform 1 0 18432 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL91080x24480
timestamp 1586547711
transform 1 0 18616 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _521_
timestamp 1586547711
transform 1 0 18708 0 1 5296
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_870
timestamp 1586547711
transform 1 0 19260 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_872
timestamp 1586547711
transform 1 0 19444 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL96140x24480
timestamp 1586547711
transform 1 0 19628 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1659
timestamp 1586547711
transform 1 0 19812 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_341
timestamp 1586547711
transform 1 0 19996 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1586547711
transform 1 0 20180 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_66
timestamp 1586547711
transform 1 0 20364 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_70
timestamp 1586547711
transform 1 0 20640 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_887
timestamp 1586547711
transform 1 0 22112 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL100740x24480
timestamp 1586547711
transform 1 0 20548 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL109480x24480
timestamp 1586547711
transform 1 0 22296 0 1 5296
box 0 -48 552 592
use sky130_fd_sc_hd__o22a_4  _525_
timestamp 1586547711
transform 1 0 20824 0 1 5296
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_8  FILL112700x24480
timestamp 1586547711
transform 1 0 22940 0 1 5296
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_878
timestamp 1586547711
transform 1 0 23768 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_628
timestamp 1586547711
transform 1 0 24596 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL116380x24480
timestamp 1586547711
transform 1 0 23676 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1586547711
transform 1 0 22848 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _522_
timestamp 1586547711
transform 1 0 23952 0 1 5296
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_873
timestamp 1586547711
transform 1 0 24780 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1034
timestamp 1586547711
transform 1 0 26160 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1182
timestamp 1586547711
transform 1 0 26344 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1190
timestamp 1586547711
transform 1 0 26712 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL125580x24480
timestamp 1586547711
transform 1 0 25516 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL122820x24480
timestamp 1586547711
transform 1 0 24964 0 1 5296
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILL130640x24480
timestamp 1586547711
transform 1 0 26528 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _632_
timestamp 1586547711
transform 1 0 25608 0 1 5296
box 0 -48 552 592
use sky130_fd_sc_hd__buf_4  _634_
timestamp 1586547711
transform 1 0 26896 0 1 5296
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_97
timestamp 1586547711
transform 1 0 27448 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1014
timestamp 1586547711
transform 1 0 27632 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1183
timestamp 1586547711
transform 1 0 27816 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1189
timestamp 1586547711
transform 1 0 28000 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1191
timestamp 1586547711
transform 1 0 28184 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1510
timestamp 1586547711
transform 1 0 29104 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL139840x24480
timestamp 1586547711
transform 1 0 28368 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1586547711
transform 1 0 28460 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _764_
timestamp 1586547711
transform 1 0 28552 0 1 5296
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL145360x24480
timestamp 1586547711
transform 1 0 29472 0 1 5296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL150880x24480
timestamp 1586547711
transform 1 0 30576 0 1 5296
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1516
timestamp 1586547711
transform 1 0 29288 0 1 5296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL154560x24480
timestamp 1586547711
transform 1 0 31312 0 1 5296
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1586547711
transform 1 0 31404 0 1 5296
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1586547711
transform 1 0 400 0 -1 6384
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_296
timestamp 1586547711
transform 1 0 676 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1669
timestamp 1586547711
transform 1 0 1136 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1482
timestamp 1586547711
transform 1 0 2516 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__conb_1  _833_
timestamp 1586547711
transform 1 0 860 0 -1 6384
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILL4600x27200
timestamp 1586547711
transform 1 0 1320 0 -1 6384
box 0 -48 552 592
use sky130_fd_sc_hd__and2_4  _754_
timestamp 1586547711
transform 1 0 1872 0 -1 6384
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  FILL14720x27200
timestamp 1586547711
transform 1 0 3344 0 -1 6384
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1586547711
transform 1 0 3252 0 -1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL11500x27200
timestamp 1586547711
transform 1 0 2700 0 -1 6384
box 0 -48 552 592
use sky130_fd_sc_hd__dfrtp_4  _903_
timestamp 1586547711
transform 1 0 3620 0 -1 6384
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_3  FILL30360x27200
timestamp 1586547711
transform 1 0 6472 0 -1 6384
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL26680x27200
timestamp 1586547711
transform 1 0 5736 0 -1 6384
box 0 -48 736 592
use sky130_fd_sc_hd__buf_4  _494_
timestamp 1586547711
transform 1 0 6748 0 -1 6384
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILL40940x27200
timestamp 1586547711
transform 1 0 8588 0 -1 6384
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL37260x27200
timestamp 1586547711
transform 1 0 7852 0 -1 6384
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1558
timestamp 1586547711
transform 1 0 7668 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL42780x27200
timestamp 1586547711
transform 1 0 8956 0 -1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1586547711
transform 1 0 8864 0 -1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL34500x27200
timestamp 1586547711
transform 1 0 7300 0 -1 6384
box 0 -48 368 592
use sky130_fd_sc_hd__dfstp_4  _873_
timestamp 1586547711
transform 1 0 9048 0 -1 6384
box 0 -48 2208 592
use sky130_fd_sc_hd__decap_4  FILL54280x27200
timestamp 1586547711
transform 1 0 11256 0 -1 6384
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL58420x27200
timestamp 1586547711
transform 1 0 12084 0 -1 6384
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_928
timestamp 1586547711
transform 1 0 11716 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1525
timestamp 1586547711
transform 1 0 11900 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL56120x27200
timestamp 1586547711
transform 1 0 11624 0 -1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _486_
timestamp 1586547711
transform 1 0 13188 0 -1 6384
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL66700x27200
timestamp 1586547711
transform 1 0 13740 0 -1 6384
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1089
timestamp 1586547711
transform 1 0 15120 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL76360x27200
timestamp 1586547711
transform 1 0 15672 0 -1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1586547711
transform 1 0 14476 0 -1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL74520x27200
timestamp 1586547711
transform 1 0 15304 0 -1 6384
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILL70840x27200
timestamp 1586547711
transform 1 0 14568 0 -1 6384
box 0 -48 552 592
use sky130_fd_sc_hd__buf_4  _570_
timestamp 1586547711
transform 1 0 15764 0 -1 6384
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL79580x27200
timestamp 1586547711
transform 1 0 16316 0 -1 6384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL85100x27200
timestamp 1586547711
transform 1 0 17420 0 -1 6384
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILL91540x27200
timestamp 1586547711
transform 1 0 18708 0 -1 6384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL97060x27200
timestamp 1586547711
transform 1 0 19812 0 -1 6384
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL88780x27200
timestamp 1586547711
transform 1 0 18156 0 -1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1586547711
transform 1 0 20088 0 -1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__dfstp_4  _887_
timestamp 1586547711
transform 1 0 20180 0 -1 6384
box 0 -48 2208 592
use sky130_fd_sc_hd__inv_4  _520_
timestamp 1586547711
transform 1 0 18248 0 -1 6384
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL109940x27200
timestamp 1586547711
transform 1 0 22388 0 -1 6384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL120060x27200
timestamp 1586547711
transform 1 0 24412 0 -1 6384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL115460x27200
timestamp 1586547711
transform 1 0 23492 0 -1 6384
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1641
timestamp 1586547711
transform 1 0 24228 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL126960x27200
timestamp 1586547711
transform 1 0 25792 0 -1 6384
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1586547711
transform 1 0 25700 0 -1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL132480x27200
timestamp 1586547711
transform 1 0 26896 0 -1 6384
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL125580x27200
timestamp 1586547711
transform 1 0 25516 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_364
timestamp 1586547711
transform 1 0 28828 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_821
timestamp 1586547711
transform 1 0 29012 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL134320x27200
timestamp 1586547711
transform 1 0 27264 0 -1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__o22ai_4  _635_ ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 27356 0 -1 6384
box 0 -48 1472 592
use sky130_fd_sc_hd__decap_12  FILL144900x27200
timestamp 1586547711
transform 1 0 29380 0 -1 6384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL150420x27200
timestamp 1586547711
transform 1 0 30484 0 -1 6384
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1130
timestamp 1586547711
transform 1 0 29196 0 -1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL154100x27200
timestamp 1586547711
transform 1 0 31220 0 -1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1586547711
transform 1 0 31312 0 -1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1586547711
transform 1 0 31404 0 -1 6384
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL1380x29920
timestamp 1586547711
transform 1 0 676 0 1 6384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1586547711
transform 1 0 400 0 1 6384
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL10580x29920
timestamp 1586547711
transform 1 0 2516 0 1 6384
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL6900x29920
timestamp 1586547711
transform 1 0 1780 0 1 6384
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1442
timestamp 1586547711
transform 1 0 2792 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1435
timestamp 1586547711
transform 1 0 3528 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1439
timestamp 1586547711
transform 1 0 3712 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1450
timestamp 1586547711
transform 1 0 3896 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1585
timestamp 1586547711
transform 1 0 4264 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL18400x29920
timestamp 1586547711
transform 1 0 4080 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _744_
timestamp 1586547711
transform 1 0 2976 0 1 6384
box 0 -48 552 592
use sky130_fd_sc_hd__buf_4  _800_
timestamp 1586547711
transform 1 0 4448 0 1 6384
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILL32200x29920
timestamp 1586547711
transform 1 0 6840 0 1 6384
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL28520x29920
timestamp 1586547711
transform 1 0 6104 0 1 6384
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1484
timestamp 1586547711
transform 1 0 5000 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_293
timestamp 1586547711
transform 1 0 5276 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_797
timestamp 1586547711
transform 1 0 5460 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_810
timestamp 1586547711
transform 1 0 5644 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL23920x29920
timestamp 1586547711
transform 1 0 5184 0 1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1586547711
transform 1 0 6012 0 1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL27140x29920
timestamp 1586547711
transform 1 0 5828 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL42780x29920
timestamp 1586547711
transform 1 0 8956 0 1 6384
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1566
timestamp 1586547711
transform 1 0 7116 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_354
timestamp 1586547711
transform 1 0 7300 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_128
timestamp 1586547711
transform 1 0 7484 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _779_
timestamp 1586547711
transform 1 0 7668 0 1 6384
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL48300x29920
timestamp 1586547711
transform 1 0 10060 0 1 6384
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_766
timestamp 1586547711
transform 1 0 11256 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_762
timestamp 1586547711
transform 1 0 11440 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL53820x29920
timestamp 1586547711
transform 1 0 11164 0 1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_326
timestamp 1586547711
transform 1 0 12360 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_756
timestamp 1586547711
transform 1 0 12544 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_761
timestamp 1586547711
transform 1 0 12728 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_768
timestamp 1586547711
transform 1 0 13648 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1586547711
transform 1 0 11624 0 1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL62560x29920
timestamp 1586547711
transform 1 0 12912 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _541_
timestamp 1586547711
transform 1 0 13096 0 1 6384
box 0 -48 552 592
use sky130_fd_sc_hd__or2_4  _485_
timestamp 1586547711
transform 1 0 11716 0 1 6384
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_924
timestamp 1586547711
transform 1 0 13832 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1015
timestamp 1586547711
transform 1 0 14476 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1010
timestamp 1586547711
transform 1 0 14660 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_109
timestamp 1586547711
transform 1 0 14844 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_106
timestamp 1586547711
transform 1 0 15764 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL69920x29920
timestamp 1586547711
transform 1 0 14384 0 1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL73140x29920
timestamp 1586547711
transform 1 0 15028 0 1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL68080x29920
timestamp 1586547711
transform 1 0 14016 0 1 6384
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _594_
timestamp 1586547711
transform 1 0 15120 0 1 6384
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL78660x29920
timestamp 1586547711
transform 1 0 16132 0 1 6384
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1011
timestamp 1586547711
transform 1 0 15948 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_997
timestamp 1586547711
transform 1 0 17972 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL87400x29920
timestamp 1586547711
transform 1 0 17880 0 1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1586547711
transform 1 0 17236 0 1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL84640x29920
timestamp 1586547711
transform 1 0 17328 0 1 6384
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1090
timestamp 1586547711
transform 1 0 18156 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1098
timestamp 1586547711
transform 1 0 18340 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1099
timestamp 1586547711
transform 1 0 18524 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_886
timestamp 1586547711
transform 1 0 18800 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL91540x29920
timestamp 1586547711
transform 1 0 18708 0 1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _524_
timestamp 1586547711
transform 1 0 18984 0 1 6384
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_868
timestamp 1586547711
transform 1 0 19536 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_883
timestamp 1586547711
transform 1 0 19720 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_340
timestamp 1586547711
transform 1 0 19904 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_64
timestamp 1586547711
transform 1 0 20088 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _527_
timestamp 1586547711
transform 1 0 20272 0 1 6384
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL105800x29920
timestamp 1586547711
transform 1 0 21560 0 1 6384
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1549
timestamp 1586547711
transform 1 0 23308 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1555
timestamp 1586547711
transform 1 0 23492 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_117
timestamp 1586547711
transform 1 0 23860 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1586547711
transform 1 0 24044 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1586547711
transform 1 0 22848 0 1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL112700x29920
timestamp 1586547711
transform 1 0 22940 0 1 6384
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL111320x29920
timestamp 1586547711
transform 1 0 22664 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL116380x29920
timestamp 1586547711
transform 1 0 23676 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__dfstp_4  _870_
timestamp 1586547711
transform 1 0 24228 0 1 6384
box 0 -48 2208 592
use sky130_fd_sc_hd__diode_2  ANTENNA_630
timestamp 1586547711
transform 1 0 26620 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1187
timestamp 1586547711
transform 1 0 26804 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL130180x29920
timestamp 1586547711
transform 1 0 26436 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1509
timestamp 1586547711
transform 1 0 26988 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1550
timestamp 1586547711
transform 1 0 27356 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1128
timestamp 1586547711
transform 1 0 27540 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_813
timestamp 1586547711
transform 1 0 27724 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_360
timestamp 1586547711
transform 1 0 27908 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL133860x29920
timestamp 1586547711
transform 1 0 27172 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_119
timestamp 1586547711
transform 1 0 28092 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_113
timestamp 1586547711
transform 1 0 28276 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1586547711
transform 1 0 28460 0 1 6384
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _784_
timestamp 1586547711
transform 1 0 28552 0 1 6384
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL148120x29920
timestamp 1586547711
transform 1 0 30024 0 1 6384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL153640x29920
timestamp 1586547711
transform 1 0 31128 0 1 6384
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1552
timestamp 1586547711
transform 1 0 29840 0 1 6384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1586547711
transform 1 0 31404 0 1 6384
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL1380x32640
timestamp 1586547711
transform 1 0 676 0 -1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL6900x32640
timestamp 1586547711
transform 1 0 1780 0 -1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1586547711
transform 1 0 400 0 -1 7472
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL18400x32640
timestamp 1586547711
transform 1 0 4080 0 -1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1586547711
transform 1 0 3252 0 -1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL12420x32640
timestamp 1586547711
transform 1 0 2884 0 -1 7472
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL14720x32640
timestamp 1586547711
transform 1 0 3344 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _745_
timestamp 1586547711
transform 1 0 3528 0 -1 7472
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL27600x32640
timestamp 1586547711
transform 1 0 5920 0 -1 7472
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_778
timestamp 1586547711
transform 1 0 6840 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_132
timestamp 1586547711
transform 1 0 7024 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL23920x32640
timestamp 1586547711
transform 1 0 5184 0 -1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL31280x32640
timestamp 1586547711
transform 1 0 6656 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _499_
timestamp 1586547711
transform 1 0 5276 0 -1 7472
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL42780x32640
timestamp 1586547711
transform 1 0 8956 0 -1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL40940x32640
timestamp 1586547711
transform 1 0 8588 0 -1 7472
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL37260x32640
timestamp 1586547711
transform 1 0 7852 0 -1 7472
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_403
timestamp 1586547711
transform 1 0 7208 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1635
timestamp 1586547711
transform 1 0 7392 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_787
timestamp 1586547711
transform 1 0 7668 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL35880x32640
timestamp 1586547711
transform 1 0 7576 0 -1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1586547711
transform 1 0 8864 0 -1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL48300x32640
timestamp 1586547711
transform 1 0 10060 0 -1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL53820x32640
timestamp 1586547711
transform 1 0 11164 0 -1 7472
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILL60260x32640
timestamp 1586547711
transform 1 0 12452 0 -1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL65780x32640
timestamp 1586547711
transform 1 0 13556 0 -1 7472
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL57500x32640
timestamp 1586547711
transform 1 0 11900 0 -1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _484_
timestamp 1586547711
transform 1 0 11992 0 -1 7472
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL75440x32640
timestamp 1586547711
transform 1 0 15488 0 -1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL70840x32640
timestamp 1586547711
transform 1 0 14568 0 -1 7472
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1586547711
transform 1 0 14476 0 -1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL69460x32640
timestamp 1586547711
transform 1 0 14292 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _568_
timestamp 1586547711
transform 1 0 14844 0 -1 7472
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL80960x32640
timestamp 1586547711
transform 1 0 16592 0 -1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL86480x32640
timestamp 1586547711
transform 1 0 17696 0 -1 7472
box 0 -48 276 592
use sky130_fd_sc_hd__and3_4  _599_
timestamp 1586547711
transform 1 0 17972 0 -1 7472
box 0 -48 828 592
use sky130_fd_sc_hd__decap_12  FILL92000x32640
timestamp 1586547711
transform 1 0 18800 0 -1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_790
timestamp 1586547711
transform 1 0 20272 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL98900x32640
timestamp 1586547711
transform 1 0 20180 0 -1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1586547711
transform 1 0 20088 0 -1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL97520x32640
timestamp 1586547711
transform 1 0 19904 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL101200x32640
timestamp 1586547711
transform 1 0 20640 0 -1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL106720x32640
timestamp 1586547711
transform 1 0 21744 0 -1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_889
timestamp 1586547711
transform 1 0 20456 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1563
timestamp 1586547711
transform 1 0 22940 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_363
timestamp 1586547711
transform 1 0 24228 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1003
timestamp 1586547711
transform 1 0 24412 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1083
timestamp 1586547711
transform 1 0 24596 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL112240x32640
timestamp 1586547711
transform 1 0 22848 0 -1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL117300x32640
timestamp 1586547711
transform 1 0 23860 0 -1 7472
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL113620x32640
timestamp 1586547711
transform 1 0 23124 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _775_
timestamp 1586547711
transform 1 0 23308 0 -1 7472
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL122820x32640
timestamp 1586547711
transform 1 0 24964 0 -1 7472
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL126960x32640
timestamp 1586547711
transform 1 0 25792 0 -1 7472
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1129
timestamp 1586547711
transform 1 0 24780 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL130640x32640
timestamp 1586547711
transform 1 0 26528 0 -1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1586547711
transform 1 0 25700 0 -1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _763_
timestamp 1586547711
transform 1 0 26620 0 -1 7472
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL134320x32640
timestamp 1586547711
transform 1 0 27264 0 -1 7472
box 0 -48 736 592
use sky130_fd_sc_hd__o22a_4  _782_
timestamp 1586547711
transform 1 0 28184 0 -1 7472
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILL138000x32640
timestamp 1586547711
transform 1 0 28000 0 -1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL145360x32640
timestamp 1586547711
transform 1 0 29472 0 -1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL150880x32640
timestamp 1586547711
transform 1 0 30576 0 -1 7472
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1586547711
transform 1 0 31312 0 -1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1586547711
transform 1 0 31404 0 -1 7472
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1586547711
transform 1 0 400 0 -1 8560
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1586547711
transform 1 0 400 0 1 7472
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_473
timestamp 1586547711
transform 1 0 676 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1670
timestamp 1586547711
transform 1 0 860 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1590
timestamp 1586547711
transform 1 0 768 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1496
timestamp 1586547711
transform 1 0 952 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL1380x35360
timestamp 1586547711
transform 1 0 676 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1498
timestamp 1586547711
transform 1 0 1136 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL3220x38080
timestamp 1586547711
transform 1 0 1044 0 -1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL4600x38080
timestamp 1586547711
transform 1 0 1320 0 -1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _805_
timestamp 1586547711
transform 1 0 1136 0 1 7472
box 0 -48 552 592
use sky130_fd_sc_hd__a21o_4  _757_
timestamp 1586547711
transform 1 0 1412 0 -1 8560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL10580x38080
timestamp 1586547711
transform 1 0 2516 0 -1 8560
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL10120x35360
timestamp 1586547711
transform 1 0 2424 0 1 7472
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_295
timestamp 1586547711
transform 1 0 1688 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_472
timestamp 1586547711
transform 1 0 1872 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1440
timestamp 1586547711
transform 1 0 2056 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1489
timestamp 1586547711
transform 1 0 2240 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL17940x38080
timestamp 1586547711
transform 1 0 3988 0 -1 8560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL16560x35360
timestamp 1586547711
transform 1 0 3712 0 1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1495
timestamp 1586547711
transform 1 0 3804 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1434
timestamp 1586547711
transform 1 0 3344 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1438
timestamp 1586547711
transform 1 0 3528 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1586547711
transform 1 0 3252 0 -1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL22080x35360
timestamp 1586547711
transform 1 0 4816 0 1 7472
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL13800x35360
timestamp 1586547711
transform 1 0 3160 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _743_
timestamp 1586547711
transform 1 0 3344 0 -1 8560
box 0 -48 460 592
use sky130_fd_sc_hd__diode_2  ANTENNA_297
timestamp 1586547711
transform 1 0 5276 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_798
timestamp 1586547711
transform 1 0 5460 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_814
timestamp 1586547711
transform 1 0 5644 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL23920x35360
timestamp 1586547711
transform 1 0 5184 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL23460x38080
timestamp 1586547711
transform 1 0 5092 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL27600x38080
timestamp 1586547711
transform 1 0 5920 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL27140x35360
timestamp 1586547711
transform 1 0 5828 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _501_
timestamp 1586547711
transform 1 0 5276 0 -1 8560
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1636
timestamp 1586547711
transform 1 0 6104 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1565
timestamp 1586547711
transform 1 0 6104 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1557
timestamp 1586547711
transform 1 0 6288 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_402
timestamp 1586547711
transform 1 0 6472 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_131
timestamp 1586547711
transform 1 0 6656 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1586547711
transform 1 0 6840 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1586547711
transform 1 0 6012 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL29440x38080
timestamp 1586547711
transform 1 0 6288 0 -1 8560
box 0 -48 552 592
use sky130_fd_sc_hd__o22a_4  _778_
timestamp 1586547711
transform 1 0 6840 0 -1 8560
box 0 -48 1288 592
use sky130_fd_sc_hd__dfstp_4  _865_
timestamp 1586547711
transform 1 0 7024 0 1 7472
box 0 -48 2208 592
use sky130_fd_sc_hd__decap_12  FILL42780x38080
timestamp 1586547711
transform 1 0 8956 0 -1 8560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL44160x35360
timestamp 1586547711
transform 1 0 9232 0 1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL38640x38080
timestamp 1586547711
transform 1 0 8128 0 -1 8560
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1586547711
transform 1 0 8864 0 -1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL48300x38080
timestamp 1586547711
transform 1 0 10060 0 -1 8560
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1586547711
transform 1 0 10796 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_135
timestamp 1586547711
transform 1 0 10980 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_401
timestamp 1586547711
transform 1 0 11164 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1634
timestamp 1586547711
transform 1 0 11348 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL51520x35360
timestamp 1586547711
transform 1 0 10704 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL49680x35360
timestamp 1586547711
transform 1 0 10336 0 1 7472
box 0 -48 368 592
use sky130_fd_sc_hd__dfstp_4  _864_
timestamp 1586547711
transform 1 0 10796 0 -1 8560
box 0 -48 2208 592
use sky130_fd_sc_hd__decap_12  FILL63020x38080
timestamp 1586547711
transform 1 0 13004 0 -1 8560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL56580x35360
timestamp 1586547711
transform 1 0 11716 0 1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL62100x35360
timestamp 1586547711
transform 1 0 12820 0 1 7472
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL55660x35360
timestamp 1586547711
transform 1 0 11532 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL65780x35360
timestamp 1586547711
transform 1 0 13556 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1586547711
transform 1 0 11624 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _505_
timestamp 1586547711
transform 1 0 13648 0 1 7472
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL70840x38080
timestamp 1586547711
transform 1 0 14568 0 -1 8560
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_327
timestamp 1586547711
transform 1 0 14200 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_822
timestamp 1586547711
transform 1 0 14384 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1586547711
transform 1 0 14476 0 -1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL68540x38080
timestamp 1586547711
transform 1 0 14108 0 -1 8560
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILL70840x35360
timestamp 1586547711
transform 1 0 14568 0 1 7472
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL76360x38080
timestamp 1586547711
transform 1 0 15672 0 -1 8560
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1007
timestamp 1586547711
transform 1 0 15580 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1009
timestamp 1586547711
transform 1 0 15764 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL72680x35360
timestamp 1586547711
transform 1 0 14936 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _567_
timestamp 1586547711
transform 1 0 15028 0 1 7472
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL77740x35360
timestamp 1586547711
transform 1 0 15948 0 1 7472
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1042
timestamp 1586547711
transform 1 0 16868 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL81880x38080
timestamp 1586547711
transform 1 0 16776 0 -1 8560
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILL81420x35360
timestamp 1586547711
transform 1 0 16684 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL86480x38080
timestamp 1586547711
transform 1 0 17696 0 -1 8560
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1043
timestamp 1586547711
transform 1 0 17328 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1045
timestamp 1586547711
transform 1 0 17512 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1016
timestamp 1586547711
transform 1 0 17052 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1586547711
transform 1 0 17236 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__and3_4  _577_
timestamp 1586547711
transform 1 0 17328 0 1 7472
box 0 -48 828 592
use sky130_fd_sc_hd__decap_12  FILL89700x35360
timestamp 1586547711
transform 1 0 18340 0 1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL95220x35360
timestamp 1586547711
transform 1 0 19444 0 1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL93840x38080
timestamp 1586547711
transform 1 0 19168 0 -1 8560
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1084
timestamp 1586547711
transform 1 0 18984 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_994
timestamp 1586547711
transform 1 0 18156 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1586547711
transform 1 0 20088 0 -1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL98900x38080
timestamp 1586547711
transform 1 0 20180 0 -1 8560
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL92000x38080
timestamp 1586547711
transform 1 0 18800 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL97520x38080
timestamp 1586547711
transform 1 0 19904 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_127
timestamp 1586547711
transform 1 0 20548 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1085
timestamp 1586547711
transform 1 0 20732 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1118
timestamp 1586547711
transform 1 0 20916 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1126
timestamp 1586547711
transform 1 0 21100 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1131
timestamp 1586547711
transform 1 0 21284 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL108100x38080
timestamp 1586547711
transform 1 0 22020 0 -1 8560
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL105340x35360
timestamp 1586547711
transform 1 0 21468 0 1 7472
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1548
timestamp 1586547711
transform 1 0 22296 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1127
timestamp 1586547711
transform 1 0 22480 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL109020x35360
timestamp 1586547711
transform 1 0 22204 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__o22ai_4  _610_
timestamp 1586547711
transform 1 0 20548 0 -1 8560
box 0 -48 1472 592
use sky130_fd_sc_hd__decap_8  FILL115000x38080
timestamp 1586547711
transform 1 0 23400 0 -1 8560
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1088
timestamp 1586547711
transform 1 0 22664 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_328
timestamp 1586547711
transform 1 0 23492 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1586547711
transform 1 0 22848 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _776_
timestamp 1586547711
transform 1 0 22940 0 1 7472
box 0 -48 552 592
use sky130_fd_sc_hd__and2_4  _774_
timestamp 1586547711
transform 1 0 22756 0 -1 8560
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  FILL118680x38080
timestamp 1586547711
transform 1 0 24136 0 -1 8560
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_817
timestamp 1586547711
transform 1 0 23768 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_362
timestamp 1586547711
transform 1 0 23952 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_116
timestamp 1586547711
transform 1 0 24136 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL116380x35360
timestamp 1586547711
transform 1 0 23676 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _593_
timestamp 1586547711
transform 1 0 24412 0 -1 8560
box 0 -48 552 592
use sky130_fd_sc_hd__o22a_4  _783_
timestamp 1586547711
transform 1 0 24320 0 1 7472
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL126040x35360
timestamp 1586547711
transform 1 0 25608 0 1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL126960x38080
timestamp 1586547711
transform 1 0 25792 0 -1 8560
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1551
timestamp 1586547711
transform 1 0 24964 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1586547711
transform 1 0 25700 0 -1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL123740x38080
timestamp 1586547711
transform 1 0 25148 0 -1 8560
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL131560x35360
timestamp 1586547711
transform 1 0 26712 0 1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1185
timestamp 1586547711
transform 1 0 26068 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1230
timestamp 1586547711
transform 1 0 26252 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_729
timestamp 1586547711
transform 1 0 26436 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1123
timestamp 1586547711
transform 1 0 26620 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1197
timestamp 1586547711
transform 1 0 26804 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL134780x38080
timestamp 1586547711
transform 1 0 27356 0 -1 8560
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1199
timestamp 1586547711
transform 1 0 26988 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1200
timestamp 1586547711
transform 1 0 27172 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILL138460x38080
timestamp 1586547711
transform 1 0 28092 0 -1 8560
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL137080x35360
timestamp 1586547711
transform 1 0 27816 0 1 7472
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1218
timestamp 1586547711
transform 1 0 28368 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1125
timestamp 1586547711
transform 1 0 28092 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1120
timestamp 1586547711
transform 1 0 28276 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_998
timestamp 1586547711
transform 1 0 29104 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL140760x38080
timestamp 1586547711
transform 1 0 28552 0 -1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1586547711
transform 1 0 28460 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _608_
timestamp 1586547711
transform 1 0 28644 0 -1 8560
box 0 -48 552 592
use sky130_fd_sc_hd__buf_4  _609_
timestamp 1586547711
transform 1 0 28552 0 1 7472
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1000
timestamp 1586547711
transform 1 0 29196 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1186
timestamp 1586547711
transform 1 0 29380 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1119
timestamp 1586547711
transform 1 0 29288 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_996
timestamp 1586547711
transform 1 0 29932 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1001
timestamp 1586547711
transform 1 0 30116 0 1 7472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL147200x35360
timestamp 1586547711
transform 1 0 29840 0 1 7472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL145820x38080
timestamp 1586547711
transform 1 0 29564 0 -1 8560
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILL145360x35360
timestamp 1586547711
transform 1 0 29472 0 1 7472
box 0 -48 368 592
use sky130_fd_sc_hd__inv_4  _565_
timestamp 1586547711
transform 1 0 29932 0 -1 8560
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL149500x35360
timestamp 1586547711
transform 1 0 30300 0 1 7472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL149960x38080
timestamp 1586547711
transform 1 0 30392 0 -1 8560
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1586547711
transform 1 0 31312 0 -1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL153640x38080
timestamp 1586547711
transform 1 0 31128 0 -1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1586547711
transform 1 0 31404 0 -1 8560
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1586547711
transform 1 0 31404 0 1 7472
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1586547711
transform 1 0 400 0 1 8560
box 0 -48 276 592
use sky130_fd_sc_hd__dfrtp_4  _908_
timestamp 1586547711
transform 1 0 676 0 1 8560
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1488
timestamp 1586547711
transform 1 0 2792 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1441
timestamp 1586547711
transform 1 0 2976 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_474
timestamp 1586547711
transform 1 0 3160 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_299
timestamp 1586547711
transform 1 0 3344 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_298
timestamp 1586547711
transform 1 0 4172 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1436
timestamp 1586547711
transform 1 0 4356 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL20700x40800
timestamp 1586547711
transform 1 0 4540 0 1 8560
box 0 -48 552 592
use sky130_fd_sc_hd__and2_4  _756_
timestamp 1586547711
transform 1 0 3528 0 1 8560
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_818
timestamp 1586547711
transform 1 0 5092 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_799
timestamp 1586547711
transform 1 0 5276 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_301
timestamp 1586547711
transform 1 0 5460 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_129
timestamp 1586547711
transform 1 0 5644 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1586547711
transform 1 0 5828 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1586547711
transform 1 0 6012 0 1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__dfstp_4  _866_
timestamp 1586547711
transform 1 0 6104 0 1 8560
box 0 -48 2208 592
use sky130_fd_sc_hd__decap_3  FILL43240x40800
timestamp 1586547711
transform 1 0 9048 0 1 8560
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL39560x40800
timestamp 1586547711
transform 1 0 8312 0 1 8560
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_122
timestamp 1586547711
transform 1 0 9324 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_358
timestamp 1586547711
transform 1 0 9508 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_809
timestamp 1586547711
transform 1 0 9692 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1560
timestamp 1586547711
transform 1 0 9876 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL49220x40800
timestamp 1586547711
transform 1 0 10244 0 1 8560
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1568
timestamp 1586547711
transform 1 0 10060 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1556
timestamp 1586547711
transform 1 0 11072 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_400
timestamp 1586547711
transform 1 0 11256 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_134
timestamp 1586547711
transform 1 0 11440 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL52900x40800
timestamp 1586547711
transform 1 0 10980 0 1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL63020x40800
timestamp 1586547711
transform 1 0 13004 0 1 8560
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1586547711
transform 1 0 11624 0 1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _777_
timestamp 1586547711
transform 1 0 11716 0 1 8560
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_3  FILL68540x40800
timestamp 1586547711
transform 1 0 14108 0 1 8560
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL75900x40800
timestamp 1586547711
transform 1 0 15580 0 1 8560
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1017
timestamp 1586547711
transform 1 0 14384 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_865
timestamp 1586547711
transform 1 0 15212 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_933
timestamp 1586547711
transform 1 0 15396 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_841
timestamp 1586547711
transform 1 0 15856 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _569_
timestamp 1586547711
transform 1 0 14568 0 1 8560
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  FILL80040x40800
timestamp 1586547711
transform 1 0 16408 0 1 8560
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_863
timestamp 1586547711
transform 1 0 16040 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_866
timestamp 1586547711
transform 1 0 16224 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1044
timestamp 1586547711
transform 1 0 16684 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1002
timestamp 1586547711
transform 1 0 16868 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_995
timestamp 1586547711
transform 1 0 17052 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_133
timestamp 1586547711
transform 1 0 17328 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1586547711
transform 1 0 17236 0 1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _564_
timestamp 1586547711
transform 1 0 17512 0 1 8560
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_722
timestamp 1586547711
transform 1 0 18064 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL99360x40800
timestamp 1586547711
transform 1 0 20272 0 1 8560
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_993
timestamp 1586547711
transform 1 0 18248 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1100
timestamp 1586547711
transform 1 0 18432 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_723
timestamp 1586547711
transform 1 0 18616 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_130
timestamp 1586547711
transform 1 0 18800 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__a211o_4  _600_
timestamp 1586547711
transform 1 0 18984 0 1 8560
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL104880x40800
timestamp 1586547711
transform 1 0 21376 0 1 8560
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1586547711
transform 1 0 22480 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_126
timestamp 1586547711
transform 1 0 22664 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_357
timestamp 1586547711
transform 1 0 22940 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1637
timestamp 1586547711
transform 1 0 23124 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1586547711
transform 1 0 22848 0 1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL114540x40800
timestamp 1586547711
transform 1 0 23308 0 1 8560
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1154
timestamp 1586547711
transform 1 0 23676 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1152
timestamp 1586547711
transform 1 0 23860 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1121
timestamp 1586547711
transform 1 0 24044 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1086
timestamp 1586547711
transform 1 0 24228 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _621_
timestamp 1586547711
transform 1 0 24412 0 1 8560
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1005
timestamp 1586547711
transform 1 0 25700 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_999
timestamp 1586547711
transform 1 0 25884 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_91
timestamp 1586547711
transform 1 0 26068 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_115
timestamp 1586547711
transform 1 0 26252 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__a211o_4  _637_
timestamp 1586547711
transform 1 0 26436 0 1 8560
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1184
timestamp 1586547711
transform 1 0 27908 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1124
timestamp 1586547711
transform 1 0 28092 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1004
timestamp 1586547711
transform 1 0 28276 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_94
timestamp 1586547711
transform 1 0 28552 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_118
timestamp 1586547711
transform 1 0 28736 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL142600x40800
timestamp 1586547711
transform 1 0 28920 0 1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1586547711
transform 1 0 28460 0 1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL136620x40800
timestamp 1586547711
transform 1 0 27724 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__and3_4  _661_
timestamp 1586547711
transform 1 0 29012 0 1 8560
box 0 -48 828 592
use sky130_fd_sc_hd__decap_12  FILL149040x40800
timestamp 1586547711
transform 1 0 30208 0 1 8560
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_88
timestamp 1586547711
transform 1 0 29840 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1246
timestamp 1586547711
transform 1 0 30024 0 1 8560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL154560x40800
timestamp 1586547711
transform 1 0 31312 0 1 8560
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1586547711
transform 1 0 31404 0 1 8560
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1586547711
transform 1 0 400 0 -1 9648
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL9200x43520
timestamp 1586547711
transform 1 0 2240 0 -1 9648
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_300
timestamp 1586547711
transform 1 0 676 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1499
timestamp 1586547711
transform 1 0 860 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1591
timestamp 1586547711
transform 1 0 1688 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1671
timestamp 1586547711
transform 1 0 2056 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL3220x43520
timestamp 1586547711
transform 1 0 1044 0 -1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL7360x43520
timestamp 1586547711
transform 1 0 1872 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _806_
timestamp 1586547711
transform 1 0 1136 0 -1 9648
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILL12880x43520
timestamp 1586547711
transform 1 0 2976 0 -1 9648
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL20240x43520
timestamp 1586547711
transform 1 0 4448 0 -1 9648
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1586547711
transform 1 0 3252 0 -1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__a21o_4  _759_
timestamp 1586547711
transform 1 0 3344 0 -1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL29440x43520
timestamp 1586547711
transform 1 0 6288 0 -1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL23920x43520
timestamp 1586547711
transform 1 0 5184 0 -1 9648
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_355
timestamp 1586547711
transform 1 0 6104 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _503_
timestamp 1586547711
transform 1 0 5460 0 -1 9648
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL34960x43520
timestamp 1586547711
transform 1 0 7392 0 -1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1638
timestamp 1586547711
transform 1 0 8956 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1586547711
transform 1 0 8864 0 -1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL40480x43520
timestamp 1586547711
transform 1 0 8496 0 -1 9648
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL43700x43520
timestamp 1586547711
transform 1 0 9140 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL51060x43520
timestamp 1586547711
transform 1 0 10612 0 -1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__o22a_4  _781_
timestamp 1586547711
transform 1 0 9324 0 -1 9648
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL58420x43520
timestamp 1586547711
transform 1 0 12084 0 -1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL63940x43520
timestamp 1586547711
transform 1 0 13188 0 -1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_929
timestamp 1586547711
transform 1 0 11716 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1564
timestamp 1586547711
transform 1 0 11900 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL71760x43520
timestamp 1586547711
transform 1 0 14752 0 -1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_914
timestamp 1586547711
transform 1 0 14568 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1586547711
transform 1 0 14476 0 -1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL69460x43520
timestamp 1586547711
transform 1 0 14292 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _519_
timestamp 1586547711
transform 1 0 15856 0 -1 9648
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL80500x43520
timestamp 1586547711
transform 1 0 16500 0 -1 9648
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL84180x43520
timestamp 1586547711
transform 1 0 17236 0 -1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__a211o_4  _578_
timestamp 1586547711
transform 1 0 17328 0 -1 9648
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL98900x43520
timestamp 1586547711
transform 1 0 20180 0 -1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL94760x43520
timestamp 1586547711
transform 1 0 19352 0 -1 9648
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_855
timestamp 1586547711
transform 1 0 18616 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_861
timestamp 1586547711
transform 1 0 18800 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_333
timestamp 1586547711
transform 1 0 18984 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1101
timestamp 1586547711
transform 1 0 19168 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1586547711
transform 1 0 20088 0 -1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL104420x43520
timestamp 1586547711
transform 1 0 21284 0 -1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL109940x43520
timestamp 1586547711
transform 1 0 22388 0 -1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__dfstp_4  _867_
timestamp 1586547711
transform 1 0 22480 0 -1 9648
box 0 -48 2208 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1155
timestamp 1586547711
transform 1 0 24688 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL122360x43520
timestamp 1586547711
transform 1 0 24872 0 -1 9648
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1153
timestamp 1586547711
transform 1 0 25792 0 -1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL126040x43520
timestamp 1586547711
transform 1 0 25608 0 -1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL127880x43520
timestamp 1586547711
transform 1 0 25976 0 -1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1586547711
transform 1 0 25700 0 -1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__a32o_4  _652_ ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 26068 0 -1 9648
box 0 -48 1564 592
use sky130_fd_sc_hd__decap_8  FILL136160x43520
timestamp 1586547711
transform 1 0 27632 0 -1 9648
box 0 -48 736 592
use sky130_fd_sc_hd__a32o_4  _645_
timestamp 1586547711
transform 1 0 28368 0 -1 9648
box 0 -48 1564 592
use sky130_fd_sc_hd__decap_12  FILL147660x43520
timestamp 1586547711
transform 1 0 29932 0 -1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL153180x43520
timestamp 1586547711
transform 1 0 31036 0 -1 9648
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1586547711
transform 1 0 31312 0 -1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1586547711
transform 1 0 31404 0 -1 9648
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1586547711
transform 1 0 400 0 1 9648
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL5060x46240
timestamp 1586547711
transform 1 0 1412 0 1 9648
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL1380x46240
timestamp 1586547711
transform 1 0 676 0 1 9648
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_475
timestamp 1586547711
transform 1 0 1688 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_303
timestamp 1586547711
transform 1 0 1872 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _909_
timestamp 1586547711
transform 1 0 2056 0 1 9648
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_12  FILL21620x46240
timestamp 1586547711
transform 1 0 4724 0 1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_302
timestamp 1586547711
transform 1 0 4172 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1437
timestamp 1586547711
transform 1 0 4356 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1494
timestamp 1586547711
transform 1 0 4540 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL28520x46240
timestamp 1586547711
transform 1 0 6104 0 1 9648
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_148
timestamp 1586547711
transform 1 0 6840 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_390
timestamp 1586547711
transform 1 0 7024 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1586547711
transform 1 0 6012 0 1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL27140x46240
timestamp 1586547711
transform 1 0 5828 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_741
timestamp 1586547711
transform 1 0 7208 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_753
timestamp 1586547711
transform 1 0 7392 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_801
timestamp 1586547711
transform 1 0 7576 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_359
timestamp 1586547711
transform 1 0 8220 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_123
timestamp 1586547711
transform 1 0 8404 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1586547711
transform 1 0 8588 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL38640x46240
timestamp 1586547711
transform 1 0 8128 0 1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL36800x46240
timestamp 1586547711
transform 1 0 7760 0 1 9648
box 0 -48 368 592
use sky130_fd_sc_hd__dfrtp_4  _868_
timestamp 1586547711
transform 1 0 8772 0 1 9648
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_8  FILL52440x46240
timestamp 1586547711
transform 1 0 10888 0 1 9648
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILL56580x46240
timestamp 1586547711
transform 1 0 11716 0 1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_986
timestamp 1586547711
transform 1 0 13280 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_988
timestamp 1586547711
transform 1 0 13464 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL63940x46240
timestamp 1586547711
transform 1 0 13188 0 1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1586547711
transform 1 0 11624 0 1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL62100x46240
timestamp 1586547711
transform 1 0 12820 0 1 9648
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILL66240x46240
timestamp 1586547711
transform 1 0 13648 0 1 9648
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1006
timestamp 1586547711
transform 1 0 14016 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_892
timestamp 1586547711
transform 1 0 14200 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_864
timestamp 1586547711
transform 1 0 14384 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_670
timestamp 1586547711
transform 1 0 15212 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_710
timestamp 1586547711
transform 1 0 15396 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL75900x46240
timestamp 1586547711
transform 1 0 15580 0 1 9648
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _530_
timestamp 1586547711
transform 1 0 14568 0 1 9648
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_987
timestamp 1586547711
transform 1 0 16040 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_991
timestamp 1586547711
transform 1 0 16224 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1046
timestamp 1586547711
transform 1 0 16408 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL77740x46240
timestamp 1586547711
transform 1 0 15948 0 1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1047
timestamp 1586547711
transform 1 0 16592 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_842
timestamp 1586547711
transform 1 0 16868 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_669
timestamp 1586547711
transform 1 0 17052 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL81880x46240
timestamp 1586547711
transform 1 0 16776 0 1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1586547711
transform 1 0 17236 0 1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _563_
timestamp 1586547711
transform 1 0 17328 0 1 9648
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_160
timestamp 1586547711
transform 1 0 18064 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL87860x46240
timestamp 1586547711
transform 1 0 17972 0 1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_332
timestamp 1586547711
transform 1 0 18248 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_772
timestamp 1586547711
transform 1 0 18432 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_162
timestamp 1586547711
transform 1 0 18616 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp 1586547711
transform 1 0 18800 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__dfstp_4  _890_
timestamp 1586547711
transform 1 0 18984 0 1 9648
box 0 -48 2208 592
use sky130_fd_sc_hd__decap_12  FILL103960x46240
timestamp 1586547711
transform 1 0 21192 0 1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1559
timestamp 1586547711
transform 1 0 22296 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_356
timestamp 1586547711
transform 1 0 22480 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL119140x46240
timestamp 1586547711
transform 1 0 24228 0 1 9648
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_125
timestamp 1586547711
transform 1 0 22664 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1586547711
transform 1 0 22848 0 1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _780_
timestamp 1586547711
transform 1 0 22940 0 1 9648
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL131560x46240
timestamp 1586547711
transform 1 0 26712 0 1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1198
timestamp 1586547711
transform 1 0 25148 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1122
timestamp 1586547711
transform 1 0 25332 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_124
timestamp 1586547711
transform 1 0 25516 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_121
timestamp 1586547711
transform 1 0 26528 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL122820x46240
timestamp 1586547711
transform 1 0 24964 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _636_ ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 25700 0 1 9648
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1247
timestamp 1586547711
transform 1 0 27908 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_731
timestamp 1586547711
transform 1 0 28092 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_112
timestamp 1586547711
transform 1 0 28276 0 1 9648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL137080x46240
timestamp 1586547711
transform 1 0 27816 0 1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1586547711
transform 1 0 28460 0 1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__a211o_4  _662_
timestamp 1586547711
transform 1 0 28552 0 1 9648
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL147200x46240
timestamp 1586547711
transform 1 0 29840 0 1 9648
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL154560x46240
timestamp 1586547711
transform 1 0 31312 0 1 9648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL152720x46240
timestamp 1586547711
transform 1 0 30944 0 1 9648
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1586547711
transform 1 0 31404 0 1 9648
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL1380x48960
timestamp 1586547711
transform 1 0 676 0 -1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1586547711
transform 1 0 400 0 -1 10736
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL6900x48960
timestamp 1586547711
transform 1 0 1780 0 -1 10736
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL9200x48960
timestamp 1586547711
transform 1 0 2240 0 -1 10736
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1504
timestamp 1586547711
transform 1 0 2056 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL19780x48960
timestamp 1586547711
transform 1 0 4356 0 -1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL12880x48960
timestamp 1586547711
transform 1 0 2976 0 -1 10736
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1586547711
transform 1 0 3252 0 -1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL14720x48960
timestamp 1586547711
transform 1 0 3344 0 -1 10736
box 0 -48 368 592
use sky130_fd_sc_hd__and2_4  _758_
timestamp 1586547711
transform 1 0 3712 0 -1 10736
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1629
timestamp 1586547711
transform 1 0 6104 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL28060x48960
timestamp 1586547711
transform 1 0 6012 0 -1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL25300x48960
timestamp 1586547711
transform 1 0 5460 0 -1 10736
box 0 -48 552 592
use sky130_fd_sc_hd__decap_6  FILL29440x48960
timestamp 1586547711
transform 1 0 6288 0 -1 10736
box 0 -48 552 592
use sky130_fd_sc_hd__o22a_4  _496_
timestamp 1586547711
transform 1 0 6840 0 -1 10736
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL43700x48960
timestamp 1586547711
transform 1 0 9140 0 -1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL38640x48960
timestamp 1586547711
transform 1 0 8128 0 -1 10736
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_780
timestamp 1586547711
transform 1 0 8956 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1586547711
transform 1 0 8864 0 -1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL49220x48960
timestamp 1586547711
transform 1 0 10244 0 -1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL54740x48960
timestamp 1586547711
transform 1 0 11348 0 -1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_922
timestamp 1586547711
transform 1 0 12452 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_921
timestamp 1586547711
transform 1 0 12636 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_989
timestamp 1586547711
transform 1 0 12820 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1049
timestamp 1586547711
transform 1 0 13004 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL63940x48960
timestamp 1586547711
transform 1 0 13188 0 -1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _561_
timestamp 1586547711
transform 1 0 13280 0 -1 10736
box 0 -48 460 592
use sky130_fd_sc_hd__decap_8  FILL66700x48960
timestamp 1586547711
transform 1 0 13740 0 -1 10736
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL74060x48960
timestamp 1586547711
transform 1 0 15212 0 -1 10736
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1586547711
transform 1 0 14476 0 -1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _566_
timestamp 1586547711
transform 1 0 14568 0 -1 10736
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  FILL85560x48960
timestamp 1586547711
transform 1 0 17512 0 -1 10736
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_992
timestamp 1586547711
transform 1 0 17328 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_860
timestamp 1586547711
transform 1 0 17788 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL77740x48960
timestamp 1586547711
transform 1 0 15948 0 -1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL84180x48960
timestamp 1586547711
transform 1 0 17236 0 -1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL87860x48960
timestamp 1586547711
transform 1 0 17972 0 -1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL82340x48960
timestamp 1586547711
transform 1 0 16868 0 -1 10736
box 0 -48 368 592
use sky130_fd_sc_hd__o22a_4  _517_
timestamp 1586547711
transform 1 0 18064 0 -1 10736
box 0 -48 1288 592
use sky130_fd_sc_hd__and3_4  _579_
timestamp 1586547711
transform 1 0 16040 0 -1 10736
box 0 -48 828 592
use sky130_fd_sc_hd__decap_12  FILL98900x48960
timestamp 1586547711
transform 1 0 20180 0 -1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1662
timestamp 1586547711
transform 1 0 19352 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1586547711
transform 1 0 20088 0 -1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL95680x48960
timestamp 1586547711
transform 1 0 19536 0 -1 10736
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL104420x48960
timestamp 1586547711
transform 1 0 21284 0 -1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILL109940x48960
timestamp 1586547711
transform 1 0 22388 0 -1 10736
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL114540x48960
timestamp 1586547711
transform 1 0 23308 0 -1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL120060x48960
timestamp 1586547711
transform 1 0 24412 0 -1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_804
timestamp 1586547711
transform 1 0 22940 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1567
timestamp 1586547711
transform 1 0 23124 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_380
timestamp 1586547711
transform 1 0 26436 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_816
timestamp 1586547711
transform 1 0 26620 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1194
timestamp 1586547711
transform 1 0 26804 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1586547711
transform 1 0 25700 0 -1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL125580x48960
timestamp 1586547711
transform 1 0 25516 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL129260x48960
timestamp 1586547711
transform 1 0 26252 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _620_
timestamp 1586547711
transform 1 0 25792 0 -1 10736
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL133860x48960
timestamp 1586547711
transform 1 0 27172 0 -1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL142600x48960
timestamp 1586547711
transform 1 0 28920 0 -1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL139380x48960
timestamp 1586547711
transform 1 0 28276 0 -1 10736
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1649
timestamp 1586547711
transform 1 0 26988 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1087
timestamp 1586547711
transform 1 0 28552 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1248
timestamp 1586547711
transform 1 0 28736 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL148120x48960
timestamp 1586547711
transform 1 0 30024 0 -1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1586547711
transform 1 0 31312 0 -1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL153640x48960
timestamp 1586547711
transform 1 0 31128 0 -1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1586547711
transform 1 0 31404 0 -1 10736
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1586547711
transform 1 0 400 0 -1 11824
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1586547711
transform 1 0 400 0 1 10736
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_196
timestamp 1586547711
transform 1 0 1228 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_201
timestamp 1586547711
transform 1 0 1412 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL1380x54400
timestamp 1586547711
transform 1 0 676 0 -1 11824
box 0 -48 552 592
use sky130_fd_sc_hd__decap_6  FILL1380x51680
timestamp 1586547711
transform 1 0 676 0 1 10736
box 0 -48 552 592
use sky130_fd_sc_hd__buf_2  _850_ ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 1228 0 -1 11824
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL5980x54400
timestamp 1586547711
transform 1 0 1596 0 -1 11824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL5980x51680
timestamp 1586547711
transform 1 0 1596 0 1 10736
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL9660x51680
timestamp 1586547711
transform 1 0 2332 0 1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _807_
timestamp 1586547711
transform 1 0 2424 0 1 10736
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL14720x54400
timestamp 1586547711
transform 1 0 3344 0 -1 11824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL20240x54400
timestamp 1586547711
transform 1 0 4448 0 -1 11824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL14720x51680
timestamp 1586547711
transform 1 0 3344 0 1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL20240x51680
timestamp 1586547711
transform 1 0 4448 0 1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1503
timestamp 1586547711
transform 1 0 2976 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1592
timestamp 1586547711
transform 1 0 3160 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1586547711
transform 1 0 3252 0 -1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL11500x54400
timestamp 1586547711
transform 1 0 2700 0 -1 11824
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_393
timestamp 1586547711
transform 1 0 5920 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_150
timestamp 1586547711
transform 1 0 5644 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1586547711
transform 1 0 5828 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL25760x51680
timestamp 1586547711
transform 1 0 5552 0 1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL25760x54400
timestamp 1586547711
transform 1 0 5552 0 -1 11824
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL32200x54400
timestamp 1586547711
transform 1 0 6840 0 -1 11824
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_391
timestamp 1586547711
transform 1 0 6104 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_392
timestamp 1586547711
transform 1 0 6288 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_754
timestamp 1586547711
transform 1 0 6472 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_806
timestamp 1586547711
transform 1 0 6656 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1586547711
transform 1 0 6012 0 1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__dfstp_4  _859_
timestamp 1586547711
transform 1 0 6104 0 1 10736
box 0 -48 2208 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1627
timestamp 1586547711
transform 1 0 8128 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL37720x54400
timestamp 1586547711
transform 1 0 7944 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILL39560x51680
timestamp 1586547711
transform 1 0 8312 0 1 10736
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_751
timestamp 1586547711
transform 1 0 8588 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_739
timestamp 1586547711
transform 1 0 8772 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_154
timestamp 1586547711
transform 1 0 8956 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_374
timestamp 1586547711
transform 1 0 9140 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1586547711
transform 1 0 8864 0 -1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL39560x54400
timestamp 1586547711
transform 1 0 8312 0 -1 11824
box 0 -48 552 592
use sky130_fd_sc_hd__o22a_4  _490_
timestamp 1586547711
transform 1 0 8956 0 -1 11824
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL50140x54400
timestamp 1586547711
transform 1 0 10428 0 -1 11824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL49220x51680
timestamp 1586547711
transform 1 0 10244 0 1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL54740x51680
timestamp 1586547711
transform 1 0 11348 0 1 10736
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1664
timestamp 1586547711
transform 1 0 10244 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_149
timestamp 1586547711
transform 1 0 9876 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1157
timestamp 1586547711
transform 1 0 10060 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL44620x51680
timestamp 1586547711
transform 1 0 9324 0 1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _622_
timestamp 1586547711
transform 1 0 9416 0 1 10736
box 0 -48 460 592
use sky130_fd_sc_hd__decap_8  FILL55660x54400
timestamp 1586547711
transform 1 0 11532 0 -1 11824
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1048
timestamp 1586547711
transform 1 0 11900 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_920
timestamp 1586547711
transform 1 0 12084 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_826
timestamp 1586547711
transform 1 0 12268 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_170
timestamp 1586547711
transform 1 0 12452 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1586547711
transform 1 0 11624 0 1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL59340x54400
timestamp 1586547711
transform 1 0 12268 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL56580x51680
timestamp 1586547711
transform 1 0 11716 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _540_
timestamp 1586547711
transform 1 0 12452 0 -1 11824
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL63480x54400
timestamp 1586547711
transform 1 0 13096 0 -1 11824
box 0 -48 1104 592
use sky130_fd_sc_hd__a211o_4  _580_
timestamp 1586547711
transform 1 0 12636 0 1 10736
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL70840x54400
timestamp 1586547711
transform 1 0 14568 0 -1 11824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL69000x54400
timestamp 1586547711
transform 1 0 14200 0 -1 11824
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_985
timestamp 1586547711
transform 1 0 14476 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1586547711
transform 1 0 14476 0 -1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL67620x51680
timestamp 1586547711
transform 1 0 13924 0 1 10736
box 0 -48 552 592
use sky130_fd_sc_hd__or2_4  _560_
timestamp 1586547711
transform 1 0 14660 0 1 10736
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL76360x51680
timestamp 1586547711
transform 1 0 15672 0 1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_668
timestamp 1586547711
transform 1 0 15304 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_932
timestamp 1586547711
transform 1 0 15488 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL76360x54400
timestamp 1586547711
transform 1 0 15672 0 -1 11824
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL80960x54400
timestamp 1586547711
transform 1 0 16592 0 -1 11824
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1052
timestamp 1586547711
transform 1 0 16224 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1053
timestamp 1586547711
transform 1 0 16408 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILL84640x54400
timestamp 1586547711
transform 1 0 17328 0 -1 11824
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL83720x51680
timestamp 1586547711
transform 1 0 17144 0 1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL84640x51680
timestamp 1586547711
transform 1 0 17328 0 1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1586547711
transform 1 0 17236 0 1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL81880x51680
timestamp 1586547711
transform 1 0 16776 0 1 10736
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILL88320x54400
timestamp 1586547711
transform 1 0 18064 0 -1 11824
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_857
timestamp 1586547711
transform 1 0 17420 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_854
timestamp 1586547711
transform 1 0 17604 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _515_
timestamp 1586547711
transform 1 0 17604 0 -1 11824
box 0 -48 460 592
use sky130_fd_sc_hd__and2_4  _516_
timestamp 1586547711
transform 1 0 17788 0 1 10736
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL92000x51680
timestamp 1586547711
transform 1 0 18800 0 1 10736
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_824
timestamp 1586547711
transform 1 0 18432 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_858
timestamp 1586547711
transform 1 0 18616 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL92000x54400
timestamp 1586547711
transform 1 0 18800 0 -1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL93380x54400
timestamp 1586547711
transform 1 0 19076 0 -1 11824
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_981
timestamp 1586547711
transform 1 0 18892 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL95680x51680
timestamp 1586547711
transform 1 0 19536 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILL97060x54400
timestamp 1586547711
transform 1 0 19812 0 -1 11824
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_990
timestamp 1586547711
transform 1 0 19720 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_717
timestamp 1586547711
transform 1 0 19904 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1586547711
transform 1 0 20088 0 -1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL98900x54400
timestamp 1586547711
transform 1 0 20180 0 -1 11824
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _562_
timestamp 1586547711
transform 1 0 20088 0 1 10736
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_750
timestamp 1586547711
transform 1 0 20640 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_158
timestamp 1586547711
transform 1 0 20732 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1586547711
transform 1 0 20916 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_159
timestamp 1586547711
transform 1 0 21100 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_353
timestamp 1586547711
transform 1 0 21284 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL100740x54400
timestamp 1586547711
transform 1 0 20548 0 -1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL102120x54400
timestamp 1586547711
transform 1 0 20824 0 -1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL106260x51680
timestamp 1586547711
transform 1 0 21652 0 1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1626
timestamp 1586547711
transform 1 0 21468 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__dfstp_4  _856_
timestamp 1586547711
transform 1 0 20916 0 -1 11824
box 0 -48 2208 592
use sky130_fd_sc_hd__decap_12  FILL112700x51680
timestamp 1586547711
transform 1 0 22940 0 1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1631
timestamp 1586547711
transform 1 0 23492 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL111780x51680
timestamp 1586547711
transform 1 0 22756 0 1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1586547711
transform 1 0 22848 0 1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL113620x54400
timestamp 1586547711
transform 1 0 23124 0 -1 11824
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL120060x54400
timestamp 1586547711
transform 1 0 24412 0 -1 11824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL118220x51680
timestamp 1586547711
transform 1 0 24044 0 1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_142
timestamp 1586547711
transform 1 0 23676 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_394
timestamp 1586547711
transform 1 0 23860 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_745
timestamp 1586547711
transform 1 0 24044 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_811
timestamp 1586547711
transform 1 0 24228 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1512
timestamp 1586547711
transform 1 0 25516 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_381
timestamp 1586547711
transform 1 0 25700 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1586547711
transform 1 0 25700 0 -1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL123740x51680
timestamp 1586547711
transform 1 0 25148 0 1 10736
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILL126960x54400
timestamp 1586547711
transform 1 0 25792 0 -1 11824
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILL125580x54400
timestamp 1586547711
transform 1 0 25516 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_93
timestamp 1586547711
transform 1 0 25884 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_92
timestamp 1586547711
transform 1 0 26068 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1586547711
transform 1 0 26252 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _772_
timestamp 1586547711
transform 1 0 26436 0 1 10736
box 0 -48 1288 592
use sky130_fd_sc_hd__dfstp_4  _878_
timestamp 1586547711
transform 1 0 26344 0 -1 11824
box 0 -48 2208 592
use sky130_fd_sc_hd__decap_8  FILL136620x51680
timestamp 1586547711
transform 1 0 27724 0 1 10736
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL140760x51680
timestamp 1586547711
transform 1 0 28552 0 1 10736
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_382
timestamp 1586547711
transform 1 0 28552 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_820
timestamp 1586547711
transform 1 0 28736 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1195
timestamp 1586547711
transform 1 0 28920 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1513
timestamp 1586547711
transform 1 0 29104 0 -1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1586547711
transform 1 0 28460 0 1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL149040x51680
timestamp 1586547711
transform 1 0 30208 0 1 10736
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_95
timestamp 1586547711
transform 1 0 29288 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_378
timestamp 1586547711
transform 1 0 29472 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_812
timestamp 1586547711
transform 1 0 29656 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1193
timestamp 1586547711
transform 1 0 29840 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1511
timestamp 1586547711
transform 1 0 30024 0 1 10736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL150880x54400
timestamp 1586547711
transform 1 0 30576 0 -1 11824
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL154560x51680
timestamp 1586547711
transform 1 0 31312 0 1 10736
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1586547711
transform 1 0 31312 0 -1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _771_
timestamp 1586547711
transform 1 0 29288 0 -1 11824
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1586547711
transform 1 0 31404 0 -1 11824
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1586547711
transform 1 0 31404 0 1 10736
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1586547711
transform 1 0 400 0 1 11824
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_178
timestamp 1586547711
transform 1 0 1504 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1505
timestamp 1586547711
transform 1 0 1688 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1593
timestamp 1586547711
transform 1 0 1872 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1594
timestamp 1586547711
transform 1 0 2516 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL10120x57120
timestamp 1586547711
transform 1 0 2424 0 1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL8280x57120
timestamp 1586547711
transform 1 0 2056 0 1 11824
box 0 -48 368 592
use sky130_fd_sc_hd__conb_1  _831_
timestamp 1586547711
transform 1 0 1228 0 1 11824
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILL1380x57120
timestamp 1586547711
transform 1 0 676 0 1 11824
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL17480x57120
timestamp 1586547711
transform 1 0 3896 0 1 11824
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_511
timestamp 1586547711
transform 1 0 3344 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1507
timestamp 1586547711
transform 1 0 3528 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1589
timestamp 1586547711
transform 1 0 3712 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_510
timestamp 1586547711
transform 1 0 4632 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1583
timestamp 1586547711
transform 1 0 4816 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL14260x57120
timestamp 1586547711
transform 1 0 3252 0 1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _809_
timestamp 1586547711
transform 1 0 2700 0 1 11824
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1630
timestamp 1586547711
transform 1 0 5092 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_742
timestamp 1586547711
transform 1 0 5276 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_147
timestamp 1586547711
transform 1 0 5460 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_145
timestamp 1586547711
transform 1 0 5644 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1586547711
transform 1 0 5828 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL23000x57120
timestamp 1586547711
transform 1 0 5000 0 1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1586547711
transform 1 0 6012 0 1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _498_
timestamp 1586547711
transform 1 0 6104 0 1 11824
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA_156
timestamp 1586547711
transform 1 0 7760 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1586547711
transform 1 0 7944 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL34960x57120
timestamp 1586547711
transform 1 0 7392 0 1 11824
box 0 -48 368 592
use sky130_fd_sc_hd__dfstp_4  _857_
timestamp 1586547711
transform 1 0 8128 0 1 11824
box 0 -48 2208 592
use sky130_fd_sc_hd__decap_8  FILL52440x57120
timestamp 1586547711
transform 1 0 10888 0 1 11824
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_40
timestamp 1586547711
transform 1 0 10336 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_168
timestamp 1586547711
transform 1 0 10520 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_407
timestamp 1586547711
transform 1 0 10704 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILL56580x57120
timestamp 1586547711
transform 1 0 11716 0 1 11824
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_919
timestamp 1586547711
transform 1 0 11992 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1586547711
transform 1 0 11624 0 1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _539_
timestamp 1586547711
transform 1 0 12176 0 1 11824
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL65320x57120
timestamp 1586547711
transform 1 0 13464 0 1 11824
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_167
timestamp 1586547711
transform 1 0 12728 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_916
timestamp 1586547711
transform 1 0 12912 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_918
timestamp 1586547711
transform 1 0 13096 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_983
timestamp 1586547711
transform 1 0 13280 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL61180x57120
timestamp 1586547711
transform 1 0 12636 0 1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_847
timestamp 1586547711
transform 1 0 14568 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_984
timestamp 1586547711
transform 1 0 14752 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1050
timestamp 1586547711
transform 1 0 14936 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1051
timestamp 1586547711
transform 1 0 15120 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_851
timestamp 1586547711
transform 1 0 15488 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_849
timestamp 1586547711
transform 1 0 15672 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL74520x57120
timestamp 1586547711
transform 1 0 15304 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _512_
timestamp 1586547711
transform 1 0 15856 0 1 11824
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  FILL88320x57120
timestamp 1586547711
transform 1 0 18064 0 1 11824
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL84640x57120
timestamp 1586547711
transform 1 0 17328 0 1 11824
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_164
timestamp 1586547711
transform 1 0 16500 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_823
timestamp 1586547711
transform 1 0 16684 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_850
timestamp 1586547711
transform 1 0 16868 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_859
timestamp 1586547711
transform 1 0 17052 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1586547711
transform 1 0 17236 0 1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1081
timestamp 1586547711
transform 1 0 18340 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_718
timestamp 1586547711
transform 1 0 18524 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_155
timestamp 1586547711
transform 1 0 18708 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_161
timestamp 1586547711
transform 1 0 19536 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_856
timestamp 1586547711
transform 1 0 19720 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_770
timestamp 1586547711
transform 1 0 20088 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_352
timestamp 1586547711
transform 1 0 20272 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL97520x57120
timestamp 1586547711
transform 1 0 19904 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _558_
timestamp 1586547711
transform 1 0 18892 0 1 11824
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_157
timestamp 1586547711
transform 1 0 20456 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_715
timestamp 1586547711
transform 1 0 21928 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_720
timestamp 1586547711
transform 1 0 22112 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL109480x57120
timestamp 1586547711
transform 1 0 22296 0 1 11824
box 0 -48 552 592
use sky130_fd_sc_hd__o22a_4  _487_
timestamp 1586547711
transform 1 0 20640 0 1 11824
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA_734
timestamp 1586547711
transform 1 0 22940 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_144
timestamp 1586547711
transform 1 0 23124 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1586547711
transform 1 0 23308 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1586547711
transform 1 0 22848 0 1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__dfstp_4  _861_
timestamp 1586547711
transform 1 0 23492 0 1 11824
box 0 -48 2208 592
use sky130_fd_sc_hd__decap_8  FILL126500x57120
timestamp 1586547711
transform 1 0 25700 0 1 11824
box 0 -48 736 592
use sky130_fd_sc_hd__buf_4  _478_
timestamp 1586547711
transform 1 0 26436 0 1 11824
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_721
timestamp 1586547711
transform 1 0 26988 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_726
timestamp 1586547711
transform 1 0 27172 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1201
timestamp 1586547711
transform 1 0 27356 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1202
timestamp 1586547711
transform 1 0 27540 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_383
timestamp 1586547711
transform 1 0 27724 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_90
timestamp 1586547711
transform 1 0 27908 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_89
timestamp 1586547711
transform 1 0 28092 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1586547711
transform 1 0 28276 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1586547711
transform 1 0 28460 0 1 11824
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _773_
timestamp 1586547711
transform 1 0 28552 0 1 11824
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL148120x57120
timestamp 1586547711
transform 1 0 30024 0 1 11824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL153640x57120
timestamp 1586547711
transform 1 0 31128 0 1 11824
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1650
timestamp 1586547711
transform 1 0 29840 0 1 11824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1586547711
transform 1 0 31404 0 1 11824
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL6440x59840
timestamp 1586547711
transform 1 0 1688 0 -1 12912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1586547711
transform 1 0 400 0 -1 12912
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILL3220x59840
timestamp 1586547711
transform 1 0 1044 0 -1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL1380x59840
timestamp 1586547711
transform 1 0 676 0 -1 12912
box 0 -48 368 592
use sky130_fd_sc_hd__buf_4  _808_
timestamp 1586547711
transform 1 0 1136 0 -1 12912
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL17480x59840
timestamp 1586547711
transform 1 0 3896 0 -1 12912
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL13800x59840
timestamp 1586547711
transform 1 0 3160 0 -1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1586547711
transform 1 0 3252 0 -1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL11960x59840
timestamp 1586547711
transform 1 0 2792 0 -1 12912
box 0 -48 368 592
use sky130_fd_sc_hd__buf_4  _804_
timestamp 1586547711
transform 1 0 3344 0 -1 12912
box 0 -48 552 592
use sky130_fd_sc_hd__buf_4  _798_
timestamp 1586547711
transform 1 0 4632 0 -1 12912
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL23920x59840
timestamp 1586547711
transform 1 0 5184 0 -1 12912
box 0 -48 736 592
use sky130_fd_sc_hd__dfstp_4  _860_
timestamp 1586547711
transform 1 0 5920 0 -1 12912
box 0 -48 2208 592
use sky130_fd_sc_hd__decap_8  FILL42780x59840
timestamp 1586547711
transform 1 0 8956 0 -1 12912
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_375
timestamp 1586547711
transform 1 0 8128 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1586547711
transform 1 0 8864 0 -1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL39560x59840
timestamp 1586547711
transform 1 0 8312 0 -1 12912
box 0 -48 552 592
use sky130_fd_sc_hd__dfrtp_4  _892_
timestamp 1586547711
transform 1 0 9876 0 -1 12912
box 0 -48 2116 592
use sky130_fd_sc_hd__fill_2  FILL46460x59840
timestamp 1586547711
transform 1 0 9692 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL64860x59840
timestamp 1586547711
transform 1 0 13372 0 -1 12912
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_925
timestamp 1586547711
transform 1 0 11992 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL58880x59840
timestamp 1586547711
transform 1 0 12176 0 -1 12912
box 0 -48 552 592
use sky130_fd_sc_hd__or2_4  _559_
timestamp 1586547711
transform 1 0 12728 0 -1 12912
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_165
timestamp 1586547711
transform 1 0 15396 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_846
timestamp 1586547711
transform 1 0 15580 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_852
timestamp 1586547711
transform 1 0 15764 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1586547711
transform 1 0 14476 0 -1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__and3_4  _581_
timestamp 1586547711
transform 1 0 14568 0 -1 12912
box 0 -48 828 592
use sky130_fd_sc_hd__decap_12  FILL85560x59840
timestamp 1586547711
transform 1 0 17512 0 -1 12912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL77740x59840
timestamp 1586547711
transform 1 0 15948 0 -1 12912
box 0 -48 276 592
use sky130_fd_sc_hd__a211o_4  _582_
timestamp 1586547711
transform 1 0 16224 0 -1 12912
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_8  FILL94760x59840
timestamp 1586547711
transform 1 0 19352 0 -1 12912
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL91080x59840
timestamp 1586547711
transform 1 0 18616 0 -1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1586547711
transform 1 0 20088 0 -1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL98900x59840
timestamp 1586547711
transform 1 0 20180 0 -1 12912
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _592_
timestamp 1586547711
transform 1 0 18708 0 -1 12912
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL107640x59840
timestamp 1586547711
transform 1 0 21928 0 -1 12912
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_738
timestamp 1586547711
transform 1 0 20640 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL100740x59840
timestamp 1586547711
transform 1 0 20548 0 -1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL104880x59840
timestamp 1586547711
transform 1 0 21376 0 -1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL102120x59840
timestamp 1586547711
transform 1 0 20824 0 -1 12912
box 0 -48 552 592
use sky130_fd_sc_hd__inv_4  _477_
timestamp 1586547711
transform 1 0 21468 0 -1 12912
box 0 -48 460 592
use sky130_fd_sc_hd__diode_2  ANTENNA_395
timestamp 1586547711
transform 1 0 23492 0 -1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL115000x59840
timestamp 1586547711
transform 1 0 23400 0 -1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL113160x59840
timestamp 1586547711
transform 1 0 23032 0 -1 12912
box 0 -48 368 592
use sky130_fd_sc_hd__o22a_4  _500_
timestamp 1586547711
transform 1 0 23676 0 -1 12912
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_3  FILL130640x59840
timestamp 1586547711
transform 1 0 26528 0 -1 12912
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL122820x59840
timestamp 1586547711
transform 1 0 24964 0 -1 12912
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL126960x59840
timestamp 1586547711
transform 1 0 25792 0 -1 12912
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1586547711
transform 1 0 25700 0 -1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _638_
timestamp 1586547711
transform 1 0 26804 0 -1 12912
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL134320x59840
timestamp 1586547711
transform 1 0 27264 0 -1 12912
box 0 -48 1104 592
use sky130_fd_sc_hd__dfstp_4  _879_
timestamp 1586547711
transform 1 0 28368 0 -1 12912
box 0 -48 2208 592
use sky130_fd_sc_hd__decap_8  FILL150880x59840
timestamp 1586547711
transform 1 0 30576 0 -1 12912
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1586547711
transform 1 0 31312 0 -1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1586547711
transform 1 0 31404 0 -1 12912
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL1380x62560
timestamp 1586547711
transform 1 0 676 0 1 12912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL6900x62560
timestamp 1586547711
transform 1 0 1780 0 1 12912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1586547711
transform 1 0 400 0 1 12912
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL18400x62560
timestamp 1586547711
transform 1 0 4080 0 1 12912
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_252
timestamp 1586547711
transform 1 0 3344 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_459
timestamp 1586547711
transform 1 0 3528 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1508
timestamp 1586547711
transform 1 0 3712 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1674
timestamp 1586547711
transform 1 0 3896 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL14260x62560
timestamp 1586547711
transform 1 0 3252 0 1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL12420x62560
timestamp 1586547711
transform 1 0 2884 0 1 12912
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL28520x62560
timestamp 1586547711
transform 1 0 6104 0 1 12912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL23920x62560
timestamp 1586547711
transform 1 0 5184 0 1 12912
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL27600x62560
timestamp 1586547711
transform 1 0 5920 0 1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1586547711
transform 1 0 6012 0 1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL34040x62560
timestamp 1586547711
transform 1 0 7208 0 1 12912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL39560x62560
timestamp 1586547711
transform 1 0 8312 0 1 12912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL45080x62560
timestamp 1586547711
transform 1 0 9416 0 1 12912
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_917
timestamp 1586547711
transform 1 0 11072 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_406
timestamp 1586547711
transform 1 0 11256 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_166
timestamp 1586547711
transform 1 0 11440 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL50600x62560
timestamp 1586547711
transform 1 0 10520 0 1 12912
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_834
timestamp 1586547711
transform 1 0 13004 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_912
timestamp 1586547711
transform 1 0 13188 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_915
timestamp 1586547711
transform 1 0 13372 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_848
timestamp 1586547711
transform 1 0 13556 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1586547711
transform 1 0 11624 0 1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _542_
timestamp 1586547711
transform 1 0 11716 0 1 12912
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA_845
timestamp 1586547711
transform 1 0 13740 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_771
timestamp 1586547711
transform 1 0 14384 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_331
timestamp 1586547711
transform 1 0 14568 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_163
timestamp 1586547711
transform 1 0 14752 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp 1586547711
transform 1 0 14936 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _513_
timestamp 1586547711
transform 1 0 15120 0 1 12912
box 0 -48 1288 592
use sky130_fd_sc_hd__inv_4  _511_
timestamp 1586547711
transform 1 0 13924 0 1 12912
box 0 -48 460 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1663
timestamp 1586547711
transform 1 0 16408 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_853
timestamp 1586547711
transform 1 0 17052 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_709
timestamp 1586547711
transform 1 0 17972 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL82800x62560
timestamp 1586547711
transform 1 0 16960 0 1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1586547711
transform 1 0 17236 0 1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL80960x62560
timestamp 1586547711
transform 1 0 16592 0 1 12912
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _514_
timestamp 1586547711
transform 1 0 17328 0 1 12912
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_833
timestamp 1586547711
transform 1 0 18156 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_951
timestamp 1586547711
transform 1 0 18432 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_982
timestamp 1586547711
transform 1 0 18616 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1054
timestamp 1586547711
transform 1 0 18800 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL89700x62560
timestamp 1586547711
transform 1 0 18340 0 1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1055
timestamp 1586547711
transform 1 0 18984 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1102
timestamp 1586547711
transform 1 0 19260 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1082
timestamp 1586547711
transform 1 0 19444 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL93840x62560
timestamp 1586547711
transform 1 0 19168 0 1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__and3_4  _601_
timestamp 1586547711
transform 1 0 19628 0 1 12912
box 0 -48 828 592
use sky130_fd_sc_hd__decap_8  FILL101200x62560
timestamp 1586547711
transform 1 0 20640 0 1 12912
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_952
timestamp 1586547711
transform 1 0 20456 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_151
timestamp 1586547711
transform 1 0 21376 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_388
timestamp 1586547711
transform 1 0 21560 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_740
timestamp 1586547711
transform 1 0 21744 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_752
timestamp 1586547711
transform 1 0 21928 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_789
timestamp 1586547711
transform 1 0 22112 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_749
timestamp 1586547711
transform 1 0 22480 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL109480x62560
timestamp 1586547711
transform 1 0 22296 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_744
timestamp 1586547711
transform 1 0 22664 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_716
timestamp 1586547711
transform 1 0 23492 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1586547711
transform 1 0 22848 0 1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _482_
timestamp 1586547711
transform 1 0 22940 0 1 12912
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_743
timestamp 1586547711
transform 1 0 23676 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1158
timestamp 1586547711
transform 1 0 23952 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1135
timestamp 1586547711
transform 1 0 24136 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_728
timestamp 1586547711
transform 1 0 24320 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL117300x62560
timestamp 1586547711
transform 1 0 23860 0 1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _623_
timestamp 1586547711
transform 1 0 24504 0 1 12912
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL129720x62560
timestamp 1586547711
transform 1 0 26344 0 1 12912
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_627
timestamp 1586547711
transform 1 0 25792 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_727
timestamp 1586547711
transform 1 0 25976 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_732
timestamp 1586547711
transform 1 0 26160 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILL138920x62560
timestamp 1586547711
transform 1 0 28184 0 1 12912
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL135240x62560
timestamp 1586547711
transform 1 0 27448 0 1 12912
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1586547711
transform 1 0 28552 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_96
timestamp 1586547711
transform 1 0 28736 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_379
timestamp 1586547711
transform 1 0 28920 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1648
timestamp 1586547711
transform 1 0 29104 0 1 12912
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1586547711
transform 1 0 28460 0 1 12912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL144440x62560
timestamp 1586547711
transform 1 0 29288 0 1 12912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL153640x62560
timestamp 1586547711
transform 1 0 31128 0 1 12912
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL149960x62560
timestamp 1586547711
transform 1 0 30392 0 1 12912
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1586547711
transform 1 0 31404 0 1 12912
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL3220x65280
timestamp 1586547711
transform 1 0 1044 0 -1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL8740x65280
timestamp 1586547711
transform 1 0 2148 0 -1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1586547711
transform 1 0 400 0 -1 14000
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_457
timestamp 1586547711
transform 1 0 676 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1672
timestamp 1586547711
transform 1 0 860 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1586547711
transform 1 0 3252 0 -1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _911_
timestamp 1586547711
transform 1 0 3344 0 -1 14000
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_12  FILL25300x65280
timestamp 1586547711
transform 1 0 5460 0 -1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL30820x65280
timestamp 1586547711
transform 1 0 6564 0 -1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL36340x65280
timestamp 1586547711
transform 1 0 7668 0 -1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL42780x65280
timestamp 1586547711
transform 1 0 8956 0 -1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL41860x65280
timestamp 1586547711
transform 1 0 8772 0 -1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1586547711
transform 1 0 8864 0 -1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL48300x65280
timestamp 1586547711
transform 1 0 10060 0 -1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILL53820x65280
timestamp 1586547711
transform 1 0 11164 0 -1 14000
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL58420x65280
timestamp 1586547711
transform 1 0 12084 0 -1 14000
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL65320x65280
timestamp 1586547711
transform 1 0 13464 0 -1 14000
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_666
timestamp 1586547711
transform 1 0 11716 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_923
timestamp 1586547711
transform 1 0 11900 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _538_
timestamp 1586547711
transform 1 0 12820 0 -1 14000
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  FILL69000x65280
timestamp 1586547711
transform 1 0 14200 0 -1 14000
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1695
timestamp 1586547711
transform 1 0 14568 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_330
timestamp 1586547711
transform 1 0 15120 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1586547711
transform 1 0 14476 0 -1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL71760x65280
timestamp 1586547711
transform 1 0 14752 0 -1 14000
box 0 -48 368 592
use sky130_fd_sc_hd__dfrtp_4  _891_
timestamp 1586547711
transform 1 0 15304 0 -1 14000
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_8  FILL85100x65280
timestamp 1586547711
transform 1 0 17420 0 -1 14000
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILL98900x65280
timestamp 1586547711
transform 1 0 20180 0 -1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL88780x65280
timestamp 1586547711
transform 1 0 18156 0 -1 14000
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL97060x65280
timestamp 1586547711
transform 1 0 19812 0 -1 14000
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_948
timestamp 1586547711
transform 1 0 19260 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1103
timestamp 1586547711
transform 1 0 19628 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1586547711
transform 1 0 20088 0 -1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL95220x65280
timestamp 1586547711
transform 1 0 19444 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__and3_4  _583_
timestamp 1586547711
transform 1 0 18432 0 -1 14000
box 0 -48 828 592
use sky130_fd_sc_hd__fill_1  FILL104420x65280
timestamp 1586547711
transform 1 0 21284 0 -1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _493_
timestamp 1586547711
transform 1 0 21376 0 -1 14000
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_8  FILL111320x65280
timestamp 1586547711
transform 1 0 22664 0 -1 14000
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1156
timestamp 1586547711
transform 1 0 24504 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1159
timestamp 1586547711
transform 1 0 24688 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL117760x65280
timestamp 1586547711
transform 1 0 23952 0 -1 14000
box 0 -48 552 592
use sky130_fd_sc_hd__buf_4  _481_
timestamp 1586547711
transform 1 0 23400 0 -1 14000
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL132020x65280
timestamp 1586547711
transform 1 0 26804 0 -1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL122360x65280
timestamp 1586547711
transform 1 0 24872 0 -1 14000
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1204
timestamp 1586547711
transform 1 0 26436 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1220
timestamp 1586547711
transform 1 0 26620 0 -1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL126040x65280
timestamp 1586547711
transform 1 0 25608 0 -1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1586547711
transform 1 0 25700 0 -1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _479_
timestamp 1586547711
transform 1 0 25792 0 -1 14000
box 0 -48 644 592
use sky130_fd_sc_hd__fill_1  FILL139380x65280
timestamp 1586547711
transform 1 0 28276 0 -1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL137540x65280
timestamp 1586547711
transform 1 0 27908 0 -1 14000
box 0 -48 368 592
use sky130_fd_sc_hd__dfstp_4  _877_
timestamp 1586547711
transform 1 0 28368 0 -1 14000
box 0 -48 2208 592
use sky130_fd_sc_hd__decap_8  FILL150880x65280
timestamp 1586547711
transform 1 0 30576 0 -1 14000
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1586547711
transform 1 0 31312 0 -1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1586547711
transform 1 0 31404 0 -1 14000
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1586547711
transform 1 0 400 0 1 14000
box 0 -48 276 592
use sky130_fd_sc_hd__dfrtp_4  _910_
timestamp 1586547711
transform 1 0 676 0 1 14000
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_8  FILL11960x68000
timestamp 1586547711
transform 1 0 2792 0 1 14000
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1427
timestamp 1586547711
transform 1 0 3620 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1423
timestamp 1586547711
transform 1 0 3804 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_458
timestamp 1586547711
transform 1 0 3988 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL15640x68000
timestamp 1586547711
transform 1 0 3528 0 1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_619
timestamp 1586547711
transform 1 0 4172 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1413
timestamp 1586547711
transform 1 0 4356 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1415
timestamp 1586547711
transform 1 0 4540 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL21620x68000
timestamp 1586547711
transform 1 0 4724 0 1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _737_
timestamp 1586547711
transform 1 0 4816 0 1 14000
box 0 -48 460 592
use sky130_fd_sc_hd__decap_8  FILL32200x68000
timestamp 1586547711
transform 1 0 6840 0 1 14000
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1425
timestamp 1586547711
transform 1 0 5276 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1426
timestamp 1586547711
transform 1 0 5460 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_249
timestamp 1586547711
transform 1 0 6288 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1419
timestamp 1586547711
transform 1 0 6472 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1422
timestamp 1586547711
transform 1 0 6656 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1586547711
transform 1 0 6012 0 1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL26220x68000
timestamp 1586547711
transform 1 0 5644 0 1 14000
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL28520x68000
timestamp 1586547711
transform 1 0 6104 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL40480x68000
timestamp 1586547711
transform 1 0 8496 0 1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1480
timestamp 1586547711
transform 1 0 8128 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1584
timestamp 1586547711
transform 1 0 8312 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _799_
timestamp 1586547711
transform 1 0 7576 0 1 14000
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL46000x68000
timestamp 1586547711
transform 1 0 9600 0 1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL51520x68000
timestamp 1586547711
transform 1 0 10704 0 1 14000
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_862
timestamp 1586547711
transform 1 0 10980 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_665
timestamp 1586547711
transform 1 0 11164 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_653
timestamp 1586547711
transform 1 0 11348 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL61640x68000
timestamp 1586547711
transform 1 0 12728 0 1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_655
timestamp 1586547711
transform 1 0 12360 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_663
timestamp 1586547711
transform 1 0 12544 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL55660x68000
timestamp 1586547711
transform 1 0 11532 0 1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1586547711
transform 1 0 11624 0 1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _463_
timestamp 1586547711
transform 1 0 11716 0 1 14000
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  FILL67160x68000
timestamp 1586547711
transform 1 0 13832 0 1 14000
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_844
timestamp 1586547711
transform 1 0 14108 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_832
timestamp 1586547711
transform 1 0 14936 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_840
timestamp 1586547711
transform 1 0 15120 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1656
timestamp 1586547711
transform 1 0 15304 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_712
timestamp 1586547711
transform 1 0 15672 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL75440x68000
timestamp 1586547711
transform 1 0 15488 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _510_
timestamp 1586547711
transform 1 0 14292 0 1 14000
box 0 -48 644 592
use sky130_fd_sc_hd__or2_4  _475_
timestamp 1586547711
transform 1 0 15856 0 1 14000
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_667
timestamp 1586547711
transform 1 0 16500 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_708
timestamp 1586547711
transform 1 0 16684 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL86480x68000
timestamp 1586547711
transform 1 0 17696 0 1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1586547711
transform 1 0 17236 0 1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL82340x68000
timestamp 1586547711
transform 1 0 16868 0 1 14000
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILL84640x68000
timestamp 1586547711
transform 1 0 17328 0 1 14000
box 0 -48 368 592
use sky130_fd_sc_hd__buf_4  _476_
timestamp 1586547711
transform 1 0 17788 0 1 14000
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_713
timestamp 1586547711
transform 1 0 18340 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_714
timestamp 1586547711
transform 1 0 18524 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_334
timestamp 1586547711
transform 1 0 18708 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_55
timestamp 1586547711
transform 1 0 18892 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _548_
timestamp 1586547711
transform 1 0 19076 0 1 14000
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL99820x68000
timestamp 1586547711
transform 1 0 20364 0 1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL105340x68000
timestamp 1586547711
transform 1 0 21468 0 1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL119600x68000
timestamp 1586547711
transform 1 0 24320 0 1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL110860x68000
timestamp 1586547711
transform 1 0 22572 0 1 14000
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_737
timestamp 1586547711
transform 1 0 23032 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_719
timestamp 1586547711
transform 1 0 23768 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_733
timestamp 1586547711
transform 1 0 23952 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1133
timestamp 1586547711
transform 1 0 24136 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL112700x68000
timestamp 1586547711
transform 1 0 22940 0 1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1586547711
transform 1 0 22848 0 1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _480_
timestamp 1586547711
transform 1 0 23216 0 1 14000
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1203
timestamp 1586547711
transform 1 0 25792 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1180
timestamp 1586547711
transform 1 0 25976 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_730
timestamp 1586547711
transform 1 0 26160 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_146
timestamp 1586547711
transform 1 0 26344 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL130640x68000
timestamp 1586547711
transform 1 0 26528 0 1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL125120x68000
timestamp 1586547711
transform 1 0 25424 0 1 14000
box 0 -48 368 592
use sky130_fd_sc_hd__and2_4  _646_
timestamp 1586547711
transform 1 0 26620 0 1 14000
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL140760x68000
timestamp 1586547711
transform 1 0 28552 0 1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL136160x68000
timestamp 1586547711
transform 1 0 27632 0 1 14000
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_143
timestamp 1586547711
transform 1 0 27264 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_724
timestamp 1586547711
transform 1 0 27448 0 1 14000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL139840x68000
timestamp 1586547711
transform 1 0 28368 0 1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1586547711
transform 1 0 28460 0 1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL146280x68000
timestamp 1586547711
transform 1 0 29656 0 1 14000
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL154560x68000
timestamp 1586547711
transform 1 0 31312 0 1 14000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL151800x68000
timestamp 1586547711
transform 1 0 30760 0 1 14000
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1586547711
transform 1 0 31404 0 1 14000
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL3220x70720
timestamp 1586547711
transform 1 0 1044 0 -1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1586547711
transform 1 0 400 0 1 15088
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL1380x73440
timestamp 1586547711
transform 1 0 676 0 1 15088
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1586547711
transform 1 0 400 0 -1 15088
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL3680x73440
timestamp 1586547711
transform 1 0 1136 0 1 15088
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_186
timestamp 1586547711
transform 1 0 952 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_246
timestamp 1586547711
transform 1 0 676 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1506
timestamp 1586547711
transform 1 0 860 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL8740x70720
timestamp 1586547711
transform 1 0 2148 0 -1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_245
timestamp 1586547711
transform 1 0 1964 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1385
timestamp 1586547711
transform 1 0 2148 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL7360x73440
timestamp 1586547711
transform 1 0 1872 0 1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL9660x73440
timestamp 1586547711
transform 1 0 2332 0 1 15088
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1414
timestamp 1586547711
transform 1 0 2792 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1407
timestamp 1586547711
transform 1 0 2976 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1408
timestamp 1586547711
transform 1 0 3344 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL11500x73440
timestamp 1586547711
transform 1 0 2700 0 1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1586547711
transform 1 0 3252 0 -1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL15640x70720
timestamp 1586547711
transform 1 0 3528 0 -1 15088
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _732_
timestamp 1586547711
transform 1 0 3160 0 1 15088
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_759
timestamp 1586547711
transform 1 0 3804 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1389
timestamp 1586547711
transform 1 0 3988 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1406
timestamp 1586547711
transform 1 0 4172 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1403
timestamp 1586547711
transform 1 0 4448 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL19780x73440
timestamp 1586547711
transform 1 0 4356 0 1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL17480x70720
timestamp 1586547711
transform 1 0 3896 0 -1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _731_
timestamp 1586547711
transform 1 0 4632 0 1 15088
box 0 -48 644 592
use sky130_fd_sc_hd__a32o_4  _738_
timestamp 1586547711
transform 1 0 3988 0 -1 15088
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA_248
timestamp 1586547711
transform 1 0 5276 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_250
timestamp 1586547711
transform 1 0 5460 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1424
timestamp 1586547711
transform 1 0 5552 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_591
timestamp 1586547711
transform 1 0 5644 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_618
timestamp 1586547711
transform 1 0 5828 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1420
timestamp 1586547711
transform 1 0 6104 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1586547711
transform 1 0 6012 0 1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL29440x73440
timestamp 1586547711
transform 1 0 6288 0 1 15088
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILL26680x70720
timestamp 1586547711
transform 1 0 5736 0 -1 15088
box 0 -48 552 592
use sky130_fd_sc_hd__or2_4  _735_
timestamp 1586547711
transform 1 0 6288 0 -1 15088
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL32660x70720
timestamp 1586547711
transform 1 0 6932 0 -1 15088
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1432
timestamp 1586547711
transform 1 0 6748 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_588
timestamp 1586547711
transform 1 0 6932 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL31280x73440
timestamp 1586547711
transform 1 0 6656 0 1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_253
timestamp 1586547711
transform 1 0 7116 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_247
timestamp 1586547711
transform 1 0 7300 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_251
timestamp 1586547711
transform 1 0 7484 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_254
timestamp 1586547711
transform 1 0 7668 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_460
timestamp 1586547711
transform 1 0 7852 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1430
timestamp 1586547711
transform 1 0 8036 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL42780x73440
timestamp 1586547711
transform 1 0 8956 0 1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL42780x70720
timestamp 1586547711
transform 1 0 8956 0 -1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL41860x70720
timestamp 1586547711
transform 1 0 8772 0 -1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1586547711
transform 1 0 8864 0 -1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL39100x70720
timestamp 1586547711
transform 1 0 8220 0 -1 15088
box 0 -48 552 592
use sky130_fd_sc_hd__o22a_4  _741_
timestamp 1586547711
transform 1 0 7668 0 1 15088
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL48300x70720
timestamp 1586547711
transform 1 0 10060 0 -1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILL48300x73440
timestamp 1586547711
transform 1 0 10060 0 1 15088
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_664
timestamp 1586547711
transform 1 0 10704 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_828
timestamp 1586547711
transform 1 0 10888 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_831
timestamp 1586547711
transform 1 0 11256 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_829
timestamp 1586547711
transform 1 0 11440 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL51060x73440
timestamp 1586547711
transform 1 0 10612 0 1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL53360x73440
timestamp 1586547711
transform 1 0 11072 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL53820x70720
timestamp 1586547711
transform 1 0 11164 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _518_
timestamp 1586547711
transform 1 0 11348 0 -1 15088
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL62560x73440
timestamp 1586547711
transform 1 0 12912 0 1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL58880x70720
timestamp 1586547711
transform 1 0 12176 0 -1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL64400x70720
timestamp 1586547711
transform 1 0 13280 0 -1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_652
timestamp 1586547711
transform 1 0 12360 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_656
timestamp 1586547711
transform 1 0 12544 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_830
timestamp 1586547711
transform 1 0 12728 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_972
timestamp 1586547711
transform 1 0 11992 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1586547711
transform 1 0 11624 0 1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _507_
timestamp 1586547711
transform 1 0 11716 0 1 15088
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1673
timestamp 1586547711
transform 1 0 14568 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1696
timestamp 1586547711
transform 1 0 14752 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL69920x70720
timestamp 1586547711
transform 1 0 14384 0 -1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1586547711
transform 1 0 14476 0 -1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_4  _CTS_buf_1_32 ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 14016 0 1 15088
box 0 -48 552 592
use sky130_fd_sc_hd__clkbuf_4  _CTS_buf_1_16
timestamp 1586547711
transform 1 0 14568 0 -1 15088
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL73600x70720
timestamp 1586547711
transform 1 0 15120 0 -1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_835
timestamp 1586547711
transform 1 0 15488 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_931
timestamp 1586547711
transform 1 0 15672 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_934
timestamp 1586547711
transform 1 0 15856 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL72680x73440
timestamp 1586547711
transform 1 0 14936 0 1 15088
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL78200x73440
timestamp 1586547711
transform 1 0 16040 0 1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL84640x73440
timestamp 1586547711
transform 1 0 17328 0 1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL79120x70720
timestamp 1586547711
transform 1 0 16224 0 -1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL84640x70720
timestamp 1586547711
transform 1 0 17328 0 -1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL83720x73440
timestamp 1586547711
transform 1 0 17144 0 1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1586547711
transform 1 0 17236 0 1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_57
timestamp 1586547711
transform 1 0 18432 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1586547711
transform 1 0 18616 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1625
timestamp 1586547711
transform 1 0 18800 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_792
timestamp 1586547711
transform 1 0 19076 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL92920x70720
timestamp 1586547711
transform 1 0 18984 0 -1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL90160x70720
timestamp 1586547711
transform 1 0 18432 0 -1 15088
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL98900x70720
timestamp 1586547711
transform 1 0 20180 0 -1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_944
timestamp 1586547711
transform 1 0 19260 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL97980x70720
timestamp 1586547711
transform 1 0 19996 0 -1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1586547711
transform 1 0 20088 0 -1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL95220x70720
timestamp 1586547711
transform 1 0 19444 0 -1 15088
box 0 -48 552 592
use sky130_fd_sc_hd__dfstp_4  _855_
timestamp 1586547711
transform 1 0 18800 0 1 15088
box 0 -48 2208 592
use sky130_fd_sc_hd__decap_12  FILL104420x70720
timestamp 1586547711
transform 1 0 21284 0 -1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL103040x73440
timestamp 1586547711
transform 1 0 21008 0 1 15088
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL109940x70720
timestamp 1586547711
transform 1 0 22388 0 -1 15088
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1586547711
transform 1 0 21836 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_153
timestamp 1586547711
transform 1 0 22020 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_389
timestamp 1586547711
transform 1 0 22204 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1628
timestamp 1586547711
transform 1 0 22388 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL106720x73440
timestamp 1586547711
transform 1 0 21744 0 1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILL110860x73440
timestamp 1586547711
transform 1 0 22572 0 1 15088
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL113620x70720
timestamp 1586547711
transform 1 0 23124 0 -1 15088
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL112700x73440
timestamp 1586547711
transform 1 0 22940 0 1 15088
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1586547711
transform 1 0 22848 0 1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _611_
timestamp 1586547711
transform 1 0 23400 0 -1 15088
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL120060x70720
timestamp 1586547711
transform 1 0 24412 0 -1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL117760x70720
timestamp 1586547711
transform 1 0 23952 0 -1 15088
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_815
timestamp 1586547711
transform 1 0 23676 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_396
timestamp 1586547711
transform 1 0 23860 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_139
timestamp 1586547711
transform 1 0 24044 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_746
timestamp 1586547711
transform 1 0 24228 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _502_
timestamp 1586547711
transform 1 0 24228 0 1 15088
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1233
timestamp 1586547711
transform 1 0 25884 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1181
timestamp 1586547711
transform 1 0 26068 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1137
timestamp 1586547711
transform 1 0 26252 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1586547711
transform 1 0 25700 0 -1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL125580x73440
timestamp 1586547711
transform 1 0 25516 0 1 15088
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILL126960x70720
timestamp 1586547711
transform 1 0 25792 0 -1 15088
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILL125580x70720
timestamp 1586547711
transform 1 0 25516 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__a211o_4  _654_
timestamp 1586547711
transform 1 0 26436 0 1 15088
box 0 -48 1288 592
use sky130_fd_sc_hd__a211o_4  _639_
timestamp 1586547711
transform 1 0 26344 0 -1 15088
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_8  FILL137080x70720
timestamp 1586547711
transform 1 0 27816 0 -1 15088
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1136
timestamp 1586547711
transform 1 0 27724 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1177
timestamp 1586547711
transform 1 0 27908 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1222
timestamp 1586547711
transform 1 0 27632 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL141680x70720
timestamp 1586547711
transform 1 0 28736 0 -1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1219
timestamp 1586547711
transform 1 0 28092 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1221
timestamp 1586547711
transform 1 0 28276 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1232
timestamp 1586547711
transform 1 0 28552 0 -1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1586547711
transform 1 0 28460 0 1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _653_
timestamp 1586547711
transform 1 0 28552 0 1 15088
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL145820x73440
timestamp 1586547711
transform 1 0 29564 0 1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL147200x70720
timestamp 1586547711
transform 1 0 29840 0 -1 15088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL151340x73440
timestamp 1586547711
transform 1 0 30668 0 1 15088
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_140
timestamp 1586547711
transform 1 0 29196 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_725
timestamp 1586547711
transform 1 0 29380 0 1 15088
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1586547711
transform 1 0 31312 0 -1 15088
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL152720x70720
timestamp 1586547711
transform 1 0 30944 0 -1 15088
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1586547711
transform 1 0 31404 0 1 15088
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1586547711
transform 1 0 31404 0 -1 15088
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1586547711
transform 1 0 400 0 -1 16176
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL1380x76160
timestamp 1586547711
transform 1 0 676 0 -1 16176
box 0 -48 276 592
use sky130_fd_sc_hd__conb_1  _845_
timestamp 1586547711
transform 1 0 952 0 -1 16176
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1387
timestamp 1586547711
transform 1 0 1320 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1395
timestamp 1586547711
transform 1 0 1504 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1398
timestamp 1586547711
transform 1 0 1688 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL4140x76160
timestamp 1586547711
transform 1 0 1228 0 -1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL7360x76160
timestamp 1586547711
transform 1 0 1872 0 -1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL10580x76160
timestamp 1586547711
transform 1 0 2516 0 -1 16176
box 0 -48 736 592
use sky130_fd_sc_hd__buf_4  _721_
timestamp 1586547711
transform 1 0 1964 0 -1 16176
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1412
timestamp 1586547711
transform 1 0 4632 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL20700x76160
timestamp 1586547711
transform 1 0 4540 0 -1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1586547711
transform 1 0 3252 0 -1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL22080x76160
timestamp 1586547711
transform 1 0 4816 0 -1 16176
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILL17940x76160
timestamp 1586547711
transform 1 0 3988 0 -1 16176
box 0 -48 552 592
use sky130_fd_sc_hd__or2_4  _728_
timestamp 1586547711
transform 1 0 3344 0 -1 16176
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL30820x76160
timestamp 1586547711
transform 1 0 6564 0 -1 16176
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL23920x76160
timestamp 1586547711
transform 1 0 5184 0 -1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__a211o_4  _736_
timestamp 1586547711
transform 1 0 5276 0 -1 16176
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_3  FILL38640x76160
timestamp 1586547711
transform 1 0 8128 0 -1 16176
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL40940x76160
timestamp 1586547711
transform 1 0 8588 0 -1 16176
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1675
timestamp 1586547711
transform 1 0 8404 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_607
timestamp 1586547711
transform 1 0 8956 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1421
timestamp 1586547711
transform 1 0 9140 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1586547711
transform 1 0 8864 0 -1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__nor2_4  _444_
timestamp 1586547711
transform 1 0 7300 0 -1 16176
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  FILL50140x76160
timestamp 1586547711
transform 1 0 10428 0 -1 16176
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL46460x76160
timestamp 1586547711
transform 1 0 9692 0 -1 16176
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL53820x76160
timestamp 1586547711
transform 1 0 11164 0 -1 16176
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1429
timestamp 1586547711
transform 1 0 9324 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1431
timestamp 1586547711
transform 1 0 9508 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _506_
timestamp 1586547711
transform 1 0 10704 0 -1 16176
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL60720x76160
timestamp 1586547711
transform 1 0 12544 0 -1 16176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL66240x76160
timestamp 1586547711
transform 1 0 13648 0 -1 16176
box 0 -48 736 592
use sky130_fd_sc_hd__or2_4  _555_
timestamp 1586547711
transform 1 0 11900 0 -1 16176
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL70840x76160
timestamp 1586547711
transform 1 0 14568 0 -1 16176
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL69920x76160
timestamp 1586547711
transform 1 0 14384 0 -1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1586547711
transform 1 0 14476 0 -1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL74520x76160
timestamp 1586547711
transform 1 0 15304 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _544_
timestamp 1586547711
transform 1 0 15488 0 -1 16176
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL78660x76160
timestamp 1586547711
transform 1 0 16132 0 -1 16176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL84180x76160
timestamp 1586547711
transform 1 0 17236 0 -1 16176
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_926
timestamp 1586547711
transform 1 0 18064 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL87860x76160
timestamp 1586547711
transform 1 0 17972 0 -1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_946
timestamp 1586547711
transform 1 0 18248 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_950
timestamp 1586547711
transform 1 0 18432 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_335
timestamp 1586547711
transform 1 0 18800 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_939
timestamp 1586547711
transform 1 0 18984 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_980
timestamp 1586547711
transform 1 0 19168 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL91080x76160
timestamp 1586547711
transform 1 0 18616 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL98900x76160
timestamp 1586547711
transform 1 0 20180 0 -1 16176
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1057
timestamp 1586547711
transform 1 0 19352 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1586547711
transform 1 0 20088 0 -1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL95680x76160
timestamp 1586547711
transform 1 0 19536 0 -1 16176
box 0 -48 552 592
use sky130_fd_sc_hd__decap_6  FILL104420x76160
timestamp 1586547711
transform 1 0 21284 0 -1 16176
box 0 -48 552 592
use sky130_fd_sc_hd__dfstp_4  _858_
timestamp 1586547711
transform 1 0 21836 0 -1 16176
box 0 -48 2208 592
use sky130_fd_sc_hd__decap_12  FILL120060x76160
timestamp 1586547711
transform 1 0 24412 0 -1 16176
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_819
timestamp 1586547711
transform 1 0 24044 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_735
timestamp 1586547711
transform 1 0 24228 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL132020x76160
timestamp 1586547711
transform 1 0 26804 0 -1 16176
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1231
timestamp 1586547711
transform 1 0 26436 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1234
timestamp 1586547711
transform 1 0 26620 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL129720x76160
timestamp 1586547711
transform 1 0 26344 0 -1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1586547711
transform 1 0 25700 0 -1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL126960x76160
timestamp 1586547711
transform 1 0 25792 0 -1 16176
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILL125580x76160
timestamp 1586547711
transform 1 0 25516 0 -1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL142140x76160
timestamp 1586547711
transform 1 0 28828 0 -1 16176
box 0 -48 1104 592
use sky130_fd_sc_hd__a211o_4  _647_
timestamp 1586547711
transform 1 0 27540 0 -1 16176
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL147660x76160
timestamp 1586547711
transform 1 0 29932 0 -1 16176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL153180x76160
timestamp 1586547711
transform 1 0 31036 0 -1 16176
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1586547711
transform 1 0 31312 0 -1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1586547711
transform 1 0 31404 0 -1 16176
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1586547711
transform 1 0 400 0 1 16176
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1287
timestamp 1586547711
transform 1 0 768 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_456
timestamp 1586547711
transform 1 0 952 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL1380x78880
timestamp 1586547711
transform 1 0 676 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__a32o_4  _730_
timestamp 1586547711
transform 1 0 1136 0 1 16176
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1399
timestamp 1586547711
transform 1 0 2700 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1409
timestamp 1586547711
transform 1 0 2884 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1405
timestamp 1586547711
transform 1 0 3068 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1402
timestamp 1586547711
transform 1 0 3252 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _727_
timestamp 1586547711
transform 1 0 3436 0 1 16176
box 0 -48 460 592
use sky130_fd_sc_hd__diode_2  ANTENNA_617
timestamp 1586547711
transform 1 0 3896 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1388
timestamp 1586547711
transform 1 0 4080 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1401
timestamp 1586547711
transform 1 0 4264 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1410
timestamp 1586547711
transform 1 0 4448 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL21160x78880
timestamp 1586547711
transform 1 0 4632 0 1 16176
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_310
timestamp 1586547711
transform 1 0 5184 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_582
timestamp 1586547711
transform 1 0 5368 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1273
timestamp 1586547711
transform 1 0 5552 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1433
timestamp 1586547711
transform 1 0 5736 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL27600x78880
timestamp 1586547711
transform 1 0 5920 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1586547711
transform 1 0 6012 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL28520x78880
timestamp 1586547711
transform 1 0 6104 0 1 16176
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1418
timestamp 1586547711
transform 1 0 6564 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL30360x78880
timestamp 1586547711
transform 1 0 6472 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_244
timestamp 1586547711
transform 1 0 6748 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _734_
timestamp 1586547711
transform 1 0 6932 0 1 16176
box 0 -48 460 592
use sky130_fd_sc_hd__diode_2  ANTENNA_589
timestamp 1586547711
transform 1 0 7392 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_592
timestamp 1586547711
transform 1 0 7576 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1417
timestamp 1586547711
transform 1 0 7760 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_461
timestamp 1586547711
transform 1 0 8036 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_255
timestamp 1586547711
transform 1 0 8220 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL37720x78880
timestamp 1586547711
transform 1 0 7944 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _912_
timestamp 1586547711
transform 1 0 8404 0 1 16176
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_12  FILL50600x78880
timestamp 1586547711
transform 1 0 10520 0 1 16176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL60720x78880
timestamp 1586547711
transform 1 0 12544 0 1 16176
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_651
timestamp 1586547711
transform 1 0 12176 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_654
timestamp 1586547711
transform 1 0 12360 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1586547711
transform 1 0 11624 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL66240x78880
timestamp 1586547711
transform 1 0 13648 0 1 16176
box 0 -48 552 592
use sky130_fd_sc_hd__inv_4  _460_
timestamp 1586547711
transform 1 0 11716 0 1 16176
box 0 -48 460 592
use sky130_fd_sc_hd__diode_2  ANTENNA_973
timestamp 1586547711
transform 1 0 14752 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_974
timestamp 1586547711
transform 1 0 14936 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1639
timestamp 1586547711
transform 1 0 15120 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1694
timestamp 1586547711
transform 1 0 15304 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL77280x78880
timestamp 1586547711
transform 1 0 15856 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL75440x78880
timestamp 1586547711
transform 1 0 15488 0 1 16176
box 0 -48 368 592
use sky130_fd_sc_hd__buf_4  _556_
timestamp 1586547711
transform 1 0 14200 0 1 16176
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_913
timestamp 1586547711
transform 1 0 15948 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_975
timestamp 1586547711
transform 1 0 16132 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_979
timestamp 1586547711
transform 1 0 16316 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL80500x78880
timestamp 1586547711
transform 1 0 16500 0 1 16176
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_936
timestamp 1586547711
transform 1 0 17052 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL84640x78880
timestamp 1586547711
transform 1 0 17328 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1586547711
transform 1 0 17236 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _547_
timestamp 1586547711
transform 1 0 17420 0 1 16176
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_49
timestamp 1586547711
transform 1 0 18064 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL87860x78880
timestamp 1586547711
transform 1 0 17972 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_408
timestamp 1586547711
transform 1 0 18248 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_56
timestamp 1586547711
transform 1 0 18524 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_52
timestamp 1586547711
transform 1 0 20180 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL90160x78880
timestamp 1586547711
transform 1 0 18432 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL97980x78880
timestamp 1586547711
transform 1 0 19996 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__a211o_4  _584_
timestamp 1586547711
transform 1 0 18708 0 1 16176
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL103500x78880
timestamp 1586547711
transform 1 0 21100 0 1 16176
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_404
timestamp 1586547711
transform 1 0 20364 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_783
timestamp 1586547711
transform 1 0 20548 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_945
timestamp 1586547711
transform 1 0 20732 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_949
timestamp 1586547711
transform 1 0 20916 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_748
timestamp 1586547711
transform 1 0 22296 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_941
timestamp 1586547711
transform 1 0 22480 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL109020x78880
timestamp 1586547711
transform 1 0 22204 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1132
timestamp 1586547711
transform 1 0 22664 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1140
timestamp 1586547711
transform 1 0 22940 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1141
timestamp 1586547711
transform 1 0 23124 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_747
timestamp 1586547711
transform 1 0 23400 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_398
timestamp 1586547711
transform 1 0 23584 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_136
timestamp 1586547711
transform 1 0 23768 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL114540x78880
timestamp 1586547711
transform 1 0 23308 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1586547711
transform 1 0 22848 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _504_
timestamp 1586547711
transform 1 0 23952 0 1 16176
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1139
timestamp 1586547711
transform 1 0 25608 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1134
timestamp 1586547711
transform 1 0 25792 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_152
timestamp 1586547711
transform 1 0 26804 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL124200x78880
timestamp 1586547711
transform 1 0 25240 0 1 16176
box 0 -48 368 592
use sky130_fd_sc_hd__nor2_4  _612_
timestamp 1586547711
transform 1 0 25976 0 1 16176
box 0 -48 828 592
use sky130_fd_sc_hd__decap_12  FILL140760x78880
timestamp 1586547711
transform 1 0 28552 0 1 16176
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1172
timestamp 1586547711
transform 1 0 27632 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1245
timestamp 1586547711
transform 1 0 27816 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1249
timestamp 1586547711
transform 1 0 28000 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1250
timestamp 1586547711
transform 1 0 28184 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL135700x78880
timestamp 1586547711
transform 1 0 27540 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL139840x78880
timestamp 1586547711
transform 1 0 28368 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1586547711
transform 1 0 28460 0 1 16176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL132940x78880
timestamp 1586547711
transform 1 0 26988 0 1 16176
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL150420x78880
timestamp 1586547711
transform 1 0 30484 0 1 16176
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_48
timestamp 1586547711
transform 1 0 30116 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_500
timestamp 1586547711
transform 1 0 30300 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL154100x78880
timestamp 1586547711
transform 1 0 31220 0 1 16176
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _417_
timestamp 1586547711
transform 1 0 29656 0 1 16176
box 0 -48 460 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1586547711
transform 1 0 31404 0 1 16176
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL8740x81600
timestamp 1586547711
transform 1 0 2148 0 -1 17264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1586547711
transform 1 0 400 0 -1 17264
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL1380x81600
timestamp 1586547711
transform 1 0 676 0 -1 17264
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1411
timestamp 1586547711
transform 1 0 952 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1397
timestamp 1586547711
transform 1 0 1136 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__nand2_4  _725_ ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 1320 0 -1 17264
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1272
timestamp 1586547711
transform 1 0 4816 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1586547711
transform 1 0 3252 0 -1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL20240x81600
timestamp 1586547711
transform 1 0 4448 0 -1 17264
box 0 -48 368 592
use sky130_fd_sc_hd__o21a_4  _729_ ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 3344 0 -1 17264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL28060x81600
timestamp 1586547711
transform 1 0 6012 0 -1 17264
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILL23000x81600
timestamp 1586547711
transform 1 0 5000 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _445_
timestamp 1586547711
transform 1 0 6748 0 -1 17264
box 0 -48 644 592
use sky130_fd_sc_hd__or3_4  _742_ ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 5184 0 -1 17264
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  FILL38640x81600
timestamp 1586547711
transform 1 0 8128 0 -1 17264
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL40940x81600
timestamp 1586547711
transform 1 0 8588 0 -1 17264
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL34960x81600
timestamp 1586547711
transform 1 0 7392 0 -1 17264
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1515
timestamp 1586547711
transform 1 0 8404 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1586547711
transform 1 0 8864 0 -1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__a21oi_4  _740_ ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 8956 0 -1 17264
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_12  FILL48760x81600
timestamp 1586547711
transform 1 0 10152 0 -1 17264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL54280x81600
timestamp 1586547711
transform 1 0 11256 0 -1 17264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL64860x81600
timestamp 1586547711
transform 1 0 13372 0 -1 17264
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_839
timestamp 1586547711
transform 1 0 12820 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_696
timestamp 1586547711
transform 1 0 13004 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_838
timestamp 1586547711
transform 1 0 13188 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL61640x81600
timestamp 1586547711
transform 1 0 12728 0 -1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL59800x81600
timestamp 1586547711
transform 1 0 12360 0 -1 17264
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILL73600x81600
timestamp 1586547711
transform 1 0 15120 0 -1 17264
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL77280x81600
timestamp 1586547711
transform 1 0 15856 0 -1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1586547711
transform 1 0 14476 0 -1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_4  _CTS_buf_1_0
timestamp 1586547711
transform 1 0 14568 0 -1 17264
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_947
timestamp 1586547711
transform 1 0 17420 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1623
timestamp 1586547711
transform 1 0 17788 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL84640x81600
timestamp 1586547711
transform 1 0 17328 0 -1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL87860x81600
timestamp 1586547711
transform 1 0 17972 0 -1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL81880x81600
timestamp 1586547711
transform 1 0 16776 0 -1 17264
box 0 -48 552 592
use sky130_fd_sc_hd__o22a_4  _550_
timestamp 1586547711
transform 1 0 18064 0 -1 17264
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILL86020x81600
timestamp 1586547711
transform 1 0 17604 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _557_
timestamp 1586547711
transform 1 0 15948 0 -1 17264
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1056
timestamp 1586547711
transform 1 0 19352 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1586547711
transform 1 0 20088 0 -1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL95680x81600
timestamp 1586547711
transform 1 0 19536 0 -1 17264
box 0 -48 552 592
use sky130_fd_sc_hd__o22a_4  _549_
timestamp 1586547711
transform 1 0 20180 0 -1 17264
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_8  FILL105340x81600
timestamp 1586547711
transform 1 0 21468 0 -1 17264
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL109020x81600
timestamp 1586547711
transform 1 0 22204 0 -1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__a211o_4  _613_
timestamp 1586547711
transform 1 0 22296 0 -1 17264
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL118680x81600
timestamp 1586547711
transform 1 0 24136 0 -1 17264
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_736
timestamp 1586547711
transform 1 0 23952 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL115920x81600
timestamp 1586547711
transform 1 0 23584 0 -1 17264
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL126960x81600
timestamp 1586547711
transform 1 0 25792 0 -1 17264
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1244
timestamp 1586547711
transform 1 0 26896 0 -1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL126040x81600
timestamp 1586547711
transform 1 0 25608 0 -1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1586547711
transform 1 0 25700 0 -1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL124200x81600
timestamp 1586547711
transform 1 0 25240 0 -1 17264
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL140300x81600
timestamp 1586547711
transform 1 0 28460 0 -1 17264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILL133400x81600
timestamp 1586547711
transform 1 0 27080 0 -1 17264
box 0 -48 552 592
use sky130_fd_sc_hd__and3_4  _663_
timestamp 1586547711
transform 1 0 27632 0 -1 17264
box 0 -48 828 592
use sky130_fd_sc_hd__decap_12  FILL145820x81600
timestamp 1586547711
transform 1 0 29564 0 -1 17264
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL154100x81600
timestamp 1586547711
transform 1 0 31220 0 -1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1586547711
transform 1 0 31312 0 -1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL151340x81600
timestamp 1586547711
transform 1 0 30668 0 -1 17264
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1586547711
transform 1 0 31404 0 -1 17264
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1586547711
transform 1 0 400 0 1 17264
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL1380x84320
timestamp 1586547711
transform 1 0 676 0 1 17264
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1396
timestamp 1586547711
transform 1 0 1412 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1386
timestamp 1586547711
transform 1 0 2240 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1394
timestamp 1586547711
transform 1 0 2424 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL11040x84320
timestamp 1586547711
transform 1 0 2608 0 1 17264
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _724_
timestamp 1586547711
transform 1 0 1596 0 1 17264
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1392
timestamp 1586547711
transform 1 0 3436 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1393
timestamp 1586547711
transform 1 0 3620 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1391
timestamp 1586547711
transform 1 0 4172 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_614
timestamp 1586547711
transform 1 0 4356 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_590
timestamp 1586547711
transform 1 0 4540 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL17020x84320
timestamp 1586547711
transform 1 0 3804 0 1 17264
box 0 -48 368 592
use sky130_fd_sc_hd__buf_4  _452_
timestamp 1586547711
transform 1 0 4724 0 1 17264
box 0 -48 552 592
use sky130_fd_sc_hd__inv_4  _723_
timestamp 1586547711
transform 1 0 2976 0 1 17264
box 0 -48 460 592
use sky130_fd_sc_hd__diode_2  ANTENNA_308
timestamp 1586547711
transform 1 0 5276 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_565
timestamp 1586547711
transform 1 0 5460 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_581
timestamp 1586547711
transform 1 0 5644 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL27140x84320
timestamp 1586547711
transform 1 0 5828 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILL28520x84320
timestamp 1586547711
transform 1 0 6104 0 1 17264
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1586547711
transform 1 0 6012 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_566
timestamp 1586547711
transform 1 0 6380 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_576
timestamp 1586547711
transform 1 0 6564 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_643
timestamp 1586547711
transform 1 0 6748 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1390
timestamp 1586547711
transform 1 0 6932 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL34500x84320
timestamp 1586547711
transform 1 0 7300 0 1 17264
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1416
timestamp 1586547711
transform 1 0 7116 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1428
timestamp 1586547711
transform 1 0 8128 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_309
timestamp 1586547711
transform 1 0 8956 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1404
timestamp 1586547711
transform 1 0 9140 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL38180x84320
timestamp 1586547711
transform 1 0 8036 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _739_
timestamp 1586547711
transform 1 0 8312 0 1 17264
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL44620x84320
timestamp 1586547711
transform 1 0 9324 0 1 17264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL50140x84320
timestamp 1586547711
transform 1 0 10428 0 1 17264
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_930
timestamp 1586547711
transform 1 0 12268 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_837
timestamp 1586547711
transform 1 0 12452 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_695
timestamp 1586547711
transform 1 0 12636 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_682
timestamp 1586547711
transform 1 0 12820 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL55660x84320
timestamp 1586547711
transform 1 0 11532 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1586547711
transform 1 0 11624 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL56580x84320
timestamp 1586547711
transform 1 0 11716 0 1 17264
box 0 -48 552 592
use sky130_fd_sc_hd__or3_4  _543_
timestamp 1586547711
transform 1 0 13004 0 1 17264
box 0 -48 828 592
use sky130_fd_sc_hd__decap_8  FILL76820x84320
timestamp 1586547711
transform 1 0 15764 0 1 17264
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_686
timestamp 1586547711
transform 1 0 13832 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_707
timestamp 1586547711
transform 1 0 14016 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_705
timestamp 1586547711
transform 1 0 14200 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_704
timestamp 1586547711
transform 1 0 14384 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_683
timestamp 1586547711
transform 1 0 15212 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_685
timestamp 1586547711
transform 1 0 15396 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_911
timestamp 1586547711
transform 1 0 15580 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _537_
timestamp 1586547711
transform 1 0 14568 0 1 17264
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_843
timestamp 1586547711
transform 1 0 16592 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_976
timestamp 1586547711
transform 1 0 16776 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1075
timestamp 1586547711
transform 1 0 16960 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL80500x84320
timestamp 1586547711
transform 1 0 16500 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_51
timestamp 1586547711
transform 1 0 17420 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1586547711
transform 1 0 17604 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL83720x84320
timestamp 1586547711
transform 1 0 17144 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL84640x84320
timestamp 1586547711
transform 1 0 17328 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1586547711
transform 1 0 17236 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__dfstp_4  _853_
timestamp 1586547711
transform 1 0 17788 0 1 17264
box 0 -48 2208 592
use sky130_fd_sc_hd__diode_2  ANTENNA_943
timestamp 1586547711
transform 1 0 19996 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_405
timestamp 1586547711
transform 1 0 20180 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL108100x84320
timestamp 1586547711
transform 1 0 22020 0 1 17264
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1586547711
transform 1 0 20364 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_54
timestamp 1586547711
transform 1 0 20548 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_629
timestamp 1586547711
transform 1 0 21468 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_938
timestamp 1586547711
transform 1 0 21652 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1624
timestamp 1586547711
transform 1 0 21836 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL101660x84320
timestamp 1586547711
transform 1 0 20732 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _546_
timestamp 1586547711
transform 1 0 20824 0 1 17264
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1632
timestamp 1586547711
transform 1 0 23400 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_141
timestamp 1586547711
transform 1 0 23584 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1586547711
transform 1 0 23768 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL111780x84320
timestamp 1586547711
transform 1 0 22756 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL114540x84320
timestamp 1586547711
transform 1 0 23308 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1586547711
transform 1 0 22848 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL112700x84320
timestamp 1586547711
transform 1 0 22940 0 1 17264
box 0 -48 368 592
use sky130_fd_sc_hd__dfstp_4  _862_
timestamp 1586547711
transform 1 0 23952 0 1 17264
box 0 -48 2208 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1179
timestamp 1586547711
transform 1 0 26252 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1176
timestamp 1586547711
transform 1 0 26436 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1077
timestamp 1586547711
transform 1 0 26620 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL128800x84320
timestamp 1586547711
transform 1 0 26160 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL132020x84320
timestamp 1586547711
transform 1 0 26804 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _660_
timestamp 1586547711
transform 1 0 26896 0 1 17264
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_137
timestamp 1586547711
transform 1 0 27540 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1138
timestamp 1586547711
transform 1 0 27724 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_501
timestamp 1586547711
transform 1 0 28000 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL137540x84320
timestamp 1586547711
transform 1 0 27908 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL142600x84320
timestamp 1586547711
transform 1 0 28920 0 1 17264
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1358
timestamp 1586547711
transform 1 0 28184 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1481
timestamp 1586547711
transform 1 0 28552 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1618
timestamp 1586547711
transform 1 0 28736 0 1 17264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL139840x84320
timestamp 1586547711
transform 1 0 28368 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1586547711
transform 1 0 28460 0 1 17264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL148120x84320
timestamp 1586547711
transform 1 0 30024 0 1 17264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL153640x84320
timestamp 1586547711
transform 1 0 31128 0 1 17264
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1586547711
transform 1 0 31404 0 1 17264
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL1380x87040
timestamp 1586547711
transform 1 0 676 0 -1 18352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL6900x87040
timestamp 1586547711
transform 1 0 1780 0 -1 18352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1586547711
transform 1 0 400 0 -1 18352
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL14720x87040
timestamp 1586547711
transform 1 0 3344 0 -1 18352
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1586547711
transform 1 0 3252 0 -1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL12420x87040
timestamp 1586547711
transform 1 0 2884 0 -1 18352
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILL20240x87040
timestamp 1586547711
transform 1 0 4448 0 -1 18352
box 0 -48 368 592
use sky130_fd_sc_hd__or4_4  _722_ ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 4816 0 -1 18352
box 0 -48 828 592
use sky130_fd_sc_hd__decap_8  FILL26220x87040
timestamp 1586547711
transform 1 0 5644 0 -1 18352
box 0 -48 736 592
use sky130_fd_sc_hd__or4_4  _733_
timestamp 1586547711
transform 1 0 6380 0 -1 18352
box 0 -48 828 592
use sky130_fd_sc_hd__decap_12  FILL34040x87040
timestamp 1586547711
transform 1 0 7208 0 -1 18352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL42780x87040
timestamp 1586547711
transform 1 0 8956 0 -1 18352
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1586547711
transform 1 0 8864 0 -1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL39560x87040
timestamp 1586547711
transform 1 0 8312 0 -1 18352
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL48300x87040
timestamp 1586547711
transform 1 0 10060 0 -1 18352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL53820x87040
timestamp 1586547711
transform 1 0 11164 0 -1 18352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL66240x87040
timestamp 1586547711
transform 1 0 13648 0 -1 18352
box 0 -48 736 592
use sky130_fd_sc_hd__decap_6  FILL59340x87040
timestamp 1586547711
transform 1 0 12268 0 -1 18352
box 0 -48 552 592
use sky130_fd_sc_hd__or3_4  _509_
timestamp 1586547711
transform 1 0 12820 0 -1 18352
box 0 -48 828 592
use sky130_fd_sc_hd__decap_12  FILL74060x87040
timestamp 1586547711
transform 1 0 15212 0 -1 18352
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL69920x87040
timestamp 1586547711
transform 1 0 14384 0 -1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1586547711
transform 1 0 14476 0 -1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _474_
timestamp 1586547711
transform 1 0 14568 0 -1 18352
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  FILL79580x87040
timestamp 1586547711
transform 1 0 16316 0 -1 18352
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_409
timestamp 1586547711
transform 1 0 17788 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL85100x87040
timestamp 1586547711
transform 1 0 17420 0 -1 18352
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILL87860x87040
timestamp 1586547711
transform 1 0 17972 0 -1 18352
box 0 -48 552 592
use sky130_fd_sc_hd__nor2_4  _590_
timestamp 1586547711
transform 1 0 16592 0 -1 18352
box 0 -48 828 592
use sky130_fd_sc_hd__decap_8  FILL94760x87040
timestamp 1586547711
transform 1 0 19352 0 -1 18352
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_935
timestamp 1586547711
transform 1 0 18984 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_937
timestamp 1586547711
transform 1 0 19168 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1586547711
transform 1 0 20088 0 -1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL98900x87040
timestamp 1586547711
transform 1 0 20180 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _545_
timestamp 1586547711
transform 1 0 18524 0 -1 18352
box 0 -48 460 592
use sky130_fd_sc_hd__dfstp_4  _854_
timestamp 1586547711
transform 1 0 20364 0 -1 18352
box 0 -48 2208 592
use sky130_fd_sc_hd__decap_12  FILL110860x87040
timestamp 1586547711
transform 1 0 22572 0 -1 18352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL118680x87040
timestamp 1586547711
transform 1 0 24136 0 -1 18352
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1633
timestamp 1586547711
transform 1 0 23768 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_397
timestamp 1586547711
transform 1 0 23952 0 -1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL116380x87040
timestamp 1586547711
transform 1 0 23676 0 -1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL126960x87040
timestamp 1586547711
transform 1 0 25792 0 -1 18352
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL126040x87040
timestamp 1586547711
transform 1 0 25608 0 -1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL130640x87040
timestamp 1586547711
transform 1 0 26528 0 -1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1586547711
transform 1 0 25700 0 -1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL124200x87040
timestamp 1586547711
transform 1 0 25240 0 -1 18352
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _631_
timestamp 1586547711
transform 1 0 26620 0 -1 18352
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL134320x87040
timestamp 1586547711
transform 1 0 27264 0 -1 18352
box 0 -48 736 592
use sky130_fd_sc_hd__dfrtp_4  _902_
timestamp 1586547711
transform 1 0 28000 0 -1 18352
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_12  FILL148580x87040
timestamp 1586547711
transform 1 0 30116 0 -1 18352
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL154100x87040
timestamp 1586547711
transform 1 0 31220 0 -1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1586547711
transform 1 0 31312 0 -1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1586547711
transform 1 0 31404 0 -1 18352
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL1380x92480
timestamp 1586547711
transform 1 0 676 0 -1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL8740x92480
timestamp 1586547711
transform 1 0 2148 0 -1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL1380x89760
timestamp 1586547711
transform 1 0 676 0 1 18352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL6900x89760
timestamp 1586547711
transform 1 0 1780 0 1 18352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1586547711
transform 1 0 400 0 -1 19440
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1586547711
transform 1 0 400 0 1 18352
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1283
timestamp 1586547711
transform 1 0 1964 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL6900x92480
timestamp 1586547711
transform 1 0 1780 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL17480x92480
timestamp 1586547711
transform 1 0 3896 0 -1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL16560x89760
timestamp 1586547711
transform 1 0 3712 0 1 18352
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_616
timestamp 1586547711
transform 1 0 3344 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1254
timestamp 1586547711
transform 1 0 3528 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL14260x89760
timestamp 1586547711
transform 1 0 3252 0 1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1586547711
transform 1 0 3252 0 -1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL12420x89760
timestamp 1586547711
transform 1 0 2884 0 1 18352
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL22080x89760
timestamp 1586547711
transform 1 0 4816 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _666_
timestamp 1586547711
transform 1 0 3344 0 -1 19440
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL25760x92480
timestamp 1586547711
transform 1 0 5552 0 -1 19440
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_615
timestamp 1586547711
transform 1 0 5000 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_620
timestamp 1586547711
transform 1 0 5184 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL27600x89760
timestamp 1586547711
transform 1 0 5920 0 1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL24840x89760
timestamp 1586547711
transform 1 0 5368 0 1 18352
box 0 -48 552 592
use sky130_fd_sc_hd__buf_4  _453_
timestamp 1586547711
transform 1 0 5000 0 -1 19440
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL31280x89760
timestamp 1586547711
transform 1 0 6656 0 1 18352
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_677
timestamp 1586547711
transform 1 0 7024 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_642
timestamp 1586547711
transform 1 0 6288 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1268
timestamp 1586547711
transform 1 0 6472 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1586547711
transform 1 0 6012 0 1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL32200x92480
timestamp 1586547711
transform 1 0 6840 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL28520x89760
timestamp 1586547711
transform 1 0 6104 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _670_
timestamp 1586547711
transform 1 0 6288 0 -1 19440
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL36800x89760
timestamp 1586547711
transform 1 0 7760 0 1 18352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL34040x92480
timestamp 1586547711
transform 1 0 7208 0 -1 19440
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL38180x92480
timestamp 1586547711
transform 1 0 8036 0 -1 19440
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_633
timestamp 1586547711
transform 1 0 7484 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_639
timestamp 1586547711
transform 1 0 7668 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_650
timestamp 1586547711
transform 1 0 7852 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILL42780x92480
timestamp 1586547711
transform 1 0 8956 0 -1 19440
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1260
timestamp 1586547711
transform 1 0 9232 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL41860x92480
timestamp 1586547711
transform 1 0 8772 0 -1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1586547711
transform 1 0 8864 0 -1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL42320x89760
timestamp 1586547711
transform 1 0 8864 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _442_
timestamp 1586547711
transform 1 0 9048 0 1 18352
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_634
timestamp 1586547711
transform 1 0 9508 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_641
timestamp 1586547711
transform 1 0 9692 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_574
timestamp 1586547711
transform 1 0 9600 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_577
timestamp 1586547711
transform 1 0 9784 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL45080x92480
timestamp 1586547711
transform 1 0 9416 0 -1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILL47840x89760
timestamp 1586547711
transform 1 0 9968 0 1 18352
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_313
timestamp 1586547711
transform 1 0 10244 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL47380x92480
timestamp 1586547711
transform 1 0 9876 0 -1 19440
box 0 -48 368 592
use sky130_fd_sc_hd__inv_4  _441_
timestamp 1586547711
transform 1 0 10244 0 -1 19440
box 0 -48 460 592
use sky130_fd_sc_hd__diode_2  ANTENNA_598
timestamp 1586547711
transform 1 0 10704 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_573
timestamp 1586547711
transform 1 0 10428 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL52440x92480
timestamp 1586547711
transform 1 0 10888 0 -1 19440
box 0 -48 552 592
use sky130_fd_sc_hd__decap_6  FILL51060x89760
timestamp 1586547711
transform 1 0 10612 0 1 18352
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_602
timestamp 1586547711
transform 1 0 11256 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_307
timestamp 1586547711
transform 1 0 11440 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL53820x89760
timestamp 1586547711
transform 1 0 11164 0 1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _448_
timestamp 1586547711
transform 1 0 11440 0 -1 19440
box 0 -48 460 592
use sky130_fd_sc_hd__diode_2  ANTENNA_580
timestamp 1586547711
transform 1 0 11900 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1365
timestamp 1586547711
transform 1 0 12084 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1586547711
transform 1 0 11624 0 1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _449_
timestamp 1586547711
transform 1 0 11716 0 1 18352
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_599
timestamp 1586547711
transform 1 0 12268 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_600
timestamp 1586547711
transform 1 0 12452 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_701
timestamp 1586547711
transform 1 0 12636 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_694
timestamp 1586547711
transform 1 0 12820 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL62100x92480
timestamp 1586547711
transform 1 0 12820 0 -1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL59340x92480
timestamp 1586547711
transform 1 0 12268 0 -1 19440
box 0 -48 552 592
use sky130_fd_sc_hd__or2_4  _473_
timestamp 1586547711
transform 1 0 12912 0 -1 19440
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL65780x92480
timestamp 1586547711
transform 1 0 13556 0 -1 19440
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_681
timestamp 1586547711
transform 1 0 13464 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_684
timestamp 1586547711
transform 1 0 13648 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _467_
timestamp 1586547711
transform 1 0 13004 0 1 18352
box 0 -48 460 592
use sky130_fd_sc_hd__decap_8  FILL68080x89760
timestamp 1586547711
transform 1 0 14016 0 1 18352
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_703
timestamp 1586547711
transform 1 0 13832 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL69460x92480
timestamp 1586547711
transform 1 0 14292 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILL70840x92480
timestamp 1586547711
transform 1 0 14568 0 -1 19440
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1514
timestamp 1586547711
transform 1 0 14844 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1596
timestamp 1586547711
transform 1 0 15028 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL71760x89760
timestamp 1586547711
transform 1 0 14752 0 1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1586547711
transform 1 0 14476 0 -1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _811_
timestamp 1586547711
transform 1 0 14844 0 -1 19440
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL74980x92480
timestamp 1586547711
transform 1 0 15396 0 -1 19440
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL74060x89760
timestamp 1586547711
transform 1 0 15212 0 1 18352
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILL82800x92480
timestamp 1586547711
transform 1 0 16960 0 -1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_706
timestamp 1586547711
transform 1 0 16132 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_977
timestamp 1586547711
transform 1 0 16316 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1145
timestamp 1586547711
transform 1 0 16500 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL81420x89760
timestamp 1586547711
transform 1 0 16684 0 1 18352
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL77740x89760
timestamp 1586547711
transform 1 0 15948 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _615_
timestamp 1586547711
transform 1 0 16132 0 -1 19440
box 0 -48 828 592
use sky130_fd_sc_hd__decap_12  FILL88320x92480
timestamp 1586547711
transform 1 0 18064 0 -1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1167
timestamp 1586547711
transform 1 0 17052 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_711
timestamp 1586547711
transform 1 0 17972 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1586547711
transform 1 0 17236 0 1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _628_
timestamp 1586547711
transform 1 0 17328 0 1 18352
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL89700x89760
timestamp 1586547711
transform 1 0 18340 0 1 18352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL95220x89760
timestamp 1586547711
transform 1 0 19444 0 1 18352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL93840x92480
timestamp 1586547711
transform 1 0 19168 0 -1 19440
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1146
timestamp 1586547711
transform 1 0 20180 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_978
timestamp 1586547711
transform 1 0 18156 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1586547711
transform 1 0 20088 0 -1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL97520x92480
timestamp 1586547711
transform 1 0 19904 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL100740x89760
timestamp 1586547711
transform 1 0 20548 0 1 18352
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1079
timestamp 1586547711
transform 1 0 20916 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1104
timestamp 1586547711
transform 1 0 21100 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1105
timestamp 1586547711
transform 1 0 21284 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL99820x92480
timestamp 1586547711
transform 1 0 20364 0 -1 19440
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILL106260x89760
timestamp 1586547711
transform 1 0 21652 0 1 18352
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL110400x92480
timestamp 1586547711
transform 1 0 22480 0 -1 19440
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_325
timestamp 1586547711
transform 1 0 21928 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_626
timestamp 1586547711
transform 1 0 22112 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL107180x92480
timestamp 1586547711
transform 1 0 21836 0 -1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL105340x92480
timestamp 1586547711
transform 1 0 21468 0 -1 19440
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILL109480x89760
timestamp 1586547711
transform 1 0 22296 0 1 18352
box 0 -48 552 592
use sky130_fd_sc_hd__buf_4  _455_
timestamp 1586547711
transform 1 0 21928 0 -1 19440
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1143
timestamp 1586547711
transform 1 0 23032 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1142
timestamp 1586547711
transform 1 0 23216 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_138
timestamp 1586547711
transform 1 0 23400 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1586547711
transform 1 0 23584 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL112700x89760
timestamp 1586547711
transform 1 0 22940 0 1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1586547711
transform 1 0 22848 0 1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _614_
timestamp 1586547711
transform 1 0 23216 0 -1 19440
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL117760x92480
timestamp 1586547711
transform 1 0 23952 0 -1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_399
timestamp 1586547711
transform 1 0 23768 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL116380x92480
timestamp 1586547711
transform 1 0 23676 0 -1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__dfstp_4  _863_
timestamp 1586547711
transform 1 0 23768 0 1 18352
box 0 -48 2208 592
use sky130_fd_sc_hd__decap_12  FILL126960x92480
timestamp 1586547711
transform 1 0 25792 0 -1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1252
timestamp 1586547711
transform 1 0 26620 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1251
timestamp 1586547711
transform 1 0 26804 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL126040x92480
timestamp 1586547711
transform 1 0 25608 0 -1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL130640x89760
timestamp 1586547711
transform 1 0 26528 0 1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1586547711
transform 1 0 25700 0 -1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL123280x92480
timestamp 1586547711
transform 1 0 25056 0 -1 19440
box 0 -48 552 592
use sky130_fd_sc_hd__decap_6  FILL127880x89760
timestamp 1586547711
transform 1 0 25976 0 1 18352
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILL132480x92480
timestamp 1586547711
transform 1 0 26896 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1243
timestamp 1586547711
transform 1 0 26988 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_970
timestamp 1586547711
transform 1 0 27632 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1169
timestamp 1586547711
transform 1 0 27816 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1175
timestamp 1586547711
transform 1 0 28000 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _630_
timestamp 1586547711
transform 1 0 27172 0 1 18352
box 0 -48 460 592
use sky130_fd_sc_hd__o21a_4  _664_
timestamp 1586547711
transform 1 0 27080 0 -1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1242
timestamp 1586547711
transform 1 0 28552 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1178
timestamp 1586547711
transform 1 0 28276 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL138920x89760
timestamp 1586547711
transform 1 0 28184 0 1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1586547711
transform 1 0 28460 0 1 18352
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL138920x92480
timestamp 1586547711
transform 1 0 28184 0 -1 19440
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL141680x92480
timestamp 1586547711
transform 1 0 28736 0 -1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _644_
timestamp 1586547711
transform 1 0 28920 0 -1 19440
box 0 -48 644 592
use sky130_fd_sc_hd__and2_4  _659_
timestamp 1586547711
transform 1 0 28552 0 1 18352
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL145820x92480
timestamp 1586547711
transform 1 0 29564 0 -1 19440
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_191
timestamp 1586547711
transform 1 0 29196 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_195
timestamp 1586547711
transform 1 0 29380 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1170
timestamp 1586547711
transform 1 0 29564 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1216
timestamp 1586547711
transform 1 0 29748 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL150880x92480
timestamp 1586547711
transform 1 0 30576 0 -1 19440
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL150420x89760
timestamp 1586547711
transform 1 0 30484 0 1 18352
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_173
timestamp 1586547711
transform 1 0 30300 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL147660x89760
timestamp 1586547711
transform 1 0 29932 0 1 18352
box 0 -48 368 592
use sky130_fd_sc_hd__conb_1  _841_
timestamp 1586547711
transform 1 0 30300 0 -1 19440
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1586547711
transform 1 0 31312 0 -1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL154100x89760
timestamp 1586547711
transform 1 0 31220 0 1 18352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1586547711
transform 1 0 31404 0 -1 19440
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1586547711
transform 1 0 31404 0 1 18352
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1586547711
transform 1 0 400 0 1 19440
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL1380x95200
timestamp 1586547711
transform 1 0 676 0 1 19440
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_189
timestamp 1586547711
transform 1 0 1228 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1297
timestamp 1586547711
transform 1 0 1412 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_637
timestamp 1586547711
transform 1 0 1596 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_430
timestamp 1586547711
transform 1 0 1780 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__conb_1  _843_
timestamp 1586547711
transform 1 0 952 0 1 19440
box 0 -48 276 592
use sky130_fd_sc_hd__o22ai_4  _679_
timestamp 1586547711
transform 1 0 1964 0 1 19440
box 0 -48 1472 592
use sky130_fd_sc_hd__decap_12  FILL17020x95200
timestamp 1586547711
transform 1 0 3804 0 1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_205
timestamp 1586547711
transform 1 0 3436 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_632
timestamp 1586547711
transform 1 0 3620 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL22540x95200
timestamp 1586547711
transform 1 0 4908 0 1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1264
timestamp 1586547711
transform 1 0 6472 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_596
timestamp 1586547711
transform 1 0 6656 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_575
timestamp 1586547711
transform 1 0 6840 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_564
timestamp 1586547711
transform 1 0 7024 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1586547711
transform 1 0 6012 0 1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL28520x95200
timestamp 1586547711
transform 1 0 6104 0 1 19440
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_532
timestamp 1586547711
transform 1 0 7300 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_675
timestamp 1586547711
transform 1 0 8772 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_579
timestamp 1586547711
transform 1 0 8956 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_572
timestamp 1586547711
transform 1 0 9140 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL34040x95200
timestamp 1586547711
transform 1 0 7208 0 1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _459_
timestamp 1586547711
transform 1 0 7484 0 1 19440
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA_534
timestamp 1586547711
transform 1 0 9324 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_478
timestamp 1586547711
transform 1 0 10796 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_543
timestamp 1586547711
transform 1 0 10980 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_569
timestamp 1586547711
transform 1 0 11164 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_578
timestamp 1586547711
transform 1 0 11348 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _466_
timestamp 1586547711
transform 1 0 9508 0 1 19440
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA_535
timestamp 1586547711
transform 1 0 12544 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL55660x95200
timestamp 1586547711
transform 1 0 11532 0 1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1586547711
transform 1 0 11624 0 1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL61640x95200
timestamp 1586547711
transform 1 0 12728 0 1 19440
box 0 -48 552 592
use sky130_fd_sc_hd__inv_4  _508_
timestamp 1586547711
transform 1 0 13280 0 1 19440
box 0 -48 460 592
use sky130_fd_sc_hd__and3_4  _709_
timestamp 1586547711
transform 1 0 11716 0 1 19440
box 0 -48 828 592
use sky130_fd_sc_hd__decap_12  FILL72680x95200
timestamp 1586547711
transform 1 0 14936 0 1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_702
timestamp 1586547711
transform 1 0 13740 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_836
timestamp 1586547711
transform 1 0 13924 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1690
timestamp 1586547711
transform 1 0 14568 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1697
timestamp 1586547711
transform 1 0 14752 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL70380x95200
timestamp 1586547711
transform 1 0 14476 0 1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL68540x95200
timestamp 1586547711
transform 1 0 14108 0 1 19440
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILL78200x95200
timestamp 1586547711
transform 1 0 16040 0 1 19440
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_44
timestamp 1586547711
transform 1 0 16500 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL80040x95200
timestamp 1586547711
transform 1 0 16408 0 1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_755
timestamp 1586547711
transform 1 0 16684 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL82340x95200
timestamp 1586547711
transform 1 0 16868 0 1 19440
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1586547711
transform 1 0 17236 0 1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL84640x95200
timestamp 1586547711
transform 1 0 17328 0 1 19440
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILL86480x95200
timestamp 1586547711
transform 1 0 17696 0 1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1530
timestamp 1586547711
transform 1 0 17788 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1598
timestamp 1586547711
transform 1 0 17972 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL88780x95200
timestamp 1586547711
transform 1 0 18156 0 1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1147
timestamp 1586547711
transform 1 0 19628 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_942
timestamp 1586547711
transform 1 0 19812 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_50
timestamp 1586547711
transform 1 0 19996 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL94300x95200
timestamp 1586547711
transform 1 0 19260 0 1 19440
box 0 -48 368 592
use sky130_fd_sc_hd__a211o_4  _616_
timestamp 1586547711
transform 1 0 20180 0 1 19440
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_8  FILL107180x95200
timestamp 1586547711
transform 1 0 21836 0 1 19440
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_53
timestamp 1586547711
transform 1 0 21468 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_940
timestamp 1586547711
transform 1 0 21652 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL117760x95200
timestamp 1586547711
transform 1 0 23952 0 1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1078
timestamp 1586547711
transform 1 0 22664 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1072
timestamp 1586547711
transform 1 0 23584 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1076
timestamp 1586547711
transform 1 0 23768 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL110860x95200
timestamp 1586547711
transform 1 0 22572 0 1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1586547711
transform 1 0 22848 0 1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _591_
timestamp 1586547711
transform 1 0 22940 0 1 19440
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL123280x95200
timestamp 1586547711
transform 1 0 25056 0 1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL132480x95200
timestamp 1586547711
transform 1 0 26896 0 1 19440
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL128800x95200
timestamp 1586547711
transform 1 0 26160 0 1 19440
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1357
timestamp 1586547711
transform 1 0 27172 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_46
timestamp 1586547711
transform 1 0 27356 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_426
timestamp 1586547711
transform 1 0 27540 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1068
timestamp 1586547711
transform 1 0 27724 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1241
timestamp 1586547711
transform 1 0 27908 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1253
timestamp 1586547711
transform 1 0 28092 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL140760x95200
timestamp 1586547711
transform 1 0 28552 0 1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1586547711
transform 1 0 28460 0 1 19440
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL139380x95200
timestamp 1586547711
transform 1 0 28276 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _422_
timestamp 1586547711
transform 1 0 28644 0 1 19440
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL145820x95200
timestamp 1586547711
transform 1 0 29564 0 1 19440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL151340x95200
timestamp 1586547711
transform 1 0 30668 0 1 19440
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1614
timestamp 1586547711
transform 1 0 29196 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1619
timestamp 1586547711
transform 1 0 29380 0 1 19440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1586547711
transform 1 0 31404 0 1 19440
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1586547711
transform 1 0 400 0 -1 20528
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_431
timestamp 1586547711
transform 1 0 676 0 -1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1682
timestamp 1586547711
transform 1 0 860 0 -1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1540
timestamp 1586547711
transform 1 0 1136 0 -1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1604
timestamp 1586547711
transform 1 0 1320 0 -1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL3220x97920
timestamp 1586547711
transform 1 0 1044 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL5520x97920
timestamp 1586547711
transform 1 0 1504 0 -1 20528
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL8740x97920
timestamp 1586547711
transform 1 0 2148 0 -1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1256
timestamp 1586547711
transform 1 0 1964 0 -1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL7360x97920
timestamp 1586547711
transform 1 0 1872 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL17020x97920
timestamp 1586547711
transform 1 0 3804 0 -1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1586547711
transform 1 0 3252 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _456_
timestamp 1586547711
transform 1 0 3344 0 -1 20528
box 0 -48 460 592
use sky130_fd_sc_hd__decap_8  FILL22540x97920
timestamp 1586547711
transform 1 0 4908 0 -1 20528
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1276
timestamp 1586547711
transform 1 0 5736 0 -1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1288
timestamp 1586547711
transform 1 0 5920 0 -1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_646
timestamp 1586547711
transform 1 0 6656 0 -1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL26220x97920
timestamp 1586547711
transform 1 0 5644 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL28520x97920
timestamp 1586547711
transform 1 0 6104 0 -1 20528
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILL32200x97920
timestamp 1586547711
transform 1 0 6840 0 -1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _669_
timestamp 1586547711
transform 1 0 7024 0 -1 20528
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  FILL42780x97920
timestamp 1586547711
transform 1 0 8956 0 -1 20528
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_645
timestamp 1586547711
transform 1 0 7852 0 -1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1262
timestamp 1586547711
transform 1 0 8680 0 -1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL40940x97920
timestamp 1586547711
transform 1 0 8588 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1586547711
transform 1 0 8864 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL38180x97920
timestamp 1586547711
transform 1 0 8036 0 -1 20528
box 0 -48 552 592
use sky130_fd_sc_hd__or2_4  _667_
timestamp 1586547711
transform 1 0 9232 0 -1 20528
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_680
timestamp 1586547711
transform 1 0 9876 0 -1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL48300x97920
timestamp 1586547711
transform 1 0 10060 0 -1 20528
box 0 -48 552 592
use sky130_fd_sc_hd__o22ai_4  _447_
timestamp 1586547711
transform 1 0 10612 0 -1 20528
box 0 -48 1472 592
use sky130_fd_sc_hd__decap_12  FILL59340x97920
timestamp 1586547711
transform 1 0 12268 0 -1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL64860x97920
timestamp 1586547711
transform 1 0 13372 0 -1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_601
timestamp 1586547711
transform 1 0 12084 0 -1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL73600x97920
timestamp 1586547711
transform 1 0 15120 0 -1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1586547711
transform 1 0 14476 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_4  _CTS_buf_1_48
timestamp 1586547711
transform 1 0 14568 0 -1 20528
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILL79120x97920
timestamp 1586547711
transform 1 0 16224 0 -1 20528
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_625
timestamp 1586547711
transform 1 0 17052 0 -1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_453
timestamp 1586547711
transform 1 0 17328 0 -1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1531
timestamp 1586547711
transform 1 0 17512 0 -1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL84180x97920
timestamp 1586547711
transform 1 0 17236 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL86480x97920
timestamp 1586547711
transform 1 0 17696 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _483_
timestamp 1586547711
transform 1 0 16500 0 -1 20528
box 0 -48 552 592
use sky130_fd_sc_hd__buf_4  _813_
timestamp 1586547711
transform 1 0 17788 0 -1 20528
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL89700x97920
timestamp 1586547711
transform 1 0 18340 0 -1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1080
timestamp 1586547711
transform 1 0 20180 0 -1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL97980x97920
timestamp 1586547711
transform 1 0 19996 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1586547711
transform 1 0 20088 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL95220x97920
timestamp 1586547711
transform 1 0 19444 0 -1 20528
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL109020x97920
timestamp 1586547711
transform 1 0 22204 0 -1 20528
box 0 -48 736 592
use sky130_fd_sc_hd__decap_6  FILL99820x97920
timestamp 1586547711
transform 1 0 20364 0 -1 20528
box 0 -48 552 592
use sky130_fd_sc_hd__a211o_4  _602_
timestamp 1586547711
transform 1 0 20916 0 -1 20528
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL114540x97920
timestamp 1586547711
transform 1 0 23308 0 -1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL120060x97920
timestamp 1586547711
transform 1 0 24412 0 -1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1144
timestamp 1586547711
transform 1 0 22940 0 -1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1148
timestamp 1586547711
transform 1 0 23124 0 -1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL126960x97920
timestamp 1586547711
transform 1 0 25792 0 -1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1586547711
transform 1 0 25700 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL132480x97920
timestamp 1586547711
transform 1 0 26896 0 -1 20528
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL125580x97920
timestamp 1586547711
transform 1 0 25516 0 -1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL143060x97920
timestamp 1586547711
transform 1 0 29012 0 -1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL134320x97920
timestamp 1586547711
transform 1 0 27264 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__o32a_4  _665_
timestamp 1586547711
transform 1 0 27356 0 -1 20528
box 0 -48 1656 592
use sky130_fd_sc_hd__decap_12  FILL148580x97920
timestamp 1586547711
transform 1 0 30116 0 -1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL154100x97920
timestamp 1586547711
transform 1 0 31220 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1586547711
transform 1 0 31312 0 -1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1586547711
transform 1 0 31404 0 -1 20528
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1586547711
transform 1 0 400 0 1 20528
box 0 -48 276 592
use sky130_fd_sc_hd__dfrtp_4  _919_
timestamp 1586547711
transform 1 0 676 0 1 20528
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1296
timestamp 1586547711
transform 1 0 3344 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1294
timestamp 1586547711
transform 1 0 3528 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_538
timestamp 1586547711
transform 1 0 3712 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_679
timestamp 1586547711
transform 1 0 3896 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1289
timestamp 1586547711
transform 1 0 4080 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1290
timestamp 1586547711
transform 1 0 4264 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL11960x100640
timestamp 1586547711
transform 1 0 2792 0 1 20528
box 0 -48 552 592
use sky130_fd_sc_hd__or2_4  _676_
timestamp 1586547711
transform 1 0 4448 0 1 20528
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_636
timestamp 1586547711
transform 1 0 5092 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1267
timestamp 1586547711
transform 1 0 5276 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1266
timestamp 1586547711
transform 1 0 5552 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_635
timestamp 1586547711
transform 1 0 5736 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL25300x100640
timestamp 1586547711
transform 1 0 5460 0 1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL27600x100640
timestamp 1586547711
transform 1 0 5920 0 1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_658
timestamp 1586547711
transform 1 0 6104 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_640
timestamp 1586547711
transform 1 0 6288 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_533
timestamp 1586547711
transform 1 0 6472 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1586547711
transform 1 0 6012 0 1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _462_
timestamp 1586547711
transform 1 0 6656 0 1 20528
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA_676
timestamp 1586547711
transform 1 0 8312 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_595
timestamp 1586547711
transform 1 0 8496 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL37720x100640
timestamp 1586547711
transform 1 0 7944 0 1 20528
box 0 -48 368 592
use sky130_fd_sc_hd__o21ai_4  _668_ ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 8680 0 1 20528
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA_621
timestamp 1586547711
transform 1 0 10336 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_314
timestamp 1586547711
transform 1 0 10520 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_446
timestamp 1586547711
transform 1 0 10704 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_571
timestamp 1586547711
transform 1 0 10888 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_586
timestamp 1586547711
transform 1 0 11072 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_594
timestamp 1586547711
transform 1 0 11256 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_597
timestamp 1586547711
transform 1 0 11440 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL49220x100640
timestamp 1586547711
transform 1 0 10244 0 1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL47380x100640
timestamp 1586547711
transform 1 0 9876 0 1 20528
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL63940x100640
timestamp 1586547711
transform 1 0 13188 0 1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_584
timestamp 1586547711
transform 1 0 12360 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_593
timestamp 1586547711
transform 1 0 12544 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_563
timestamp 1586547711
transform 1 0 12820 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_567
timestamp 1586547711
transform 1 0 13004 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL61640x100640
timestamp 1586547711
transform 1 0 12728 0 1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1586547711
transform 1 0 11624 0 1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _446_
timestamp 1586547711
transform 1 0 11716 0 1 20528
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL69460x100640
timestamp 1586547711
transform 1 0 14292 0 1 20528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL74980x100640
timestamp 1586547711
transform 1 0 15396 0 1 20528
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1379
timestamp 1586547711
transform 1 0 16132 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_971
timestamp 1586547711
transform 1 0 16316 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_758
timestamp 1586547711
transform 1 0 16500 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_452
timestamp 1586547711
transform 1 0 16684 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_324
timestamp 1586547711
transform 1 0 16868 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_322
timestamp 1586547711
transform 1 0 17052 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1586547711
transform 1 0 17236 0 1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _914_
timestamp 1586547711
transform 1 0 17328 0 1 20528
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1575
timestamp 1586547711
transform 1 0 19996 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL95220x100640
timestamp 1586547711
transform 1 0 19444 0 1 20528
box 0 -48 552 592
use sky130_fd_sc_hd__or2_4  _786_
timestamp 1586547711
transform 1 0 20180 0 1 20528
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_323
timestamp 1586547711
transform 1 0 20824 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_631
timestamp 1586547711
transform 1 0 21008 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1354
timestamp 1586547711
transform 1 0 21376 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL103960x100640
timestamp 1586547711
transform 1 0 21192 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1064
timestamp 1586547711
transform 1 0 21560 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_256
timestamp 1586547711
transform 1 0 21744 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_412
timestamp 1586547711
transform 1 0 21928 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_967
timestamp 1586547711
transform 1 0 22112 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1058
timestamp 1586547711
transform 1 0 22296 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_968
timestamp 1586547711
transform 1 0 22480 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_260
timestamp 1586547711
transform 1 0 22664 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1074
timestamp 1586547711
transform 1 0 24228 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1206
timestamp 1586547711
transform 1 0 24412 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1586547711
transform 1 0 22848 0 1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL120980x100640
timestamp 1586547711
transform 1 0 24596 0 1 20528
box 0 -48 368 592
use sky130_fd_sc_hd__o22a_4  _617_
timestamp 1586547711
transform 1 0 22940 0 1 20528
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_8  FILL127420x100640
timestamp 1586547711
transform 1 0 25884 0 1 20528
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_961
timestamp 1586547711
transform 1 0 25516 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_966
timestamp 1586547711
transform 1 0 25700 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1224
timestamp 1586547711
transform 1 0 26804 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL131100x100640
timestamp 1586547711
transform 1 0 26620 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _554_
timestamp 1586547711
transform 1 0 24964 0 1 20528
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_269
timestamp 1586547711
transform 1 0 26988 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_964
timestamp 1586547711
transform 1 0 27172 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1208
timestamp 1586547711
transform 1 0 27356 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1217
timestamp 1586547711
transform 1 0 27540 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1223
timestamp 1586547711
transform 1 0 27724 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1479
timestamp 1586547711
transform 1 0 27908 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_427
timestamp 1586547711
transform 1 0 28092 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_47
timestamp 1586547711
transform 1 0 28276 0 1 20528
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1586547711
transform 1 0 28460 0 1 20528
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _901_
timestamp 1586547711
transform 1 0 28552 0 1 20528
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_8  FILL151340x100640
timestamp 1586547711
transform 1 0 30668 0 1 20528
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1586547711
transform 1 0 31404 0 1 20528
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL6440x103360
timestamp 1586547711
transform 1 0 1688 0 -1 21616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1586547711
transform 1 0 400 0 -1 21616
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_207
timestamp 1586547711
transform 1 0 676 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1541
timestamp 1586547711
transform 1 0 860 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL3220x103360
timestamp 1586547711
transform 1 0 1044 0 -1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _819_
timestamp 1586547711
transform 1 0 1136 0 -1 21616
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1299
timestamp 1586547711
transform 1 0 3344 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1301
timestamp 1586547711
transform 1 0 3528 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL13800x103360
timestamp 1586547711
transform 1 0 3160 0 -1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1586547711
transform 1 0 3252 0 -1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL11960x103360
timestamp 1586547711
transform 1 0 2792 0 -1 21616
box 0 -48 368 592
use sky130_fd_sc_hd__o22a_4  _678_
timestamp 1586547711
transform 1 0 3712 0 -1 21616
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_8  FILL23000x103360
timestamp 1586547711
transform 1 0 5000 0 -1 21616
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_662
timestamp 1586547711
transform 1 0 6840 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL33120x103360
timestamp 1586547711
transform 1 0 7024 0 -1 21616
box 0 -48 368 592
use sky130_fd_sc_hd__o21a_4  _675_
timestamp 1586547711
transform 1 0 5736 0 -1 21616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL35880x103360
timestamp 1586547711
transform 1 0 7576 0 -1 21616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL42780x103360
timestamp 1586547711
transform 1 0 8956 0 -1 21616
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_638
timestamp 1586547711
transform 1 0 7392 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1261
timestamp 1586547711
transform 1 0 8680 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1586547711
transform 1 0 8864 0 -1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL50140x103360
timestamp 1586547711
transform 1 0 10428 0 -1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL48300x103360
timestamp 1586547711
transform 1 0 10060 0 -1 21616
box 0 -48 368 592
use sky130_fd_sc_hd__a32o_4  _454_
timestamp 1586547711
transform 1 0 10520 0 -1 21616
box 0 -48 1564 592
use sky130_fd_sc_hd__decap_8  FILL58420x103360
timestamp 1586547711
transform 1 0 12084 0 -1 21616
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL65780x103360
timestamp 1586547711
transform 1 0 13556 0 -1 21616
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1691
timestamp 1586547711
transform 1 0 13372 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _440_
timestamp 1586547711
transform 1 0 12820 0 -1 21616
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL72220x103360
timestamp 1586547711
transform 1 0 14844 0 -1 21616
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1573
timestamp 1586547711
transform 1 0 14660 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL70840x103360
timestamp 1586547711
transform 1 0 14568 0 -1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1586547711
transform 1 0 14476 0 -1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL69460x103360
timestamp 1586547711
transform 1 0 14292 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL77740x103360
timestamp 1586547711
transform 1 0 15948 0 -1 21616
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1677
timestamp 1586547711
transform 1 0 16868 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL81420x103360
timestamp 1586547711
transform 1 0 16684 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__a32o_4  _717_
timestamp 1586547711
transform 1 0 17052 0 -1 21616
box 0 -48 1564 592
use sky130_fd_sc_hd__decap_12  FILL91080x103360
timestamp 1586547711
transform 1 0 18616 0 -1 21616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL98900x103360
timestamp 1586547711
transform 1 0 20180 0 -1 21616
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1586547711
transform 1 0 20088 0 -1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL96600x103360
timestamp 1586547711
transform 1 0 19720 0 -1 21616
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILL106260x103360
timestamp 1586547711
transform 1 0 21652 0 -1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL104420x103360
timestamp 1586547711
transform 1 0 21284 0 -1 21616
box 0 -48 368 592
use sky130_fd_sc_hd__a32o_4  _587_
timestamp 1586547711
transform 1 0 21744 0 -1 21616
box 0 -48 1564 592
use sky130_fd_sc_hd__decap_8  FILL115460x103360
timestamp 1586547711
transform 1 0 23492 0 -1 21616
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1149
timestamp 1586547711
transform 1 0 23308 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _640_
timestamp 1586547711
transform 1 0 24228 0 -1 21616
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILL131560x103360
timestamp 1586547711
transform 1 0 26712 0 -1 21616
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL121900x103360
timestamp 1586547711
transform 1 0 24780 0 -1 21616
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL127880x103360
timestamp 1586547711
transform 1 0 25976 0 -1 21616
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1207
timestamp 1586547711
transform 1 0 25792 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1586547711
transform 1 0 25700 0 -1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL125580x103360
timestamp 1586547711
transform 1 0 25516 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1620
timestamp 1586547711
transform 1 0 29012 0 -1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__a32oi_4  _648_
timestamp 1586547711
transform 1 0 26988 0 -1 21616
box 0 -48 2024 592
use sky130_fd_sc_hd__decap_12  FILL143980x103360
timestamp 1586547711
transform 1 0 29196 0 -1 21616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL153180x103360
timestamp 1586547711
transform 1 0 31036 0 -1 21616
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL149500x103360
timestamp 1586547711
transform 1 0 30300 0 -1 21616
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1586547711
transform 1 0 31312 0 -1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1586547711
transform 1 0 31404 0 -1 21616
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL5520x108800
timestamp 1586547711
transform 1 0 1504 0 -1 22704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL1380x106080
timestamp 1586547711
transform 1 0 676 0 1 21616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1586547711
transform 1 0 400 0 -1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1586547711
transform 1 0 400 0 1 21616
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_433
timestamp 1586547711
transform 1 0 676 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1683
timestamp 1586547711
transform 1 0 860 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1542
timestamp 1586547711
transform 1 0 1136 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1605
timestamp 1586547711
transform 1 0 1320 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL3220x108800
timestamp 1586547711
transform 1 0 1044 0 -1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1293
timestamp 1586547711
transform 1 0 2240 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1291
timestamp 1586547711
transform 1 0 2424 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL8740x106080
timestamp 1586547711
transform 1 0 2148 0 1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL6900x106080
timestamp 1586547711
transform 1 0 1780 0 1 21616
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILL11040x108800
timestamp 1586547711
transform 1 0 2608 0 -1 22704
box 0 -48 552 592
use sky130_fd_sc_hd__inv_4  _677_
timestamp 1586547711
transform 1 0 2608 0 1 21616
box 0 -48 460 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1277
timestamp 1586547711
transform 1 0 3160 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_206
timestamp 1586547711
transform 1 0 3344 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_546
timestamp 1586547711
transform 1 0 3528 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL13800x108800
timestamp 1586547711
transform 1 0 3160 0 -1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL13340x106080
timestamp 1586547711
transform 1 0 3068 0 1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL16560x106080
timestamp 1586547711
transform 1 0 3712 0 1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1586547711
transform 1 0 3252 0 -1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_647
timestamp 1586547711
transform 1 0 4448 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1292
timestamp 1586547711
transform 1 0 4632 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1300
timestamp 1586547711
transform 1 0 4816 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _681_
timestamp 1586547711
transform 1 0 3804 0 1 21616
box 0 -48 644 592
use sky130_fd_sc_hd__a32oi_4  _682_
timestamp 1586547711
transform 1 0 3344 0 -1 22704
box 0 -48 2024 592
use sky130_fd_sc_hd__decap_8  FILL24840x108800
timestamp 1586547711
transform 1 0 5368 0 -1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1304
timestamp 1586547711
transform 1 0 5000 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1275
timestamp 1586547711
transform 1 0 5276 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1263
timestamp 1586547711
transform 1 0 5460 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_757
timestamp 1586547711
transform 1 0 5644 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_545
timestamp 1586547711
transform 1 0 5828 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL23920x106080
timestamp 1586547711
transform 1 0 5184 0 1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1255
timestamp 1586547711
transform 1 0 6104 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1265
timestamp 1586547711
transform 1 0 6288 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1280
timestamp 1586547711
transform 1 0 6472 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_536
timestamp 1586547711
transform 1 0 6840 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1586547711
transform 1 0 6012 0 1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL33120x108800
timestamp 1586547711
transform 1 0 7024 0 -1 22704
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL31280x108800
timestamp 1586547711
transform 1 0 6656 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__a32oi_4  _672_
timestamp 1586547711
transform 1 0 6104 0 1 21616
box 0 -48 2024 592
use sky130_fd_sc_hd__decap_12  FILL39560x106080
timestamp 1586547711
transform 1 0 8312 0 1 21616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL37720x108800
timestamp 1586547711
transform 1 0 7944 0 -1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL42780x108800
timestamp 1586547711
transform 1 0 8956 0 -1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_318
timestamp 1586547711
transform 1 0 8128 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1586547711
transform 1 0 8864 0 -1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL41400x108800
timestamp 1586547711
transform 1 0 8680 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _457_
timestamp 1586547711
transform 1 0 7392 0 -1 22704
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILL46460x108800
timestamp 1586547711
transform 1 0 9692 0 -1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL51520x106080
timestamp 1586547711
transform 1 0 10704 0 1 21616
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_311
timestamp 1586547711
transform 1 0 9968 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_447
timestamp 1586547711
transform 1 0 10152 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1572
timestamp 1586547711
transform 1 0 10336 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1689
timestamp 1586547711
transform 1 0 10520 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL45080x106080
timestamp 1586547711
transform 1 0 9416 0 1 21616
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILL55200x106080
timestamp 1586547711
transform 1 0 11440 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__dfstp_4  _926_
timestamp 1586547711
transform 1 0 9968 0 -1 22704
box 0 -48 2208 592
use sky130_fd_sc_hd__decap_8  FILL56580x106080
timestamp 1586547711
transform 1 0 11716 0 1 21616
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_698
timestamp 1586547711
transform 1 0 12176 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1586547711
transform 1 0 11624 0 1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL59800x108800
timestamp 1586547711
transform 1 0 12360 0 -1 22704
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILL60260x106080
timestamp 1586547711
transform 1 0 12452 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL65780x108800
timestamp 1586547711
transform 1 0 13556 0 -1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1574
timestamp 1586547711
transform 1 0 13372 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_583
timestamp 1586547711
transform 1 0 12636 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_568
timestamp 1586547711
transform 1 0 12820 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_479
timestamp 1586547711
transform 1 0 13004 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_316
timestamp 1586547711
transform 1 0 13188 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _443_
timestamp 1586547711
transform 1 0 12912 0 -1 22704
box 0 -48 460 592
use sky130_fd_sc_hd__dfrtp_4  _927_
timestamp 1586547711
transform 1 0 13372 0 1 21616
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_12  FILL74060x108800
timestamp 1586547711
transform 1 0 15212 0 -1 22704
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_512
timestamp 1586547711
transform 1 0 15488 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL70840x108800
timestamp 1586547711
transform 1 0 14568 0 -1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1586547711
transform 1 0 14476 0 -1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL76360x106080
timestamp 1586547711
transform 1 0 15672 0 1 21616
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILL69460x108800
timestamp 1586547711
transform 1 0 14292 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _828_
timestamp 1586547711
transform 1 0 14660 0 -1 22704
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_43
timestamp 1586547711
transform 1 0 16316 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_697
timestamp 1586547711
transform 1 0 16500 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_587
timestamp 1586547711
transform 1 0 16868 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL79120x106080
timestamp 1586547711
transform 1 0 16224 0 1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL81880x108800
timestamp 1586547711
transform 1 0 16776 0 -1 22704
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILL81420x106080
timestamp 1586547711
transform 1 0 16684 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _471_
timestamp 1586547711
transform 1 0 16316 0 -1 22704
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL85560x108800
timestamp 1586547711
transform 1 0 17512 0 -1 22704
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1576
timestamp 1586547711
transform 1 0 17328 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_476
timestamp 1586547711
transform 1 0 17052 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1586547711
transform 1 0 17236 0 1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__and3_4  _787_
timestamp 1586547711
transform 1 0 17328 0 1 21616
box 0 -48 828 592
use sky130_fd_sc_hd__decap_8  FILL93840x108800
timestamp 1586547711
transform 1 0 19168 0 -1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_329
timestamp 1586547711
transform 1 0 18616 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_499
timestamp 1586547711
transform 1 0 18800 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1449
timestamp 1586547711
transform 1 0 18984 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_315
timestamp 1586547711
transform 1 0 18156 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1378
timestamp 1586547711
transform 1 0 18708 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL89700x106080
timestamp 1586547711
transform 1 0 18340 0 1 21616
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _716_
timestamp 1586547711
transform 1 0 18892 0 1 21616
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL98900x108800
timestamp 1586547711
transform 1 0 20180 0 -1 22704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL97520x106080
timestamp 1586547711
transform 1 0 19904 0 1 21616
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_605
timestamp 1586547711
transform 1 0 19536 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1211
timestamp 1586547711
transform 1 0 19720 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1586547711
transform 1 0 20088 0 -1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL97520x108800
timestamp 1586547711
transform 1 0 19904 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL104420x108800
timestamp 1586547711
transform 1 0 21284 0 -1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1106
timestamp 1586547711
transform 1 0 21652 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1070
timestamp 1586547711
transform 1 0 21836 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_259
timestamp 1586547711
transform 1 0 22020 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_414
timestamp 1586547711
transform 1 0 22204 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_516
timestamp 1586547711
transform 1 0 22388 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL105800x106080
timestamp 1586547711
transform 1 0 21560 0 1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL103040x106080
timestamp 1586547711
transform 1 0 21008 0 1 21616
box 0 -48 552 592
use sky130_fd_sc_hd__a32o_4  _603_
timestamp 1586547711
transform 1 0 22020 0 -1 22704
box 0 -48 1564 592
use sky130_fd_sc_hd__decap_12  FILL118680x108800
timestamp 1586547711
transform 1 0 24136 0 -1 22704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL112700x106080
timestamp 1586547711
transform 1 0 22940 0 1 21616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL118220x106080
timestamp 1586547711
transform 1 0 24044 0 1 21616
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1162
timestamp 1586547711
transform 1 0 23952 0 -1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1065
timestamp 1586547711
transform 1 0 22572 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL111780x106080
timestamp 1586547711
transform 1 0 22756 0 1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1586547711
transform 1 0 22848 0 1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL115920x108800
timestamp 1586547711
transform 1 0 23584 0 -1 22704
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1212
timestamp 1586547711
transform 1 0 25240 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1205
timestamp 1586547711
transform 1 0 25424 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1174
timestamp 1586547711
transform 1 0 25608 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_266
timestamp 1586547711
transform 1 0 25792 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL126040x108800
timestamp 1586547711
transform 1 0 25608 0 -1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL123740x106080
timestamp 1586547711
transform 1 0 25148 0 1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1586547711
transform 1 0 25700 0 -1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL124200x108800
timestamp 1586547711
transform 1 0 25240 0 -1 22704
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_969
timestamp 1586547711
transform 1 0 25976 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1173
timestamp 1586547711
transform 1 0 26160 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _629_
timestamp 1586547711
transform 1 0 26344 0 1 21616
box 0 -48 644 592
use sky130_fd_sc_hd__a32oi_4  _641_
timestamp 1586547711
transform 1 0 25792 0 -1 22704
box 0 -48 2024 592
use sky130_fd_sc_hd__decap_12  FILL134780x106080
timestamp 1586547711
transform 1 0 27356 0 1 21616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL137080x108800
timestamp 1586547711
transform 1 0 27816 0 -1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_197
timestamp 1586547711
transform 1 0 26988 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1168
timestamp 1586547711
transform 1 0 27172 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL143520x106080
timestamp 1586547711
transform 1 0 29104 0 1 21616
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_275
timestamp 1586547711
transform 1 0 28552 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1210
timestamp 1586547711
transform 1 0 28736 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1240
timestamp 1586547711
transform 1 0 28920 0 1 21616
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1586547711
transform 1 0 28460 0 1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _658_
timestamp 1586547711
transform 1 0 28552 0 -1 22704
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL143980x108800
timestamp 1586547711
transform 1 0 29196 0 -1 22704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL149040x106080
timestamp 1586547711
transform 1 0 30208 0 1 21616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL153180x108800
timestamp 1586547711
transform 1 0 31036 0 -1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL149500x108800
timestamp 1586547711
transform 1 0 30300 0 -1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL154560x106080
timestamp 1586547711
transform 1 0 31312 0 1 21616
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1586547711
transform 1 0 31312 0 -1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1586547711
transform 1 0 31404 0 -1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1586547711
transform 1 0 31404 0 1 21616
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1586547711
transform 1 0 400 0 1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__dfrtp_4  _920_
timestamp 1586547711
transform 1 0 676 0 1 22704
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_8  FILL20700x111520
timestamp 1586547711
transform 1 0 4540 0 1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1298
timestamp 1586547711
transform 1 0 2976 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_644
timestamp 1586547711
transform 1 0 3160 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_208
timestamp 1586547711
transform 1 0 3344 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_209
timestamp 1586547711
transform 1 0 4172 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1295
timestamp 1586547711
transform 1 0 4356 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL11960x111520
timestamp 1586547711
transform 1 0 2792 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _680_
timestamp 1586547711
transform 1 0 3528 0 1 22704
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1281
timestamp 1586547711
transform 1 0 5460 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_610
timestamp 1586547711
transform 1 0 5644 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_428
timestamp 1586547711
transform 1 0 5828 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1586547711
transform 1 0 6012 0 1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL24380x111520
timestamp 1586547711
transform 1 0 5276 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__o22ai_4  _673_
timestamp 1586547711
transform 1 0 6104 0 1 22704
box 0 -48 1472 592
use sky130_fd_sc_hd__decap_12  FILL36800x111520
timestamp 1586547711
transform 1 0 7760 0 1 22704
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_531
timestamp 1586547711
transform 1 0 7576 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_672
timestamp 1586547711
transform 1 0 9048 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_674
timestamp 1586547711
transform 1 0 9232 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL42320x111520
timestamp 1586547711
transform 1 0 8864 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL45080x111520
timestamp 1586547711
transform 1 0 9416 0 1 22704
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_410
timestamp 1586547711
transform 1 0 10520 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_544
timestamp 1586547711
transform 1 0 10704 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_570
timestamp 1586547711
transform 1 0 10888 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_585
timestamp 1586547711
transform 1 0 11072 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_609
timestamp 1586547711
transform 1 0 11256 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL55200x111520
timestamp 1586547711
transform 1 0 11440 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL65320x111520
timestamp 1586547711
transform 1 0 13464 0 1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_529
timestamp 1586547711
transform 1 0 11808 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_320
timestamp 1586547711
transform 1 0 11992 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL56580x111520
timestamp 1586547711
transform 1 0 11716 0 1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1586547711
transform 1 0 11624 0 1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _472_
timestamp 1586547711
transform 1 0 12176 0 1 22704
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL73600x111520
timestamp 1586547711
transform 1 0 15120 0 1 22704
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1693
timestamp 1586547711
transform 1 0 14752 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1698
timestamp 1586547711
transform 1 0 14936 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_4  _CTS_buf_1_64
timestamp 1586547711
transform 1 0 14200 0 1 22704
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILL82800x111520
timestamp 1586547711
transform 1 0 16960 0 1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL79120x111520
timestamp 1586547711
transform 1 0 16224 0 1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_513
timestamp 1586547711
transform 1 0 17880 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_477
timestamp 1586547711
transform 1 0 18064 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1586547711
transform 1 0 17236 0 1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL84640x111520
timestamp 1586547711
transform 1 0 17328 0 1 22704
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_312
timestamp 1586547711
transform 1 0 18248 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_304
timestamp 1586547711
transform 1 0 18432 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _893_
timestamp 1586547711
transform 1 0 18616 0 1 22704
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1071
timestamp 1586547711
transform 1 0 21192 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_960
timestamp 1586547711
transform 1 0 21376 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_958
timestamp 1586547711
transform 1 0 22112 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_959
timestamp 1586547711
transform 1 0 22296 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL103500x111520
timestamp 1586547711
transform 1 0 21100 0 1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL101660x111520
timestamp 1586547711
transform 1 0 20732 0 1 22704
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILL110400x111520
timestamp 1586547711
transform 1 0 22480 0 1 22704
box 0 -48 368 592
use sky130_fd_sc_hd__buf_4  _553_
timestamp 1586547711
transform 1 0 21560 0 1 22704
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_257
timestamp 1586547711
transform 1 0 22940 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_962
timestamp 1586547711
transform 1 0 23124 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1069
timestamp 1586547711
transform 1 0 23308 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1073
timestamp 1586547711
transform 1 0 23584 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_963
timestamp 1586547711
transform 1 0 23768 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL115460x111520
timestamp 1586547711
transform 1 0 23492 0 1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1586547711
transform 1 0 22848 0 1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _625_
timestamp 1586547711
transform 1 0 23952 0 1 22704
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1353
timestamp 1586547711
transform 1 0 25792 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_514
timestamp 1586547711
transform 1 0 26528 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_272
timestamp 1586547711
transform 1 0 26804 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL131560x111520
timestamp 1586547711
transform 1 0 26712 0 1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL124200x111520
timestamp 1586547711
transform 1 0 25240 0 1 22704
box 0 -48 552 592
use sky130_fd_sc_hd__buf_4  _419_
timestamp 1586547711
transform 1 0 25976 0 1 22704
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL140760x111520
timestamp 1586547711
transform 1 0 28552 0 1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_965
timestamp 1586547711
transform 1 0 26988 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1209
timestamp 1586547711
transform 1 0 27172 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1229
timestamp 1586547711
transform 1 0 27356 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1235
timestamp 1586547711
transform 1 0 27540 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1236
timestamp 1586547711
transform 1 0 27724 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1586547711
transform 1 0 28460 0 1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL137540x111520
timestamp 1586547711
transform 1 0 27908 0 1 22704
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILL144440x111520
timestamp 1586547711
transform 1 0 29288 0 1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL150880x111520
timestamp 1586547711
transform 1 0 30576 0 1 22704
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_193
timestamp 1586547711
transform 1 0 29564 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_174
timestamp 1586547711
transform 1 0 30024 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1171
timestamp 1586547711
transform 1 0 30208 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1228
timestamp 1586547711
transform 1 0 30392 0 1 22704
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL154560x111520
timestamp 1586547711
transform 1 0 31312 0 1 22704
box 0 -48 92 592
use sky130_fd_sc_hd__conb_1  _840_
timestamp 1586547711
transform 1 0 29748 0 1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1586547711
transform 1 0 31404 0 1 22704
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1586547711
transform 1 0 400 0 -1 23792
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL9200x114240
timestamp 1586547711
transform 1 0 2240 0 -1 23792
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_210
timestamp 1586547711
transform 1 0 676 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1543
timestamp 1586547711
transform 1 0 860 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1257
timestamp 1586547711
transform 1 0 2056 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL3220x114240
timestamp 1586547711
transform 1 0 1044 0 -1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL6440x114240
timestamp 1586547711
transform 1 0 1688 0 -1 23792
box 0 -48 368 592
use sky130_fd_sc_hd__buf_4  _820_
timestamp 1586547711
transform 1 0 1136 0 -1 23792
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL17020x114240
timestamp 1586547711
transform 1 0 3804 0 -1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL12880x114240
timestamp 1586547711
transform 1 0 2976 0 -1 23792
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1586547711
transform 1 0 3252 0 -1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _458_
timestamp 1586547711
transform 1 0 3344 0 -1 23792
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL22540x114240
timestamp 1586547711
transform 1 0 4908 0 -1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_678
timestamp 1586547711
transform 1 0 6104 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL28060x114240
timestamp 1586547711
transform 1 0 6012 0 -1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL29440x114240
timestamp 1586547711
transform 1 0 6288 0 -1 23792
box 0 -48 552 592
use sky130_fd_sc_hd__buf_4  _434_
timestamp 1586547711
transform 1 0 6840 0 -1 23792
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL37720x114240
timestamp 1586547711
transform 1 0 7944 0 -1 23792
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1538
timestamp 1586547711
transform 1 0 7576 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1603
timestamp 1586547711
transform 1 0 7760 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL42780x114240
timestamp 1586547711
transform 1 0 8956 0 -1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1586547711
transform 1 0 8864 0 -1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL34960x114240
timestamp 1586547711
transform 1 0 7392 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL41400x114240
timestamp 1586547711
transform 1 0 8680 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _465_
timestamp 1586547711
transform 1 0 9048 0 -1 23792
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL46000x114240
timestamp 1586547711
transform 1 0 9600 0 -1 23792
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILL49680x114240
timestamp 1586547711
transform 1 0 10336 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__o22ai_4  _451_
timestamp 1586547711
transform 1 0 10520 0 -1 23792
box 0 -48 1472 592
use sky130_fd_sc_hd__decap_12  FILL64860x114240
timestamp 1586547711
transform 1 0 13372 0 -1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_673
timestamp 1586547711
transform 1 0 12176 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_700
timestamp 1586547711
transform 1 0 12360 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1692
timestamp 1586547711
transform 1 0 13188 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL63480x114240
timestamp 1586547711
transform 1 0 13096 0 -1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL60720x114240
timestamp 1586547711
transform 1 0 12544 0 -1 23792
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILL57960x114240
timestamp 1586547711
transform 1 0 11992 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL70840x114240
timestamp 1586547711
transform 1 0 14568 0 -1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL76360x114240
timestamp 1586547711
transform 1 0 15672 0 -1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1586547711
transform 1 0 14476 0 -1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL81880x114240
timestamp 1586547711
transform 1 0 16776 0 -1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILL87400x114240
timestamp 1586547711
transform 1 0 17880 0 -1 23792
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL98900x114240
timestamp 1586547711
transform 1 0 20180 0 -1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL93840x114240
timestamp 1586547711
transform 1 0 19168 0 -1 23792
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL90160x114240
timestamp 1586547711
transform 1 0 18432 0 -1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1586547711
transform 1 0 20088 0 -1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL97520x114240
timestamp 1586547711
transform 1 0 19904 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _418_
timestamp 1586547711
transform 1 0 18524 0 -1 23792
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  FILL104420x114240
timestamp 1586547711
transform 1 0 21284 0 -1 23792
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL108100x114240
timestamp 1586547711
transform 1 0 22020 0 -1 23792
box 0 -48 736 592
use sky130_fd_sc_hd__inv_4  _589_
timestamp 1586547711
transform 1 0 21560 0 -1 23792
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL119600x114240
timestamp 1586547711
transform 1 0 24320 0 -1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1160
timestamp 1586547711
transform 1 0 23952 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1163
timestamp 1586547711
transform 1 0 24136 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL115920x114240
timestamp 1586547711
transform 1 0 23584 0 -1 23792
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILL111780x114240
timestamp 1586547711
transform 1 0 22756 0 -1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _588_
timestamp 1586547711
transform 1 0 22940 0 -1 23792
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  FILL125120x114240
timestamp 1586547711
transform 1 0 25424 0 -1 23792
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL130640x114240
timestamp 1586547711
transform 1 0 26528 0 -1 23792
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL126960x114240
timestamp 1586547711
transform 1 0 25792 0 -1 23792
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1586547711
transform 1 0 25700 0 -1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__a32oi_4  _655_
timestamp 1586547711
transform 1 0 26804 0 -1 23792
box 0 -48 2024 592
use sky130_fd_sc_hd__decap_8  FILL142140x114240
timestamp 1586547711
transform 1 0 28828 0 -1 23792
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILL149040x114240
timestamp 1586547711
transform 1 0 30208 0 -1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1586547711
transform 1 0 31312 0 -1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _651_
timestamp 1586547711
transform 1 0 29564 0 -1 23792
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1586547711
transform 1 0 31404 0 -1 23792
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1586547711
transform 1 0 400 0 1 23792
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL1380x116960
timestamp 1586547711
transform 1 0 676 0 1 23792
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1305
timestamp 1586547711
transform 1 0 1504 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_611
timestamp 1586547711
transform 1 0 1688 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_432
timestamp 1586547711
transform 1 0 1872 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL5060x116960
timestamp 1586547711
transform 1 0 1412 0 1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__o22ai_4  _683_
timestamp 1586547711
transform 1 0 2056 0 1 23792
box 0 -48 1472 592
use sky130_fd_sc_hd__decap_12  FILL19780x116960
timestamp 1586547711
transform 1 0 4356 0 1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_659
timestamp 1586547711
transform 1 0 3620 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1270
timestamp 1586547711
transform 1 0 3804 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1302
timestamp 1586547711
transform 1 0 3988 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1306
timestamp 1586547711
transform 1 0 4172 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL15640x116960
timestamp 1586547711
transform 1 0 3528 0 1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILL28520x116960
timestamp 1586547711
transform 1 0 6104 0 1 23792
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1681
timestamp 1586547711
transform 1 0 6380 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_429
timestamp 1586547711
transform 1 0 6564 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_204
timestamp 1586547711
transform 1 0 6748 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1586547711
transform 1 0 6012 0 1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL25300x116960
timestamp 1586547711
transform 1 0 5460 0 1 23792
box 0 -48 552 592
use sky130_fd_sc_hd__dfrtp_4  _918_
timestamp 1586547711
transform 1 0 6932 0 1 23792
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA_203
timestamp 1586547711
transform 1 0 9232 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL43240x116960
timestamp 1586547711
transform 1 0 9048 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL51520x116960
timestamp 1586547711
transform 1 0 10704 0 1 23792
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_671
timestamp 1586547711
transform 1 0 9416 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_604
timestamp 1586547711
transform 1 0 10336 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1282
timestamp 1586547711
transform 1 0 10520 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL46000x116960
timestamp 1586547711
transform 1 0 9600 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL55200x116960
timestamp 1586547711
transform 1 0 11440 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _674_
timestamp 1586547711
transform 1 0 9784 0 1 23792
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_527
timestamp 1586547711
transform 1 0 12268 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_530
timestamp 1586547711
transform 1 0 12452 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_411
timestamp 1586547711
transform 1 0 12820 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_321
timestamp 1586547711
transform 1 0 13004 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1586547711
transform 1 0 11624 0 1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _928_
timestamp 1586547711
transform 1 0 13188 0 1 23792
box 0 -48 2116 592
use sky130_fd_sc_hd__fill_2  FILL61180x116960
timestamp 1586547711
transform 1 0 12636 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _433_
timestamp 1586547711
transform 1 0 11716 0 1 23792
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILL74520x116960
timestamp 1586547711
transform 1 0 15304 0 1 23792
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_699
timestamp 1586547711
transform 1 0 15580 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1381
timestamp 1586547711
transform 1 0 15764 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL78660x116960
timestamp 1586547711
transform 1 0 16132 0 1 23792
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1383
timestamp 1586547711
transform 1 0 15948 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_305
timestamp 1586547711
transform 1 0 16960 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL82340x116960
timestamp 1586547711
transform 1 0 16868 0 1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL87400x116960
timestamp 1586547711
transform 1 0 17880 0 1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_454
timestamp 1586547711
transform 1 0 17328 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1382
timestamp 1586547711
transform 1 0 17512 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1384
timestamp 1586547711
transform 1 0 17696 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL83720x116960
timestamp 1586547711
transform 1 0 17144 0 1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1586547711
transform 1 0 17236 0 1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILL92920x116960
timestamp 1586547711
transform 1 0 18984 0 1 23792
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL98900x116960
timestamp 1586547711
transform 1 0 20180 0 1 23792
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_481
timestamp 1586547711
transform 1 0 19812 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1448
timestamp 1586547711
transform 1 0 19996 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _788_
timestamp 1586547711
transform 1 0 19260 0 1 23792
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL106260x116960
timestamp 1586547711
transform 1 0 21652 0 1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_258
timestamp 1586547711
transform 1 0 20916 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_413
timestamp 1586547711
transform 1 0 21100 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_497
timestamp 1586547711
transform 1 0 21284 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1457
timestamp 1586547711
transform 1 0 21468 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL112700x116960
timestamp 1586547711
transform 1 0 22940 0 1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL118220x116960
timestamp 1586547711
transform 1 0 24044 0 1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL111780x116960
timestamp 1586547711
transform 1 0 22756 0 1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1586547711
transform 1 0 22848 0 1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILL132480x116960
timestamp 1586547711
transform 1 0 26896 0 1 23792
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL128800x116960
timestamp 1586547711
transform 1 0 26160 0 1 23792
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_515
timestamp 1586547711
transform 1 0 25792 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1059
timestamp 1586547711
transform 1 0 25976 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL126500x116960
timestamp 1586547711
transform 1 0 25700 0 1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL123740x116960
timestamp 1586547711
transform 1 0 25148 0 1 23792
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILL140760x116960
timestamp 1586547711
transform 1 0 28552 0 1 23792
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_420
timestamp 1586547711
transform 1 0 27172 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1110
timestamp 1586547711
transform 1 0 27356 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1213
timestamp 1586547711
transform 1 0 27540 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1215
timestamp 1586547711
transform 1 0 27724 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1356
timestamp 1586547711
transform 1 0 27908 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1586547711
transform 1 0 28460 0 1 23792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL138460x116960
timestamp 1586547711
transform 1 0 28092 0 1 23792
box 0 -48 368 592
use sky130_fd_sc_hd__inv_4  _642_
timestamp 1586547711
transform 1 0 28828 0 1 23792
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL148120x116960
timestamp 1586547711
transform 1 0 30024 0 1 23792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL153640x116960
timestamp 1586547711
transform 1 0 31128 0 1 23792
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_268
timestamp 1586547711
transform 1 0 29288 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1214
timestamp 1586547711
transform 1 0 29472 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1478
timestamp 1586547711
transform 1 0 29656 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1582
timestamp 1586547711
transform 1 0 29840 0 1 23792
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1586547711
transform 1 0 31404 0 1 23792
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1586547711
transform 1 0 400 0 -1 24880
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL5060x119680
timestamp 1586547711
transform 1 0 1412 0 -1 24880
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL1380x119680
timestamp 1586547711
transform 1 0 676 0 -1 24880
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL9200x119680
timestamp 1586547711
transform 1 0 2240 0 -1 24880
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1284
timestamp 1586547711
transform 1 0 1688 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_648
timestamp 1586547711
transform 1 0 2056 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL7360x119680
timestamp 1586547711
transform 1 0 1872 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL21620x119680
timestamp 1586547711
transform 1 0 4724 0 -1 24880
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL12880x119680
timestamp 1586547711
transform 1 0 2976 0 -1 24880
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1312
timestamp 1586547711
transform 1 0 3344 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL15640x119680
timestamp 1586547711
transform 1 0 3528 0 -1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1586547711
transform 1 0 3252 0 -1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__o21a_4  _684_
timestamp 1586547711
transform 1 0 3620 0 -1 24880
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL27140x119680
timestamp 1586547711
transform 1 0 5828 0 -1 24880
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1539
timestamp 1586547711
transform 1 0 6932 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILL42780x119680
timestamp 1586547711
transform 1 0 8956 0 -1 24880
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL38640x119680
timestamp 1586547711
transform 1 0 8128 0 -1 24880
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL35420x119680
timestamp 1586547711
transform 1 0 7484 0 -1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1586547711
transform 1 0 8864 0 -1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL33580x119680
timestamp 1586547711
transform 1 0 7116 0 -1 24880
box 0 -48 368 592
use sky130_fd_sc_hd__buf_4  _818_
timestamp 1586547711
transform 1 0 7576 0 -1 24880
box 0 -48 552 592
use sky130_fd_sc_hd__inv_4  _464_
timestamp 1586547711
transform 1 0 9232 0 -1 24880
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL46460x119680
timestamp 1586547711
transform 1 0 9692 0 -1 24880
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL51980x119680
timestamp 1586547711
transform 1 0 10796 0 -1 24880
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL57500x119680
timestamp 1586547711
transform 1 0 11900 0 -1 24880
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL64860x119680
timestamp 1586547711
transform 1 0 13372 0 -1 24880
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_485
timestamp 1586547711
transform 1 0 13188 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL63020x119680
timestamp 1586547711
transform 1 0 13004 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILL74520x119680
timestamp 1586547711
transform 1 0 15304 0 -1 24880
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL70840x119680
timestamp 1586547711
transform 1 0 14568 0 -1 24880
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1586547711
transform 1 0 14476 0 -1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _719_
timestamp 1586547711
transform 1 0 15580 0 -1 24880
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL79120x119680
timestamp 1586547711
transform 1 0 16224 0 -1 24880
box 0 -48 736 592
use sky130_fd_sc_hd__a21bo_4  _720_ ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 16960 0 -1 24880
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_12  FILL90620x119680
timestamp 1586547711
transform 1 0 18524 0 -1 24880
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL98900x119680
timestamp 1586547711
transform 1 0 20180 0 -1 24880
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_550
timestamp 1586547711
transform 1 0 18156 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_957
timestamp 1586547711
transform 1 0 18340 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL97980x119680
timestamp 1586547711
transform 1 0 19996 0 -1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1586547711
transform 1 0 20088 0 -1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL96140x119680
timestamp 1586547711
transform 1 0 19628 0 -1 24880
box 0 -48 368 592
use sky130_fd_sc_hd__dfrtp_4  _894_
timestamp 1586547711
transform 1 0 20916 0 -1 24880
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_12  FILL117300x119680
timestamp 1586547711
transform 1 0 23860 0 -1 24880
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1150
timestamp 1586547711
transform 1 0 23676 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL115920x119680
timestamp 1586547711
transform 1 0 23584 0 -1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL113160x119680
timestamp 1586547711
transform 1 0 23032 0 -1 24880
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL122820x119680
timestamp 1586547711
transform 1 0 24964 0 -1 24880
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL129260x119680
timestamp 1586547711
transform 1 0 26252 0 -1 24880
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1586547711
transform 1 0 25700 0 -1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _585_
timestamp 1586547711
transform 1 0 25792 0 -1 24880
box 0 -48 460 592
use sky130_fd_sc_hd__decap_8  FILL142140x119680
timestamp 1586547711
transform 1 0 28828 0 -1 24880
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1469
timestamp 1586547711
transform 1 0 28644 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL132940x119680
timestamp 1586547711
transform 1 0 26988 0 -1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__o22ai_4  _643_
timestamp 1586547711
transform 1 0 27172 0 -1 24880
box 0 -48 1472 592
use sky130_fd_sc_hd__decap_12  FILL148580x119680
timestamp 1586547711
transform 1 0 30116 0 -1 24880
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL154100x119680
timestamp 1586547711
transform 1 0 31220 0 -1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1586547711
transform 1 0 31312 0 -1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _797_
timestamp 1586547711
transform 1 0 29564 0 -1 24880
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1586547711
transform 1 0 31404 0 -1 24880
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1586547711
transform 1 0 400 0 1 24880
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1315
timestamp 1586547711
transform 1 0 1136 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_661
timestamp 1586547711
transform 1 0 1320 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_434
timestamp 1586547711
transform 1 0 1504 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL3220x122400
timestamp 1586547711
transform 1 0 1044 0 1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL1380x122400
timestamp 1586547711
transform 1 0 676 0 1 24880
box 0 -48 368 592
use sky130_fd_sc_hd__o22ai_4  _688_
timestamp 1586547711
transform 1 0 1688 0 1 24880
box 0 -48 1472 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1308
timestamp 1586547711
transform 1 0 3160 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_539
timestamp 1586547711
transform 1 0 3344 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_649
timestamp 1586547711
transform 1 0 3528 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1307
timestamp 1586547711
transform 1 0 3712 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_660
timestamp 1586547711
transform 1 0 4540 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1303
timestamp 1586547711
transform 1 0 4724 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _685_
timestamp 1586547711
transform 1 0 3896 0 1 24880
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1314
timestamp 1586547711
transform 1 0 4908 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_542
timestamp 1586547711
transform 1 0 5552 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_537
timestamp 1586547711
transform 1 0 5736 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL25300x122400
timestamp 1586547711
transform 1 0 5460 0 1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL27600x122400
timestamp 1586547711
transform 1 0 5920 0 1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL23460x122400
timestamp 1586547711
transform 1 0 5092 0 1 24880
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL33120x122400
timestamp 1586547711
transform 1 0 7024 0 1 24880
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1269
timestamp 1586547711
transform 1 0 6656 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1274
timestamp 1586547711
transform 1 0 6840 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1586547711
transform 1 0 6012 0 1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _671_
timestamp 1586547711
transform 1 0 6104 0 1 24880
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL38640x122400
timestamp 1586547711
transform 1 0 8128 0 1 24880
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL44160x122400
timestamp 1586547711
transform 1 0 9232 0 1 24880
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_603
timestamp 1586547711
transform 1 0 10888 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_608
timestamp 1586547711
transform 1 0 11072 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL54280x122400
timestamp 1586547711
transform 1 0 11256 0 1 24880
box 0 -48 368 592
use sky130_fd_sc_hd__buf_4  _450_
timestamp 1586547711
transform 1 0 10336 0 1 24880
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILL58420x122400
timestamp 1586547711
transform 1 0 12084 0 1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1586547711
transform 1 0 11624 0 1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL56580x122400
timestamp 1586547711
transform 1 0 11716 0 1 24880
box 0 -48 368 592
use sky130_fd_sc_hd__inv_4  _432_
timestamp 1586547711
transform 1 0 12176 0 1 24880
box 0 -48 460 592
use sky130_fd_sc_hd__diode_2  ANTENNA_317
timestamp 1586547711
transform 1 0 12636 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_526
timestamp 1586547711
transform 1 0 12820 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1699
timestamp 1586547711
transform 1 0 13096 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_42
timestamp 1586547711
transform 1 0 13280 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL63020x122400
timestamp 1586547711
transform 1 0 13004 0 1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_16  _CTS_root ${PDK_PATH}/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1586547711
transform 1 0 13464 0 1 24880
box 0 -48 1840 592
use sky130_fd_sc_hd__fill_1  FILL77280x122400
timestamp 1586547711
transform 1 0 15856 0 1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL74520x122400
timestamp 1586547711
transform 1 0 15304 0 1 24880
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1380
timestamp 1586547711
transform 1 0 15948 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_236
timestamp 1586547711
transform 1 0 16132 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_241
timestamp 1586547711
transform 1 0 16316 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_606
timestamp 1586547711
transform 1 0 16500 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_955
timestamp 1586547711
transform 1 0 16684 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_455
timestamp 1586547711
transform 1 0 16868 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_306
timestamp 1586547711
transform 1 0 17052 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1586547711
transform 1 0 17236 0 1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _913_
timestamp 1586547711
transform 1 0 17328 0 1 24880
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1456
timestamp 1586547711
transform 1 0 19904 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_525
timestamp 1586547711
transform 1 0 20088 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL97060x122400
timestamp 1586547711
transform 1 0 19812 0 1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL95220x122400
timestamp 1586547711
transform 1 0 19444 0 1 24880
box 0 -48 368 592
use sky130_fd_sc_hd__buf_4  _789_
timestamp 1586547711
transform 1 0 20272 0 1 24880
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_482
timestamp 1586547711
transform 1 0 20824 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_498
timestamp 1586547711
transform 1 0 21008 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_495
timestamp 1586547711
transform 1 0 21192 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_483
timestamp 1586547711
transform 1 0 21376 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_261
timestamp 1586547711
transform 1 0 22112 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_415
timestamp 1586547711
transform 1 0 22296 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1460
timestamp 1586547711
transform 1 0 22480 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _790_
timestamp 1586547711
transform 1 0 21560 0 1 24880
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1461
timestamp 1586547711
transform 1 0 22664 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1355
timestamp 1586547711
transform 1 0 23124 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_416
timestamp 1586547711
transform 1 0 23308 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_262
timestamp 1586547711
transform 1 0 23492 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1586547711
transform 1 0 22848 0 1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _618_
timestamp 1586547711
transform 1 0 23676 0 1 24880
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILL112700x122400
timestamp 1586547711
transform 1 0 22940 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_263
timestamp 1586547711
transform 1 0 24964 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1161
timestamp 1586547711
transform 1 0 25148 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1060
timestamp 1586547711
transform 1 0 26344 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1063
timestamp 1586547711
transform 1 0 26528 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1061
timestamp 1586547711
transform 1 0 26712 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1225
timestamp 1586547711
transform 1 0 26896 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL126500x122400
timestamp 1586547711
transform 1 0 25700 0 1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL124660x122400
timestamp 1586547711
transform 1 0 25332 0 1 24880
box 0 -48 368 592
use sky130_fd_sc_hd__buf_4  _586_
timestamp 1586547711
transform 1 0 25792 0 1 24880
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1226
timestamp 1586547711
transform 1 0 27080 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1617
timestamp 1586547711
transform 1 0 27724 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_488
timestamp 1586547711
transform 1 0 27908 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_421
timestamp 1586547711
transform 1 0 28092 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_270
timestamp 1586547711
transform 1 0 28276 0 1 24880
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL136160x122400
timestamp 1586547711
transform 1 0 27632 0 1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1586547711
transform 1 0 28460 0 1 24880
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL134320x122400
timestamp 1586547711
transform 1 0 27264 0 1 24880
box 0 -48 368 592
use sky130_fd_sc_hd__dfrtp_4  _898_
timestamp 1586547711
transform 1 0 28552 0 1 24880
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_8  FILL151340x122400
timestamp 1586547711
transform 1 0 30668 0 1 24880
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1586547711
transform 1 0 31404 0 1 24880
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL7360x125120
timestamp 1586547711
transform 1 0 1872 0 -1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1586547711
transform 1 0 400 0 1 25968
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1586547711
transform 1 0 400 0 -1 25968
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_435
timestamp 1586547711
transform 1 0 676 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1684
timestamp 1586547711
transform 1 0 860 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1258
timestamp 1586547711
transform 1 0 1688 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL5980x125120
timestamp 1586547711
transform 1 0 1596 0 -1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL3220x125120
timestamp 1586547711
transform 1 0 1044 0 -1 25968
box 0 -48 552 592
use sky130_fd_sc_hd__dfrtp_4  _921_
timestamp 1586547711
transform 1 0 676 0 1 25968
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_3  FILL12880x125120
timestamp 1586547711
transform 1 0 2976 0 -1 25968
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1309
timestamp 1586547711
transform 1 0 3344 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1311
timestamp 1586547711
transform 1 0 3528 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1586547711
transform 1 0 3252 0 -1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL11960x127840
timestamp 1586547711
transform 1 0 2792 0 1 25968
box 0 -48 552 592
use sky130_fd_sc_hd__decap_6  FILL16560x127840
timestamp 1586547711
transform 1 0 3712 0 1 25968
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL21160x125120
timestamp 1586547711
transform 1 0 4632 0 -1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_211
timestamp 1586547711
transform 1 0 4724 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _461_
timestamp 1586547711
transform 1 0 4264 0 1 25968
box 0 -48 460 592
use sky130_fd_sc_hd__o22a_4  _687_
timestamp 1586547711
transform 1 0 3344 0 -1 25968
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA_657
timestamp 1586547711
transform 1 0 4908 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_687
timestamp 1586547711
transform 1 0 5644 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_319
timestamp 1586547711
transform 1 0 5828 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL23460x127840
timestamp 1586547711
transform 1 0 5092 0 1 25968
box 0 -48 552 592
use sky130_fd_sc_hd__buf_4  _435_
timestamp 1586547711
transform 1 0 5736 0 -1 25968
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL32660x125120
timestamp 1586547711
transform 1 0 6932 0 -1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL29440x125120
timestamp 1586547711
transform 1 0 6288 0 -1 25968
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_212
timestamp 1586547711
transform 1 0 6748 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_214
timestamp 1586547711
transform 1 0 6932 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_691
timestamp 1586547711
transform 1 0 6564 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_693
timestamp 1586547711
transform 1 0 6748 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1586547711
transform 1 0 6012 0 1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _468_
timestamp 1586547711
transform 1 0 6104 0 1 25968
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_218
timestamp 1586547711
transform 1 0 7116 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_688
timestamp 1586547711
transform 1 0 7300 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1363
timestamp 1586547711
transform 1 0 8036 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL35420x127840
timestamp 1586547711
transform 1 0 7484 0 1 25968
box 0 -48 552 592
use sky130_fd_sc_hd__decap_6  FILL38180x125120
timestamp 1586547711
transform 1 0 8036 0 -1 25968
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILL42780x125120
timestamp 1586547711
transform 1 0 8956 0 -1 25968
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1279
timestamp 1586547711
transform 1 0 8220 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_228
timestamp 1586547711
transform 1 0 8404 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1362
timestamp 1586547711
transform 1 0 8588 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_624
timestamp 1586547711
transform 1 0 9232 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL41860x125120
timestamp 1586547711
transform 1 0 8772 0 -1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1586547711
transform 1 0 8864 0 -1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__a211o_4  _707_
timestamp 1586547711
transform 1 0 8588 0 1 25968
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILL50140x127840
timestamp 1586547711
transform 1 0 10428 0 1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL46920x125120
timestamp 1586547711
transform 1 0 9784 0 -1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL52440x125120
timestamp 1586547711
transform 1 0 10888 0 -1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_229
timestamp 1586547711
transform 1 0 9876 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_442
timestamp 1586547711
transform 1 0 10060 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1364
timestamp 1586547711
transform 1 0 10244 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_692
timestamp 1586547711
transform 1 0 9416 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1286
timestamp 1586547711
transform 1 0 9600 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL61180x127840
timestamp 1586547711
transform 1 0 12636 0 1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL57960x125120
timestamp 1586547711
transform 1 0 11992 0 -1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL63480x125120
timestamp 1586547711
transform 1 0 13096 0 -1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1571
timestamp 1586547711
transform 1 0 12268 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1612
timestamp 1586547711
transform 1 0 12452 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL55660x127840
timestamp 1586547711
transform 1 0 11532 0 1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1586547711
transform 1 0 11624 0 1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _827_
timestamp 1586547711
transform 1 0 11716 0 1 25968
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILL69000x125120
timestamp 1586547711
transform 1 0 14200 0 -1 25968
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_552
timestamp 1586547711
transform 1 0 13832 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_242
timestamp 1586547711
transform 1 0 14016 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_237
timestamp 1586547711
transform 1 0 14200 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1400
timestamp 1586547711
transform 1 0 14568 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL66700x127840
timestamp 1586547711
transform 1 0 13740 0 1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL71760x125120
timestamp 1586547711
transform 1 0 14752 0 -1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1586547711
transform 1 0 14476 0 -1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL74980x125120
timestamp 1586547711
transform 1 0 15396 0 -1 25968
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_549
timestamp 1586547711
transform 1 0 15672 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_554
timestamp 1586547711
transform 1 0 14844 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_559
timestamp 1586547711
transform 1 0 15028 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_562
timestamp 1586547711
transform 1 0 15212 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL77280x127840
timestamp 1586547711
transform 1 0 15856 0 1 25968
box 0 -48 552 592
use sky130_fd_sc_hd__o22a_4  _726_
timestamp 1586547711
transform 1 0 14384 0 1 25968
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA_555
timestamp 1586547711
transform 1 0 16408 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_560
timestamp 1586547711
transform 1 0 16592 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _718_
timestamp 1586547711
transform 1 0 16132 0 -1 25968
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  FILL82800x127840
timestamp 1586547711
transform 1 0 16960 0 1 25968
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_953
timestamp 1586547711
transform 1 0 16776 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1523
timestamp 1586547711
transform 1 0 17328 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1676
timestamp 1586547711
transform 1 0 17512 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1586547711
transform 1 0 17236 0 1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL84640x127840
timestamp 1586547711
transform 1 0 17328 0 1 25968
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILL82800x125120
timestamp 1586547711
transform 1 0 16960 0 -1 25968
box 0 -48 368 592
use sky130_fd_sc_hd__buf_4  _812_
timestamp 1586547711
transform 1 0 17696 0 1 25968
box 0 -48 552 592
use sky130_fd_sc_hd__and2_4  _552_
timestamp 1586547711
transform 1 0 17696 0 -1 25968
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL91080x127840
timestamp 1586547711
transform 1 0 18616 0 1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL90620x125120
timestamp 1586547711
transform 1 0 18524 0 -1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1522
timestamp 1586547711
transform 1 0 18248 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1597
timestamp 1586547711
transform 1 0 18432 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_954
timestamp 1586547711
transform 1 0 18340 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL96600x127840
timestamp 1586547711
transform 1 0 19720 0 1 25968
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL97980x125120
timestamp 1586547711
transform 1 0 19996 0 -1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1586547711
transform 1 0 20088 0 -1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL96140x125120
timestamp 1586547711
transform 1 0 19628 0 -1 25968
box 0 -48 368 592
use sky130_fd_sc_hd__buf_4  _431_
timestamp 1586547711
transform 1 0 20180 0 -1 25968
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL101660x125120
timestamp 1586547711
transform 1 0 20732 0 -1 25968
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_524
timestamp 1586547711
transform 1 0 20548 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_494
timestamp 1586547711
transform 1 0 21284 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL100280x127840
timestamp 1586547711
transform 1 0 20456 0 1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _430_
timestamp 1586547711
transform 1 0 20732 0 1 25968
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL107180x127840
timestamp 1586547711
transform 1 0 21836 0 1 25968
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_496
timestamp 1586547711
transform 1 0 21468 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_523
timestamp 1586547711
transform 1 0 21652 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL105340x125120
timestamp 1586547711
transform 1 0 21468 0 -1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _895_
timestamp 1586547711
transform 1 0 21560 0 -1 25968
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_12  FILL112700x127840
timestamp 1586547711
transform 1 0 22940 0 1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL110860x127840
timestamp 1586547711
transform 1 0 22572 0 1 25968
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1586547711
transform 1 0 22848 0 1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1165
timestamp 1586547711
transform 1 0 24504 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1108
timestamp 1586547711
transform 1 0 23676 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL120060x127840
timestamp 1586547711
transform 1 0 24412 0 1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL120060x125120
timestamp 1586547711
transform 1 0 24412 0 -1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL118220x127840
timestamp 1586547711
transform 1 0 24044 0 1 25968
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILL117300x125120
timestamp 1586547711
transform 1 0 23860 0 -1 25968
box 0 -48 552 592
use sky130_fd_sc_hd__inv_4  _624_
timestamp 1586547711
transform 1 0 24504 0 -1 25968
box 0 -48 460 592
use sky130_fd_sc_hd__or2_4  _626_
timestamp 1586547711
transform 1 0 24688 0 1 25968
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL122820x125120
timestamp 1586547711
transform 1 0 24964 0 -1 25968
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1067
timestamp 1586547711
transform 1 0 25332 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL126960x125120
timestamp 1586547711
transform 1 0 25792 0 -1 25968
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1164
timestamp 1586547711
transform 1 0 25516 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1066
timestamp 1586547711
transform 1 0 25792 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1107
timestamp 1586547711
transform 1 0 25976 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL126500x127840
timestamp 1586547711
transform 1 0 25700 0 1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1586547711
transform 1 0 25700 0 -1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL128800x127840
timestamp 1586547711
transform 1 0 26160 0 1 25968
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1238
timestamp 1586547711
transform 1 0 26804 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL131560x127840
timestamp 1586547711
transform 1 0 26712 0 1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL130640x125120
timestamp 1586547711
transform 1 0 26528 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _649_
timestamp 1586547711
transform 1 0 26712 0 -1 25968
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILL134780x125120
timestamp 1586547711
transform 1 0 27356 0 -1 25968
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1062
timestamp 1586547711
transform 1 0 27632 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1237
timestamp 1586547711
transform 1 0 27816 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL138000x127840
timestamp 1586547711
transform 1 0 28000 0 1 25968
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _656_
timestamp 1586547711
transform 1 0 26988 0 1 25968
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL142140x125120
timestamp 1586547711
transform 1 0 28828 0 -1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_194
timestamp 1586547711
transform 1 0 28552 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_200
timestamp 1586547711
transform 1 0 28736 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_489
timestamp 1586547711
transform 1 0 28644 0 -1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL139840x127840
timestamp 1586547711
transform 1 0 28368 0 1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1586547711
transform 1 0 28460 0 1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL142600x127840
timestamp 1586547711
transform 1 0 28920 0 1 25968
box 0 -48 368 592
use sky130_fd_sc_hd__buf_4  _425_
timestamp 1586547711
transform 1 0 28092 0 -1 25968
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL149500x127840
timestamp 1586547711
transform 1 0 30300 0 1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL147660x125120
timestamp 1586547711
transform 1 0 29932 0 -1 25968
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL153180x125120
timestamp 1586547711
transform 1 0 31036 0 -1 25968
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1468
timestamp 1586547711
transform 1 0 29932 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1579
timestamp 1586547711
transform 1 0 30116 0 1 25968
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL144440x127840
timestamp 1586547711
transform 1 0 29288 0 1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1586547711
transform 1 0 31312 0 -1 25968
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _794_
timestamp 1586547711
transform 1 0 29380 0 1 25968
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1586547711
transform 1 0 31404 0 1 25968
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1586547711
transform 1 0 31404 0 -1 25968
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL3220x130560
timestamp 1586547711
transform 1 0 1044 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1586547711
transform 1 0 400 0 -1 27056
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_213
timestamp 1586547711
transform 1 0 676 0 -1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1545
timestamp 1586547711
transform 1 0 860 0 -1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1328
timestamp 1586547711
transform 1 0 2608 0 -1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL10580x130560
timestamp 1586547711
transform 1 0 2516 0 -1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL8740x130560
timestamp 1586547711
transform 1 0 2148 0 -1 27056
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL17020x130560
timestamp 1586547711
transform 1 0 3804 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL13800x130560
timestamp 1586547711
transform 1 0 3160 0 -1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1586547711
transform 1 0 3252 0 -1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL11960x130560
timestamp 1586547711
transform 1 0 2792 0 -1 27056
box 0 -48 368 592
use sky130_fd_sc_hd__inv_4  _686_
timestamp 1586547711
transform 1 0 3344 0 -1 27056
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL22540x130560
timestamp 1586547711
transform 1 0 4908 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILL28060x130560
timestamp 1586547711
transform 1 0 6012 0 -1 27056
box 0 -48 552 592
use sky130_fd_sc_hd__or4_4  _470_
timestamp 1586547711
transform 1 0 6564 0 -1 27056
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  FILL39560x130560
timestamp 1586547711
transform 1 0 8312 0 -1 27056
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL42780x130560
timestamp 1586547711
transform 1 0 8956 0 -1 27056
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL35880x130560
timestamp 1586547711
transform 1 0 7576 0 -1 27056
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1359
timestamp 1586547711
transform 1 0 7392 0 -1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1350
timestamp 1586547711
transform 1 0 8588 0 -1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL41860x130560
timestamp 1586547711
transform 1 0 8772 0 -1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1586547711
transform 1 0 8864 0 -1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__a32o_4  _708_
timestamp 1586547711
transform 1 0 9232 0 -1 27056
box 0 -48 1564 592
use sky130_fd_sc_hd__decap_8  FILL51980x130560
timestamp 1586547711
transform 1 0 10796 0 -1 27056
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILL57500x130560
timestamp 1586547711
transform 1 0 11900 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL63020x130560
timestamp 1586547711
transform 1 0 13004 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_528
timestamp 1586547711
transform 1 0 11716 0 -1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL55660x130560
timestamp 1586547711
transform 1 0 11532 0 -1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILL76360x130560
timestamp 1586547711
transform 1 0 15672 0 -1 27056
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_956
timestamp 1586547711
transform 1 0 14568 0 -1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL71760x130560
timestamp 1586547711
transform 1 0 14752 0 -1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1586547711
transform 1 0 14476 0 -1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL68540x130560
timestamp 1586547711
transform 1 0 14108 0 -1 27056
box 0 -48 368 592
use sky130_fd_sc_hd__or3_4  _439_
timestamp 1586547711
transform 1 0 14844 0 -1 27056
box 0 -48 828 592
use sky130_fd_sc_hd__decap_12  FILL83260x130560
timestamp 1586547711
transform 1 0 17052 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__and2_4  _551_
timestamp 1586547711
transform 1 0 16408 0 -1 27056
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL88780x130560
timestamp 1586547711
transform 1 0 18156 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL94300x130560
timestamp 1586547711
transform 1 0 19260 0 -1 27056
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL98900x130560
timestamp 1586547711
transform 1 0 20180 0 -1 27056
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL97980x130560
timestamp 1586547711
transform 1 0 19996 0 -1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1586547711
transform 1 0 20088 0 -1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL106720x130560
timestamp 1586547711
transform 1 0 21744 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL102580x130560
timestamp 1586547711
transform 1 0 20916 0 -1 27056
box 0 -48 276 592
use sky130_fd_sc_hd__buf_4  _429_
timestamp 1586547711
transform 1 0 21192 0 -1 27056
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL113620x130560
timestamp 1586547711
transform 1 0 23124 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL120520x130560
timestamp 1586547711
transform 1 0 24504 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1463
timestamp 1586547711
transform 1 0 22940 0 -1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1613
timestamp 1586547711
transform 1 0 24320 0 -1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL112240x130560
timestamp 1586547711
transform 1 0 22848 0 -1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL119140x130560
timestamp 1586547711
transform 1 0 24228 0 -1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL129720x130560
timestamp 1586547711
transform 1 0 26344 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL126040x130560
timestamp 1586547711
transform 1 0 25608 0 -1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1586547711
transform 1 0 25700 0 -1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _604_
timestamp 1586547711
transform 1 0 25792 0 -1 27056
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL135240x130560
timestamp 1586547711
transform 1 0 27448 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL142600x130560
timestamp 1586547711
transform 1 0 28920 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__buf_2  _851_
timestamp 1586547711
transform 1 0 28552 0 -1 27056
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL148120x130560
timestamp 1586547711
transform 1 0 30024 0 -1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1586547711
transform 1 0 31312 0 -1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL153640x130560
timestamp 1586547711
transform 1 0 31128 0 -1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1586547711
transform 1 0 31404 0 -1 27056
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1586547711
transform 1 0 400 0 1 27056
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL1380x133280
timestamp 1586547711
transform 1 0 676 0 1 27056
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1606
timestamp 1586547711
transform 1 0 952 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _821_
timestamp 1586547711
transform 1 0 1136 0 1 27056
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1544
timestamp 1586547711
transform 1 0 1688 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1310
timestamp 1586547711
transform 1 0 1872 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1317
timestamp 1586547711
transform 1 0 2056 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1320
timestamp 1586547711
transform 1 0 2240 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_689
timestamp 1586547711
transform 1 0 2424 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _693_
timestamp 1586547711
transform 1 0 2608 0 1 27056
box 0 -48 828 592
use sky130_fd_sc_hd__decap_8  FILL17940x133280
timestamp 1586547711
transform 1 0 3988 0 1 27056
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_216
timestamp 1586547711
transform 1 0 3436 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1313
timestamp 1586547711
transform 1 0 3620 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1324
timestamp 1586547711
transform 1 0 3804 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1271
timestamp 1586547711
transform 1 0 4816 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL21620x133280
timestamp 1586547711
transform 1 0 4724 0 1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1322
timestamp 1586547711
transform 1 0 5000 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1331
timestamp 1586547711
transform 1 0 5184 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1334
timestamp 1586547711
transform 1 0 5368 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL27600x133280
timestamp 1586547711
transform 1 0 5920 0 1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL25760x133280
timestamp 1586547711
transform 1 0 5552 0 1 27056
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1586547711
transform 1 0 6012 0 1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL28520x133280
timestamp 1586547711
transform 1 0 6104 0 1 27056
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1349
timestamp 1586547711
transform 1 0 6656 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_547
timestamp 1586547711
transform 1 0 6840 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_220
timestamp 1586547711
transform 1 0 7024 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_227
timestamp 1586547711
transform 1 0 9232 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__a32oi_4  _704_
timestamp 1586547711
transform 1 0 7208 0 1 27056
box 0 -48 2024 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1339
timestamp 1586547711
transform 1 0 9416 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1361
timestamp 1586547711
transform 1 0 9600 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL46920x133280
timestamp 1586547711
transform 1 0 9784 0 1 27056
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1688
timestamp 1586547711
transform 1 0 10336 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_230
timestamp 1586547711
transform 1 0 10520 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_443
timestamp 1586547711
transform 1 0 10704 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1570
timestamp 1586547711
transform 1 0 10888 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_690
timestamp 1586547711
transform 1 0 11072 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_226
timestamp 1586547711
transform 1 0 11256 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_222
timestamp 1586547711
transform 1 0 11440 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL62100x133280
timestamp 1586547711
transform 1 0 12820 0 1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1586547711
transform 1 0 11624 0 1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__a21o_4  _469_
timestamp 1586547711
transform 1 0 11716 0 1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL67620x133280
timestamp 1586547711
transform 1 0 13924 0 1 27056
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1368
timestamp 1586547711
transform 1 0 14660 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1366
timestamp 1586547711
transform 1 0 14844 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_239
timestamp 1586547711
transform 1 0 15488 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_548
timestamp 1586547711
transform 1 0 15672 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_556
timestamp 1586547711
transform 1 0 15856 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _436_
timestamp 1586547711
transform 1 0 15028 0 1 27056
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL84640x133280
timestamp 1586547711
transform 1 0 17328 0 1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_233
timestamp 1586547711
transform 1 0 16500 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_558
timestamp 1586547711
transform 1 0 16684 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL80040x133280
timestamp 1586547711
transform 1 0 16408 0 1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1586547711
transform 1 0 17236 0 1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL78200x133280
timestamp 1586547711
transform 1 0 16040 0 1 27056
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILL82340x133280
timestamp 1586547711
transform 1 0 16868 0 1 27056
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL90160x133280
timestamp 1586547711
transform 1 0 18432 0 1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_508
timestamp 1586547711
transform 1 0 19720 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL95680x133280
timestamp 1586547711
transform 1 0 19536 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _416_
timestamp 1586547711
transform 1 0 19904 0 1 27056
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL103040x133280
timestamp 1586547711
transform 1 0 21008 0 1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_41
timestamp 1586547711
transform 1 0 20456 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_480
timestamp 1586547711
transform 1 0 20640 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_517
timestamp 1586547711
transform 1 0 20824 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1462
timestamp 1586547711
transform 1 0 22112 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_484
timestamp 1586547711
transform 1 0 22296 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_417
timestamp 1586547711
transform 1 0 22480 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_264
timestamp 1586547711
transform 1 0 22664 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1586547711
transform 1 0 22848 0 1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _896_
timestamp 1586547711
transform 1 0 22940 0 1 27056
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_12  FILL124200x133280
timestamp 1586547711
transform 1 0 25240 0 1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_518
timestamp 1586547711
transform 1 0 25056 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL132480x133280
timestamp 1586547711
transform 1 0 26896 0 1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL129720x133280
timestamp 1586547711
transform 1 0 26344 0 1 27056
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL140760x133280
timestamp 1586547711
transform 1 0 28552 0 1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL136620x133280
timestamp 1586547711
transform 1 0 27724 0 1 27056
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_271
timestamp 1586547711
transform 1 0 26988 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_422
timestamp 1586547711
transform 1 0 27172 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1111
timestamp 1586547711
transform 1 0 27356 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1227
timestamp 1586547711
transform 1 0 27540 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1586547711
transform 1 0 28460 0 1 27056
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL148120x133280
timestamp 1586547711
transform 1 0 30024 0 1 27056
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL153640x133280
timestamp 1586547711
transform 1 0 31128 0 1 27056
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1586547711
transform 1 0 29656 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_169
timestamp 1586547711
transform 1 0 29840 0 1 27056
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1586547711
transform 1 0 31404 0 1 27056
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL1380x136000
timestamp 1586547711
transform 1 0 676 0 -1 28144
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1586547711
transform 1 0 400 0 -1 28144
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1327
timestamp 1586547711
transform 1 0 2608 0 -1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL6900x136000
timestamp 1586547711
transform 1 0 1780 0 -1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL10580x136000
timestamp 1586547711
transform 1 0 2516 0 -1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _690_
timestamp 1586547711
transform 1 0 1872 0 -1 28144
box 0 -48 644 592
use sky130_fd_sc_hd__fill_1  FILL13800x136000
timestamp 1586547711
transform 1 0 3160 0 -1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1586547711
transform 1 0 3252 0 -1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL11960x136000
timestamp 1586547711
transform 1 0 2792 0 -1 28144
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _691_
timestamp 1586547711
transform 1 0 3344 0 -1 28144
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1335
timestamp 1586547711
transform 1 0 3988 0 -1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1343
timestamp 1586547711
transform 1 0 4172 0 -1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1344
timestamp 1586547711
transform 1 0 4448 0 -1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_622
timestamp 1586547711
transform 1 0 4632 0 -1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL19780x136000
timestamp 1586547711
transform 1 0 4356 0 -1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__o21a_4  _696_
timestamp 1586547711
transform 1 0 4816 0 -1 28144
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL27600x136000
timestamp 1586547711
transform 1 0 5920 0 -1 28144
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILL33120x136000
timestamp 1586547711
transform 1 0 7024 0 -1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1278
timestamp 1586547711
transform 1 0 7208 0 -1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1352
timestamp 1586547711
transform 1 0 7392 0 -1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1347
timestamp 1586547711
transform 1 0 8036 0 -1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL37720x136000
timestamp 1586547711
transform 1 0 7944 0 -1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL41860x136000
timestamp 1586547711
transform 1 0 8772 0 -1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1586547711
transform 1 0 8864 0 -1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL35880x136000
timestamp 1586547711
transform 1 0 7576 0 -1 28144
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILL39100x136000
timestamp 1586547711
transform 1 0 8220 0 -1 28144
box 0 -48 552 592
use sky130_fd_sc_hd__nor2_4  _706_
timestamp 1586547711
transform 1 0 8956 0 -1 28144
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1348
timestamp 1586547711
transform 1 0 10244 0 -1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL48760x136000
timestamp 1586547711
transform 1 0 10152 0 -1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL50140x136000
timestamp 1586547711
transform 1 0 10428 0 -1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL46920x136000
timestamp 1586547711
transform 1 0 9784 0 -1 28144
box 0 -48 368 592
use sky130_fd_sc_hd__dfrtp_4  _925_
timestamp 1586547711
transform 1 0 10520 0 -1 28144
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_12  FILL61180x136000
timestamp 1586547711
transform 1 0 12636 0 -1 28144
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL66700x136000
timestamp 1586547711
transform 1 0 13740 0 -1 28144
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1375
timestamp 1586547711
transform 1 0 15764 0 -1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1586547711
transform 1 0 14476 0 -1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL70840x136000
timestamp 1586547711
transform 1 0 14568 0 -1 28144
box 0 -48 552 592
use sky130_fd_sc_hd__or2_4  _710_
timestamp 1586547711
transform 1 0 15120 0 -1 28144
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILL82800x136000
timestamp 1586547711
transform 1 0 16960 0 -1 28144
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1533
timestamp 1586547711
transform 1 0 18064 0 -1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL77740x136000
timestamp 1586547711
transform 1 0 15948 0 -1 28144
box 0 -48 552 592
use sky130_fd_sc_hd__inv_4  _438_
timestamp 1586547711
transform 1 0 16500 0 -1 28144
box 0 -48 460 592
use sky130_fd_sc_hd__decap_8  FILL94300x136000
timestamp 1586547711
transform 1 0 19260 0 -1 28144
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_231
timestamp 1586547711
transform 1 0 18892 0 -1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_553
timestamp 1586547711
transform 1 0 19076 0 -1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL92000x136000
timestamp 1586547711
transform 1 0 18800 0 -1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL97980x136000
timestamp 1586547711
transform 1 0 19996 0 -1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1586547711
transform 1 0 20088 0 -1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL89240x136000
timestamp 1586547711
transform 1 0 18248 0 -1 28144
box 0 -48 552 592
use sky130_fd_sc_hd__inv_4  _420_
timestamp 1586547711
transform 1 0 20180 0 -1 28144
box 0 -48 460 592
use sky130_fd_sc_hd__decap_12  FILL101200x136000
timestamp 1586547711
transform 1 0 20640 0 -1 28144
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL109480x136000
timestamp 1586547711
transform 1 0 22296 0 -1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL106720x136000
timestamp 1586547711
transform 1 0 21744 0 -1 28144
box 0 -48 552 592
use sky130_fd_sc_hd__buf_4  _791_
timestamp 1586547711
transform 1 0 22388 0 -1 28144
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL113620x136000
timestamp 1586547711
transform 1 0 23124 0 -1 28144
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_493
timestamp 1586547711
transform 1 0 22940 0 -1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL119140x136000
timestamp 1586547711
transform 1 0 24228 0 -1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _421_
timestamp 1586547711
transform 1 0 24320 0 -1 28144
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL126960x136000
timestamp 1586547711
transform 1 0 25792 0 -1 28144
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1166
timestamp 1586547711
transform 1 0 24872 0 -1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL126040x136000
timestamp 1586547711
transform 1 0 25608 0 -1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL132480x136000
timestamp 1586547711
transform 1 0 26896 0 -1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1586547711
transform 1 0 25700 0 -1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL123280x136000
timestamp 1586547711
transform 1 0 25056 0 -1 28144
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL141680x136000
timestamp 1586547711
transform 1 0 28736 0 -1 28144
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1112
timestamp 1586547711
transform 1 0 28552 0 -1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL138920x136000
timestamp 1586547711
transform 1 0 28184 0 -1 28144
box 0 -48 368 592
use sky130_fd_sc_hd__a21bo_4  _650_
timestamp 1586547711
transform 1 0 26988 0 -1 28144
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_12  FILL148580x136000
timestamp 1586547711
transform 1 0 30116 0 -1 28144
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL154100x136000
timestamp 1586547711
transform 1 0 31220 0 -1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1586547711
transform 1 0 31312 0 -1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL145360x136000
timestamp 1586547711
transform 1 0 29472 0 -1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _785_
timestamp 1586547711
transform 1 0 29656 0 -1 28144
box 0 -48 460 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1586547711
transform 1 0 31404 0 -1 28144
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1586547711
transform 1 0 400 0 1 28144
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1318
timestamp 1586547711
transform 1 0 1228 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_612
timestamp 1586547711
transform 1 0 1412 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_436
timestamp 1586547711
transform 1 0 1596 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL1380x138720
timestamp 1586547711
transform 1 0 676 0 1 28144
box 0 -48 552 592
use sky130_fd_sc_hd__o22ai_4  _694_
timestamp 1586547711
transform 1 0 1780 0 1 28144
box 0 -48 1472 592
use sky130_fd_sc_hd__diode_2  ANTENNA_215
timestamp 1586547711
transform 1 0 3344 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1316
timestamp 1586547711
transform 1 0 3528 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_541
timestamp 1586547711
transform 1 0 3804 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL14260x138720
timestamp 1586547711
transform 1 0 3252 0 1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL16560x138720
timestamp 1586547711
transform 1 0 3712 0 1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _699_
timestamp 1586547711
transform 1 0 3988 0 1 28144
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA_438
timestamp 1586547711
transform 1 0 5276 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_613
timestamp 1586547711
transform 1 0 5460 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1332
timestamp 1586547711
transform 1 0 5644 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1323
timestamp 1586547711
transform 1 0 5828 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_219
timestamp 1586547711
transform 1 0 6840 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1330
timestamp 1586547711
transform 1 0 7024 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL31740x138720
timestamp 1586547711
transform 1 0 6748 0 1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1586547711
transform 1 0 6012 0 1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _697_
timestamp 1586547711
transform 1 0 6104 0 1 28144
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  FILL34040x138720
timestamp 1586547711
transform 1 0 7208 0 1 28144
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1360
timestamp 1586547711
transform 1 0 7484 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_623
timestamp 1586547711
transform 1 0 7668 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_440
timestamp 1586547711
transform 1 0 7852 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__o22ai_4  _705_
timestamp 1586547711
transform 1 0 8036 0 1 28144
box 0 -48 1472 592
use sky130_fd_sc_hd__diode_2  ANTENNA_224
timestamp 1586547711
transform 1 0 9508 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1342
timestamp 1586547711
transform 1 0 9692 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1346
timestamp 1586547711
transform 1 0 9876 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1345
timestamp 1586547711
transform 1 0 10060 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_223
timestamp 1586547711
transform 1 0 10888 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1338
timestamp 1586547711
transform 1 0 11072 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL54280x138720
timestamp 1586547711
transform 1 0 11256 0 1 28144
box 0 -48 368 592
use sky130_fd_sc_hd__or2_4  _702_
timestamp 1586547711
transform 1 0 10244 0 1 28144
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1569
timestamp 1586547711
transform 1 0 11808 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1611
timestamp 1586547711
transform 1 0 11992 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1602
timestamp 1586547711
transform 1 0 12820 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_505
timestamp 1586547711
transform 1 0 13556 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL56580x138720
timestamp 1586547711
transform 1 0 11716 0 1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL61640x138720
timestamp 1586547711
transform 1 0 12728 0 1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1586547711
transform 1 0 11624 0 1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL58880x138720
timestamp 1586547711
transform 1 0 12176 0 1 28144
box 0 -48 552 592
use sky130_fd_sc_hd__buf_4  _817_
timestamp 1586547711
transform 1 0 13004 0 1 28144
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILL68540x138720
timestamp 1586547711
transform 1 0 14108 0 1 28144
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1536
timestamp 1586547711
transform 1 0 13740 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1601
timestamp 1586547711
transform 1 0 13924 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1377
timestamp 1586547711
transform 1 0 14384 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_235
timestamp 1586547711
transform 1 0 14568 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_240
timestamp 1586547711
transform 1 0 14752 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_450
timestamp 1586547711
transform 1 0 14936 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_551
timestamp 1586547711
transform 1 0 15120 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1374
timestamp 1586547711
transform 1 0 15304 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL75440x138720
timestamp 1586547711
transform 1 0 15488 0 1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _713_
timestamp 1586547711
transform 1 0 15580 0 1 28144
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  FILL80960x138720
timestamp 1586547711
transform 1 0 16592 0 1 28144
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_561
timestamp 1586547711
transform 1 0 16224 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1370
timestamp 1586547711
transform 1 0 16408 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_444
timestamp 1586547711
transform 1 0 16868 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_557
timestamp 1586547711
transform 1 0 17052 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1367
timestamp 1586547711
transform 1 0 17328 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1372
timestamp 1586547711
transform 1 0 17512 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_445
timestamp 1586547711
transform 1 0 17696 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_232
timestamp 1586547711
transform 1 0 17880 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1586547711
transform 1 0 17236 0 1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _915_
timestamp 1586547711
transform 1 0 18064 0 1 28144
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1532
timestamp 1586547711
transform 1 0 20180 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILL104420x138720
timestamp 1586547711
transform 1 0 21284 0 1 28144
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL100740x138720
timestamp 1586547711
transform 1 0 20548 0 1 28144
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1599
timestamp 1586547711
transform 1 0 20364 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_519
timestamp 1586547711
transform 1 0 22112 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_520
timestamp 1586547711
transform 1 0 22296 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL110400x138720
timestamp 1586547711
transform 1 0 22480 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _426_
timestamp 1586547711
transform 1 0 21560 0 1 28144
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_522
timestamp 1586547711
transform 1 0 22664 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1586547711
transform 1 0 22848 0 1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _428_
timestamp 1586547711
transform 1 0 22940 0 1 28144
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_492
timestamp 1586547711
transform 1 0 23492 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_509
timestamp 1586547711
transform 1 0 23676 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1577
timestamp 1586547711
transform 1 0 23860 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL118220x138720
timestamp 1586547711
transform 1 0 24044 0 1 28144
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_418
timestamp 1586547711
transform 1 0 24504 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_265
timestamp 1586547711
transform 1 0 24688 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL120060x138720
timestamp 1586547711
transform 1 0 24412 0 1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILL128340x138720
timestamp 1586547711
transform 1 0 26068 0 1 28144
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_273
timestamp 1586547711
transform 1 0 26896 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL132020x138720
timestamp 1586547711
transform 1 0 26804 0 1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__a21bo_4  _627_
timestamp 1586547711
transform 1 0 24872 0 1 28144
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_3  FILL136160x138720
timestamp 1586547711
transform 1 0 27632 0 1 28144
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_423
timestamp 1586547711
transform 1 0 27080 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_487
timestamp 1586547711
transform 1 0 27264 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1473
timestamp 1586547711
transform 1 0 27448 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1239
timestamp 1586547711
transform 1 0 27908 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_424
timestamp 1586547711
transform 1 0 28092 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_274
timestamp 1586547711
transform 1 0 28276 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1586547711
transform 1 0 28460 0 1 28144
box 0 -48 92 592
use sky130_fd_sc_hd__a21bo_4  _657_
timestamp 1586547711
transform 1 0 28552 0 1 28144
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_12  FILL148580x138720
timestamp 1586547711
transform 1 0 30116 0 1 28144
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_192
timestamp 1586547711
transform 1 0 29748 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_199
timestamp 1586547711
transform 1 0 29932 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL154100x138720
timestamp 1586547711
transform 1 0 31220 0 1 28144
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1586547711
transform 1 0 31404 0 1 28144
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1586547711
transform 1 0 400 0 1 29232
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1586547711
transform 1 0 400 0 -1 29232
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL1380x141440
timestamp 1586547711
transform 1 0 676 0 -1 29232
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_217
timestamp 1586547711
transform 1 0 768 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1547
timestamp 1586547711
transform 1 0 952 0 -1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL1380x144160
timestamp 1586547711
transform 1 0 676 0 1 29232
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL3680x141440
timestamp 1586547711
transform 1 0 1136 0 -1 29232
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL8740x141440
timestamp 1586547711
transform 1 0 2148 0 -1 29232
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1259
timestamp 1586547711
transform 1 0 1780 0 -1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1329
timestamp 1586547711
transform 1 0 1964 0 -1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL6440x141440
timestamp 1586547711
transform 1 0 1688 0 -1 29232
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _922_
timestamp 1586547711
transform 1 0 952 0 1 29232
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1546
timestamp 1586547711
transform 1 0 3068 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1326
timestamp 1586547711
transform 1 0 3252 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1321
timestamp 1586547711
transform 1 0 3436 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_540
timestamp 1586547711
transform 1 0 3620 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1586547711
transform 1 0 3252 0 -1 29232
box 0 -48 92 592
use sky130_fd_sc_hd__inv_4  _689_
timestamp 1586547711
transform 1 0 3344 0 -1 29232
box 0 -48 460 592
use sky130_fd_sc_hd__diode_2  ANTENNA_221
timestamp 1586547711
transform 1 0 4632 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_439
timestamp 1586547711
transform 1 0 4816 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1325
timestamp 1586547711
transform 1 0 3804 0 -1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1319
timestamp 1586547711
transform 1 0 3988 0 -1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1341
timestamp 1586547711
transform 1 0 4172 0 -1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1333
timestamp 1586547711
transform 1 0 4448 0 -1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL19780x141440
timestamp 1586547711
transform 1 0 4356 0 -1 29232
box 0 -48 92 592
use sky130_fd_sc_hd__and3_4  _692_
timestamp 1586547711
transform 1 0 3804 0 1 29232
box 0 -48 828 592
use sky130_fd_sc_hd__o22ai_4  _700_
timestamp 1586547711
transform 1 0 4632 0 -1 29232
box 0 -48 1472 592
use sky130_fd_sc_hd__decap_12  FILL28520x144160
timestamp 1586547711
transform 1 0 6104 0 1 29232
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1554
timestamp 1586547711
transform 1 0 5000 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1686
timestamp 1586547711
transform 1 0 5184 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1336
timestamp 1586547711
transform 1 0 6104 0 -1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL27600x144160
timestamp 1586547711
transform 1 0 5920 0 1 29232
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1586547711
transform 1 0 6012 0 1 29232
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL24840x144160
timestamp 1586547711
transform 1 0 5368 0 1 29232
box 0 -48 552 592
use sky130_fd_sc_hd__decap_6  FILL29440x141440
timestamp 1586547711
transform 1 0 6288 0 -1 29232
box 0 -48 552 592
use sky130_fd_sc_hd__inv_4  _695_
timestamp 1586547711
transform 1 0 6840 0 -1 29232
box 0 -48 460 592
use sky130_fd_sc_hd__decap_8  FILL34500x141440
timestamp 1586547711
transform 1 0 7300 0 -1 29232
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_181
timestamp 1586547711
transform 1 0 7668 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _698_
timestamp 1586547711
transform 1 0 7208 0 1 29232
box 0 -48 460 592
use sky130_fd_sc_hd__decap_8  FILL39100x144160
timestamp 1586547711
transform 1 0 8220 0 1 29232
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1337
timestamp 1586547711
transform 1 0 7852 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1340
timestamp 1586547711
transform 1 0 8036 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1285
timestamp 1586547711
transform 1 0 8036 0 -1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL39100x141440
timestamp 1586547711
transform 1 0 8220 0 -1 29232
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_225
timestamp 1586547711
transform 1 0 8956 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_441
timestamp 1586547711
transform 1 0 9140 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL41860x141440
timestamp 1586547711
transform 1 0 8772 0 -1 29232
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1586547711
transform 1 0 8864 0 -1 29232
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _703_
timestamp 1586547711
transform 1 0 8956 0 -1 29232
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  FILL46460x144160
timestamp 1586547711
transform 1 0 9692 0 1 29232
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1562
timestamp 1586547711
transform 1 0 9324 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1687
timestamp 1586547711
transform 1 0 9508 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1351
timestamp 1586547711
transform 1 0 9600 0 -1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL46920x141440
timestamp 1586547711
transform 1 0 9784 0 -1 29232
box 0 -48 552 592
use sky130_fd_sc_hd__buf_4  _825_
timestamp 1586547711
transform 1 0 9968 0 1 29232
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1561
timestamp 1586547711
transform 1 0 10520 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1610
timestamp 1586547711
transform 1 0 10704 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__inv_4  _701_
timestamp 1586547711
transform 1 0 10336 0 -1 29232
box 0 -48 460 592
use sky130_fd_sc_hd__decap_8  FILL52440x144160
timestamp 1586547711
transform 1 0 10888 0 1 29232
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL51980x141440
timestamp 1586547711
transform 1 0 10796 0 -1 29232
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILL55660x141440
timestamp 1586547711
transform 1 0 11532 0 -1 29232
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL59800x141440
timestamp 1586547711
transform 1 0 12360 0 -1 29232
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_190
timestamp 1586547711
transform 1 0 11992 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1607
timestamp 1586547711
transform 1 0 12268 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_506
timestamp 1586547711
transform 1 0 12452 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL58880x144160
timestamp 1586547711
transform 1 0 12176 0 1 29232
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1586547711
transform 1 0 11624 0 1 29232
box 0 -48 92 592
use sky130_fd_sc_hd__conb_1  _834_
timestamp 1586547711
transform 1 0 11716 0 1 29232
box 0 -48 276 592
use sky130_fd_sc_hd__buf_4  _826_
timestamp 1586547711
transform 1 0 11808 0 -1 29232
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL66240x141440
timestamp 1586547711
transform 1 0 13648 0 -1 29232
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_451
timestamp 1586547711
transform 1 0 12636 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_243
timestamp 1586547711
transform 1 0 12820 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _816_
timestamp 1586547711
transform 1 0 13096 0 -1 29232
box 0 -48 552 592
use sky130_fd_sc_hd__dfrtp_4  _917_
timestamp 1586547711
transform 1 0 13004 0 1 29232
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1679
timestamp 1586547711
transform 1 0 15488 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1371
timestamp 1586547711
transform 1 0 15672 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL69920x141440
timestamp 1586547711
transform 1 0 14384 0 -1 29232
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1586547711
transform 1 0 14476 0 -1 29232
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL73600x144160
timestamp 1586547711
transform 1 0 15120 0 1 29232
box 0 -48 368 592
use sky130_fd_sc_hd__inv_4  _711_
timestamp 1586547711
transform 1 0 15856 0 1 29232
box 0 -48 460 592
use sky130_fd_sc_hd__a32o_4  _715_
timestamp 1586547711
transform 1 0 14568 0 -1 29232
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA_238
timestamp 1586547711
transform 1 0 16316 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_449
timestamp 1586547711
transform 1 0 16500 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1369
timestamp 1586547711
transform 1 0 16684 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_448
timestamp 1586547711
transform 1 0 16868 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1535
timestamp 1586547711
transform 1 0 16132 0 -1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL79580x141440
timestamp 1586547711
transform 1 0 16316 0 -1 29232
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_234
timestamp 1586547711
transform 1 0 17052 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1376
timestamp 1586547711
transform 1 0 18064 0 -1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1586547711
transform 1 0 17236 0 1 29232
box 0 -48 92 592
use sky130_fd_sc_hd__o21a_4  _714_
timestamp 1586547711
transform 1 0 17328 0 1 29232
box 0 -48 1104 592
use sky130_fd_sc_hd__a21oi_4  _712_
timestamp 1586547711
transform 1 0 16868 0 -1 29232
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1373
timestamp 1586547711
transform 1 0 18432 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1678
timestamp 1586547711
transform 1 0 18248 0 -1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL92000x141440
timestamp 1586547711
transform 1 0 18800 0 -1 29232
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL91080x144160
timestamp 1586547711
transform 1 0 18616 0 1 29232
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILL90160x141440
timestamp 1586547711
transform 1 0 18432 0 -1 29232
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILL94760x141440
timestamp 1586547711
transform 1 0 19352 0 -1 29232
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_179
timestamp 1586547711
transform 1 0 18984 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1595
timestamp 1586547711
transform 1 0 19352 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL93840x144160
timestamp 1586547711
transform 1 0 19168 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _810_
timestamp 1586547711
transform 1 0 19536 0 1 29232
box 0 -48 552 592
use sky130_fd_sc_hd__inv_4  _437_
timestamp 1586547711
transform 1 0 18892 0 -1 29232
box 0 -48 460 592
use sky130_fd_sc_hd__diode_2  ANTENNA_504
timestamp 1586547711
transform 1 0 20088 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL99360x144160
timestamp 1586547711
transform 1 0 20272 0 1 29232
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1586547711
transform 1 0 20088 0 -1 29232
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _814_
timestamp 1586547711
transform 1 0 20180 0 -1 29232
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL106720x144160
timestamp 1586547711
transform 1 0 21744 0 1 29232
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL101660x141440
timestamp 1586547711
transform 1 0 20732 0 -1 29232
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL107180x141440
timestamp 1586547711
transform 1 0 21836 0 -1 29232
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_45
timestamp 1586547711
transform 1 0 20364 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_502
timestamp 1586547711
transform 1 0 20548 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_503
timestamp 1586547711
transform 1 0 21376 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_507
timestamp 1586547711
transform 1 0 21560 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL101660x144160
timestamp 1586547711
transform 1 0 20732 0 1 29232
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _415_
timestamp 1586547711
transform 1 0 20824 0 1 29232
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_521
timestamp 1586547711
transform 1 0 22940 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_182
timestamp 1586547711
transform 1 0 23400 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_490
timestamp 1586547711
transform 1 0 23584 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1586547711
transform 1 0 22848 0 1 29232
box 0 -48 92 592
use sky130_fd_sc_hd__conb_1  _836_
timestamp 1586547711
transform 1 0 23124 0 1 29232
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILL112700x141440
timestamp 1586547711
transform 1 0 22940 0 -1 29232
box 0 -48 552 592
use sky130_fd_sc_hd__buf_4  _792_
timestamp 1586547711
transform 1 0 23492 0 -1 29232
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_267
timestamp 1586547711
transform 1 0 23768 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_198
timestamp 1586547711
transform 1 0 23952 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_491
timestamp 1586547711
transform 1 0 24136 0 -1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_202
timestamp 1586547711
transform 1 0 24320 0 -1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1467
timestamp 1586547711
transform 1 0 24504 0 -1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL118220x141440
timestamp 1586547711
transform 1 0 24044 0 -1 29232
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL121440x141440
timestamp 1586547711
transform 1 0 24688 0 -1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _897_
timestamp 1586547711
transform 1 0 24136 0 1 29232
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_12  FILL126960x141440
timestamp 1586547711
transform 1 0 25792 0 -1 29232
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1109
timestamp 1586547711
transform 1 0 24872 0 -1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL126040x141440
timestamp 1586547711
transform 1 0 25608 0 -1 29232
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1586547711
transform 1 0 25700 0 -1 29232
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL123280x141440
timestamp 1586547711
transform 1 0 25056 0 -1 29232
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1466
timestamp 1586547711
transform 1 0 26252 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1578
timestamp 1586547711
transform 1 0 26436 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1616
timestamp 1586547711
transform 1 0 26804 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILL131100x144160
timestamp 1586547711
transform 1 0 26620 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _899_
timestamp 1586547711
transform 1 0 26896 0 -1 29232
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_3  FILL143060x141440
timestamp 1586547711
transform 1 0 29012 0 -1 29232
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_486
timestamp 1586547711
transform 1 0 27540 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1580
timestamp 1586547711
transform 1 0 27724 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1472
timestamp 1586547711
transform 1 0 27908 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_425
timestamp 1586547711
transform 1 0 28092 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_276
timestamp 1586547711
transform 1 0 28276 0 1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1586547711
transform 1 0 28460 0 1 29232
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _900_
timestamp 1586547711
transform 1 0 28552 0 1 29232
box 0 -48 2116 592
use sky130_fd_sc_hd__buf_4  _424_
timestamp 1586547711
transform 1 0 26988 0 1 29232
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL148580x141440
timestamp 1586547711
transform 1 0 30116 0 -1 29232
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL151340x144160
timestamp 1586547711
transform 1 0 30668 0 1 29232
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1474
timestamp 1586547711
transform 1 0 29288 0 -1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1581
timestamp 1586547711
transform 1 0 29472 0 -1 29232
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL146280x141440
timestamp 1586547711
transform 1 0 29656 0 -1 29232
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILL154100x141440
timestamp 1586547711
transform 1 0 31220 0 -1 29232
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1586547711
transform 1 0 31312 0 -1 29232
box 0 -48 92 592
use sky130_fd_sc_hd__buf_2  _852_
timestamp 1586547711
transform 1 0 29748 0 -1 29232
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1586547711
transform 1 0 31404 0 1 29232
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1586547711
transform 1 0 31404 0 -1 29232
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL4600x146880
timestamp 1586547711
transform 1 0 1320 0 -1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1586547711
transform 1 0 400 0 -1 30320
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILL1380x146880
timestamp 1586547711
transform 1 0 676 0 -1 30320
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILL10120x146880
timestamp 1586547711
transform 1 0 2424 0 -1 30320
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_437
timestamp 1586547711
transform 1 0 952 0 -1 30320
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1685
timestamp 1586547711
transform 1 0 1136 0 -1 30320
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1608
timestamp 1586547711
transform 1 0 3896 0 -1 30320
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL13800x146880
timestamp 1586547711
transform 1 0 3160 0 -1 30320
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1586547711
transform 1 0 3252 0 -1 30320
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL18400x146880
timestamp 1586547711
transform 1 0 4080 0 -1 30320
box 0 -48 552 592
use sky130_fd_sc_hd__dfrtp_4  _923_
timestamp 1586547711
transform 1 0 4632 0 -1 30320
box 0 -48 2116 592
use sky130_fd_sc_hd__buf_4  _823_
timestamp 1586547711
transform 1 0 3344 0 -1 30320
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILL31740x146880
timestamp 1586547711
transform 1 0 6748 0 -1 30320
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILL36800x146880
timestamp 1586547711
transform 1 0 7760 0 -1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1586547711
transform 1 0 8864 0 -1 30320
box 0 -48 92 592
use sky130_fd_sc_hd__conb_1  _829_
timestamp 1586547711
transform 1 0 7484 0 -1 30320
box 0 -48 276 592
use sky130_fd_sc_hd__dfrtp_4  _924_
timestamp 1586547711
transform 1 0 8956 0 -1 30320
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_12  FILL53360x146880
timestamp 1586547711
transform 1 0 11072 0 -1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL65320x146880
timestamp 1586547711
transform 1 0 13464 0 -1 30320
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1537
timestamp 1586547711
transform 1 0 13096 0 -1 30320
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1680
timestamp 1586547711
transform 1 0 13280 0 -1 30320
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL58880x146880
timestamp 1586547711
transform 1 0 12176 0 -1 30320
box 0 -48 368 592
use sky130_fd_sc_hd__buf_4  _822_
timestamp 1586547711
transform 1 0 12544 0 -1 30320
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL70840x146880
timestamp 1586547711
transform 1 0 14568 0 -1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL69000x146880
timestamp 1586547711
transform 1 0 14200 0 -1 30320
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1586547711
transform 1 0 14476 0 -1 30320
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL76360x146880
timestamp 1586547711
transform 1 0 15672 0 -1 30320
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILL78200x146880
timestamp 1586547711
transform 1 0 16040 0 -1 30320
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _916_
timestamp 1586547711
transform 1 0 16132 0 -1 30320
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_8  FILL89240x146880
timestamp 1586547711
transform 1 0 18248 0 -1 30320
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILL94300x146880
timestamp 1586547711
transform 1 0 19260 0 -1 30320
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILL97980x146880
timestamp 1586547711
transform 1 0 19996 0 -1 30320
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1586547711
transform 1 0 20088 0 -1 30320
box 0 -48 92 592
use sky130_fd_sc_hd__conb_1  _837_
timestamp 1586547711
transform 1 0 18984 0 -1 30320
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILL98900x146880
timestamp 1586547711
transform 1 0 20180 0 -1 30320
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL102120x146880
timestamp 1586547711
transform 1 0 20824 0 -1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL107640x146880
timestamp 1586547711
transform 1 0 21928 0 -1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__inv_4  _414_
timestamp 1586547711
transform 1 0 20364 0 -1 30320
box 0 -48 460 592
use sky130_fd_sc_hd__decap_8  FILL121440x146880
timestamp 1586547711
transform 1 0 24688 0 -1 30320
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_419
timestamp 1586547711
transform 1 0 24136 0 -1 30320
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILL115920x146880
timestamp 1586547711
transform 1 0 23584 0 -1 30320
box 0 -48 552 592
use sky130_fd_sc_hd__buf_4  _427_
timestamp 1586547711
transform 1 0 23032 0 -1 30320
box 0 -48 552 592
use sky130_fd_sc_hd__buf_2  _849_
timestamp 1586547711
transform 1 0 24320 0 -1 30320
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL129720x146880
timestamp 1586547711
transform 1 0 26344 0 -1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILL125120x146880
timestamp 1586547711
transform 1 0 25424 0 -1 30320
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1586547711
transform 1 0 25700 0 -1 30320
box 0 -48 92 592
use sky130_fd_sc_hd__buf_4  _793_
timestamp 1586547711
transform 1 0 25792 0 -1 30320
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1475
timestamp 1586547711
transform 1 0 28552 0 -1 30320
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1622
timestamp 1586547711
transform 1 0 28736 0 -1 30320
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILL142600x146880
timestamp 1586547711
transform 1 0 28920 0 -1 30320
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILL135240x146880
timestamp 1586547711
transform 1 0 27448 0 -1 30320
box 0 -48 552 592
use sky130_fd_sc_hd__buf_4  _795_
timestamp 1586547711
transform 1 0 28000 0 -1 30320
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL147200x146880
timestamp 1586547711
transform 1 0 29840 0 -1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1586547711
transform 1 0 31312 0 -1 30320
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL152720x146880
timestamp 1586547711
transform 1 0 30944 0 -1 30320
box 0 -48 368 592
use sky130_fd_sc_hd__buf_4  _796_
timestamp 1586547711
transform 1 0 29288 0 -1 30320
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1586547711
transform 1 0 31404 0 -1 30320
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL1380x149600
timestamp 1586547711
transform 1 0 676 0 1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL6900x149600
timestamp 1586547711
transform 1 0 1780 0 1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1586547711
transform 1 0 400 0 1 30320
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL12420x149600
timestamp 1586547711
transform 1 0 2884 0 1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL17940x149600
timestamp 1586547711
transform 1 0 3988 0 1 30320
box 0 -48 736 592
use sky130_fd_sc_hd__buf_4  _824_
timestamp 1586547711
transform 1 0 4724 0 1 30320
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL28520x149600
timestamp 1586547711
transform 1 0 6104 0 1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1553
timestamp 1586547711
transform 1 0 5276 0 1 30320
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1609
timestamp 1586547711
transform 1 0 5460 0 1 30320
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1586547711
transform 1 0 6012 0 1 30320
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL26220x149600
timestamp 1586547711
transform 1 0 5644 0 1 30320
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL34040x149600
timestamp 1586547711
transform 1 0 7208 0 1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL39560x149600
timestamp 1586547711
transform 1 0 8312 0 1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL45080x149600
timestamp 1586547711
transform 1 0 9416 0 1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL50600x149600
timestamp 1586547711
transform 1 0 10520 0 1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL56580x149600
timestamp 1586547711
transform 1 0 11716 0 1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL62100x149600
timestamp 1586547711
transform 1 0 12820 0 1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1586547711
transform 1 0 11624 0 1 30320
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL67620x149600
timestamp 1586547711
transform 1 0 13924 0 1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL73140x149600
timestamp 1586547711
transform 1 0 15028 0 1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL78660x149600
timestamp 1586547711
transform 1 0 16132 0 1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1534
timestamp 1586547711
transform 1 0 18064 0 1 30320
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1586547711
transform 1 0 17236 0 1 30320
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILL84640x149600
timestamp 1586547711
transform 1 0 17328 0 1 30320
box 0 -48 184 592
use sky130_fd_sc_hd__buf_4  _815_
timestamp 1586547711
transform 1 0 17512 0 1 30320
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL90160x149600
timestamp 1586547711
transform 1 0 18432 0 1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL98900x149600
timestamp 1586547711
transform 1 0 20180 0 1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1600
timestamp 1586547711
transform 1 0 18248 0 1 30320
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_188
timestamp 1586547711
transform 1 0 19996 0 1 30320
box 0 -48 184 592
use sky130_fd_sc_hd__conb_1  _835_
timestamp 1586547711
transform 1 0 19720 0 1 30320
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILL95680x149600
timestamp 1586547711
transform 1 0 19536 0 1 30320
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILL104420x149600
timestamp 1586547711
transform 1 0 21284 0 1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILL109940x149600
timestamp 1586547711
transform 1 0 22388 0 1 30320
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL112700x149600
timestamp 1586547711
transform 1 0 22940 0 1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL118220x149600
timestamp 1586547711
transform 1 0 24044 0 1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILL111780x149600
timestamp 1586547711
transform 1 0 22756 0 1 30320
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1586547711
transform 1 0 22848 0 1 30320
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL123740x149600
timestamp 1586547711
transform 1 0 25148 0 1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL129260x149600
timestamp 1586547711
transform 1 0 26252 0 1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_176
timestamp 1586547711
transform 1 0 27632 0 1 30320
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1615
timestamp 1586547711
transform 1 0 29104 0 1 30320
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL139840x149600
timestamp 1586547711
transform 1 0 28368 0 1 30320
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1586547711
transform 1 0 28460 0 1 30320
box 0 -48 92 592
use sky130_fd_sc_hd__conb_1  _832_
timestamp 1586547711
transform 1 0 27356 0 1 30320
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILL137080x149600
timestamp 1586547711
transform 1 0 27816 0 1 30320
box 0 -48 552 592
use sky130_fd_sc_hd__buf_4  _423_
timestamp 1586547711
transform 1 0 28552 0 1 30320
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL145360x149600
timestamp 1586547711
transform 1 0 29472 0 1 30320
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILL150880x149600
timestamp 1586547711
transform 1 0 30576 0 1 30320
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1621
timestamp 1586547711
transform 1 0 29288 0 1 30320
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILL154560x149600
timestamp 1586547711
transform 1 0 31312 0 1 30320
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1586547711
transform 1 0 31404 0 1 30320
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL1380x152320
timestamp 1586547711
transform 1 0 676 0 -1 31408
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL6900x152320
timestamp 1586547711
transform 1 0 1780 0 -1 31408
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1586547711
transform 1 0 400 0 -1 31408
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILL14720x152320
timestamp 1586547711
transform 1 0 3344 0 -1 31408
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL20240x152320
timestamp 1586547711
transform 1 0 4448 0 -1 31408
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1586547711
transform 1 0 3252 0 -1 31408
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILL12420x152320
timestamp 1586547711
transform 1 0 2884 0 -1 31408
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILL28980x152320
timestamp 1586547711
transform 1 0 6196 0 -1 31408
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1586547711
transform 1 0 6104 0 -1 31408
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL25760x152320
timestamp 1586547711
transform 1 0 5552 0 -1 31408
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL34500x152320
timestamp 1586547711
transform 1 0 7300 0 -1 31408
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL43240x152320
timestamp 1586547711
transform 1 0 9048 0 -1 31408
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1586547711
transform 1 0 8956 0 -1 31408
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL40020x152320
timestamp 1586547711
transform 1 0 8404 0 -1 31408
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL48760x152320
timestamp 1586547711
transform 1 0 10152 0 -1 31408
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILL54280x152320
timestamp 1586547711
transform 1 0 11256 0 -1 31408
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL57500x152320
timestamp 1586547711
transform 1 0 11900 0 -1 31408
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL63020x152320
timestamp 1586547711
transform 1 0 13004 0 -1 31408
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1586547711
transform 1 0 11808 0 -1 31408
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL71760x152320
timestamp 1586547711
transform 1 0 14752 0 -1 31408
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL77280x152320
timestamp 1586547711
transform 1 0 15856 0 -1 31408
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1586547711
transform 1 0 14660 0 -1 31408
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL68540x152320
timestamp 1586547711
transform 1 0 14108 0 -1 31408
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL86020x152320
timestamp 1586547711
transform 1 0 17604 0 -1 31408
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1586547711
transform 1 0 17512 0 -1 31408
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL82800x152320
timestamp 1586547711
transform 1 0 16960 0 -1 31408
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL91540x152320
timestamp 1586547711
transform 1 0 18708 0 -1 31408
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILL97060x152320
timestamp 1586547711
transform 1 0 19812 0 -1 31408
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL100280x152320
timestamp 1586547711
transform 1 0 20456 0 -1 31408
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL105800x152320
timestamp 1586547711
transform 1 0 21560 0 -1 31408
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1586547711
transform 1 0 20364 0 -1 31408
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILL114540x152320
timestamp 1586547711
transform 1 0 23308 0 -1 31408
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL120060x152320
timestamp 1586547711
transform 1 0 24412 0 -1 31408
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1586547711
transform 1 0 23216 0 -1 31408
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL111320x152320
timestamp 1586547711
transform 1 0 22664 0 -1 31408
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL128800x152320
timestamp 1586547711
transform 1 0 26160 0 -1 31408
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1586547711
transform 1 0 26068 0 -1 31408
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL125580x152320
timestamp 1586547711
transform 1 0 25516 0 -1 31408
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL134320x152320
timestamp 1586547711
transform 1 0 27264 0 -1 31408
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILL143060x152320
timestamp 1586547711
transform 1 0 29012 0 -1 31408
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1586547711
transform 1 0 28920 0 -1 31408
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILL139840x152320
timestamp 1586547711
transform 1 0 28368 0 -1 31408
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILL148580x152320
timestamp 1586547711
transform 1 0 30116 0 -1 31408
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILL154100x152320
timestamp 1586547711
transform 1 0 31220 0 -1 31408
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1586547711
transform 1 0 31404 0 -1 31408
box 0 -48 276 592
<< labels >>
rlabel metal3 s 0 28636 440 28876 4 RSTB
port 0 nsew default input
rlabel metal3 s 0 24556 440 24796 4 SCK
port 1 nsew default input
rlabel metal2 s 27990 0 28102 424 8 SDI
port 2 nsew default input
rlabel metal2 s 20446 31664 20558 32088 6 CSB
port 3 nsew default input
rlabel metal2 s 25230 0 25342 424 8 SDO
port 4 nsew default tristate
rlabel metal3 s 31648 9052 32088 9292 6 sdo_enb
port 5 nsew default tristate
rlabel metal2 s 14926 31664 15038 32088 6 xtal_ena
port 6 nsew default tristate
rlabel metal2 s 21918 31664 22030 32088 6 reg_ena
port 7 nsew default tristate
rlabel metal2 s 5910 0 6022 424 8 pll_dco_ena
port 8 nsew default tristate
rlabel metal2 s 22470 0 22582 424 8 pll_div[4]
port 9 nsew default tristate
rlabel metal2 s 20998 0 21110 424 8 pll_div[3]
port 10 nsew default tristate
rlabel metal3 s 0 14492 440 14732 4 pll_div[2]
port 11 nsew default tristate
rlabel metal3 s 31648 7148 32088 7388 6 pll_div[1]
port 12 nsew default tristate
rlabel metal2 s 24678 31664 24790 32088 6 pll_div[0]
port 13 nsew default tristate
rlabel metal2 s 1126 31664 1238 32088 6 pll_sel[2]
port 14 nsew default tristate
rlabel metal3 s 0 30812 440 31052 4 pll_sel[1]
port 15 nsew default tristate
rlabel metal2 s 18238 0 18350 424 8 pll_sel[0]
port 16 nsew default tristate
rlabel metal2 s 26518 0 26630 424 8 pll_trim[25]
port 17 nsew default tristate
rlabel metal3 s 31648 892 32088 1132 6 pll_trim[24]
port 18 nsew default tristate
rlabel metal2 s 30198 31664 30310 32088 6 pll_trim[23]
port 19 nsew default tristate
rlabel metal2 s 16398 31664 16510 32088 6 pll_trim[22]
port 20 nsew default tristate
rlabel metal2 s 28726 31664 28838 32088 6 pll_trim[21]
port 21 nsew default tristate
rlabel metal3 s 31648 3068 32088 3308 6 pll_trim[20]
port 22 nsew default tristate
rlabel metal2 s 30750 0 30862 424 8 pll_trim[19]
port 23 nsew default tristate
rlabel metal2 s 7198 0 7310 424 8 pll_trim[18]
port 24 nsew default tristate
rlabel metal2 s 9406 31664 9518 32088 6 pll_trim[17]
port 25 nsew default tristate
rlabel metal2 s 3886 31664 3998 32088 6 pll_trim[16]
port 26 nsew default tristate
rlabel metal2 s 29278 0 29390 424 8 pll_trim[15]
port 27 nsew default tristate
rlabel metal2 s 19710 0 19822 424 8 pll_trim[14]
port 28 nsew default tristate
rlabel metal2 s 12718 0 12830 424 8 pll_trim[13]
port 29 nsew default tristate
rlabel metal2 s 8118 31664 8230 32088 6 pll_trim[12]
port 30 nsew default tristate
rlabel metal2 s 31486 31664 31598 32088 6 pll_trim[11]
port 31 nsew default tristate
rlabel metal3 s 0 22652 440 22892 4 pll_trim[10]
port 32 nsew default tristate
rlabel metal2 s 2598 31664 2710 32088 6 pll_trim[9]
port 33 nsew default tristate
rlabel metal2 s 8670 0 8782 424 8 pll_trim[8]
port 34 nsew default tristate
rlabel metal2 s 13638 31664 13750 32088 6 pll_trim[7]
port 35 nsew default tristate
rlabel metal2 s 25966 31664 26078 32088 6 pll_trim[6]
port 36 nsew default tristate
rlabel metal2 s 390 0 502 424 8 pll_trim[5]
port 37 nsew default tristate
rlabel metal3 s 0 18572 440 18812 4 pll_trim[4]
port 38 nsew default tristate
rlabel metal2 s 1678 0 1790 424 8 pll_trim[3]
port 39 nsew default tristate
rlabel metal3 s 31648 17212 32088 17452 6 pll_trim[2]
port 40 nsew default tristate
rlabel metal3 s 0 8236 440 8476 4 pll_trim[1]
port 41 nsew default tristate
rlabel metal3 s 31648 13132 32088 13372 6 pll_trim[0]
port 42 nsew default tristate
rlabel metal3 s 31648 4972 32088 5212 6 pll_bypass
port 43 nsew default tristate
rlabel metal3 s 31648 15308 32088 15548 6 irq
port 44 nsew default tristate
rlabel metal2 s 12166 31664 12278 32088 6 reset
port 45 nsew default tristate
rlabel metal3 s 31648 27548 32088 27788 6 RST
port 46 nsew default tristate
rlabel metal2 s 9958 0 10070 424 8 trap
port 47 nsew default input
rlabel metal2 s 16950 0 17062 424 8 mfgr_id[11]
port 48 nsew default tristate
rlabel metal3 s 0 6332 440 6572 4 mfgr_id[10]
port 49 nsew default tristate
rlabel metal3 s 31648 19388 32088 19628 6 mfgr_id[9]
port 50 nsew default tristate
rlabel metal3 s 31648 23468 32088 23708 6 mfgr_id[8]
port 51 nsew default tristate
rlabel metal3 s 0 2252 440 2492 4 mfgr_id[7]
port 52 nsew default tristate
rlabel metal2 s 27438 31664 27550 32088 6 mfgr_id[6]
port 53 nsew default tristate
rlabel metal2 s 11430 0 11542 424 8 mfgr_id[5]
port 54 nsew default tristate
rlabel metal3 s 0 12316 440 12556 4 mfgr_id[4]
port 55 nsew default tristate
rlabel metal2 s 17686 31664 17798 32088 6 mfgr_id[3]
port 56 nsew default tristate
rlabel metal3 s 0 4156 440 4396 4 mfgr_id[2]
port 57 nsew default tristate
rlabel metal2 s 6646 31664 6758 32088 6 mfgr_id[1]
port 58 nsew default tristate
rlabel metal2 s 23206 31664 23318 32088 6 mfgr_id[0]
port 59 nsew default tristate
rlabel metal2 s 3150 0 3262 424 8 prod_id[7]
port 60 nsew default tristate
rlabel metal2 s 4438 0 4550 424 8 prod_id[6]
port 61 nsew default tristate
rlabel metal2 s 23758 0 23870 424 8 prod_id[5]
port 62 nsew default tristate
rlabel metal3 s 0 16396 440 16636 4 prod_id[4]
port 63 nsew default tristate
rlabel metal2 s 15478 0 15590 424 8 prod_id[3]
port 64 nsew default tristate
rlabel metal2 s 19158 31664 19270 32088 6 prod_id[2]
port 65 nsew default tristate
rlabel metal3 s 0 20476 440 20716 4 prod_id[1]
port 66 nsew default tristate
rlabel metal2 s 10878 31664 10990 32088 6 prod_id[0]
port 67 nsew default tristate
rlabel metal2 s 14190 0 14302 424 8 mask_rev_in[3]
port 68 nsew default input
rlabel metal3 s 31648 25372 32088 25612 6 mask_rev_in[2]
port 69 nsew default input
rlabel metal3 s 31648 11228 32088 11468 6 mask_rev_in[1]
port 70 nsew default input
rlabel metal3 s 31648 21292 32088 21532 6 mask_rev_in[0]
port 71 nsew default input
rlabel metal3 s 31648 29452 32088 29692 6 mask_rev[3]
port 72 nsew default tristate
rlabel metal3 s 0 26732 440 26972 4 mask_rev[2]
port 73 nsew default tristate
rlabel metal3 s 0 10412 440 10652 4 mask_rev[1]
port 74 nsew default tristate
rlabel metal2 s 5358 31664 5470 32088 6 mask_rev[0]
port 75 nsew default tristate
flabel metal4 s 3536 504 3784 728 0 FreeSans 1600 0 0 0 vdd
port 76 nsew
flabel metal4 s 18888 512 19136 736 0 FreeSans 1600 0 0 0 vss
port 77 nsew
<< properties >>
string FIXED_BBOX 0 0 32088 32088
<< end >>
